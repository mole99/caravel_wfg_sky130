// This is the unpowered netlist.
module wfg_top (csb1,
    io_wbs_ack,
    io_wbs_clk,
    io_wbs_cyc,
    io_wbs_rst,
    io_wbs_stb,
    io_wbs_we,
    wfg_drive_spi_cs_no,
    wfg_drive_spi_sclk_o,
    wfg_drive_spi_sdo_o,
    addr1,
    dout1,
    io_oeb,
    io_wbs_adr,
    io_wbs_datrd,
    io_wbs_datwr,
    wfg_drive_pat_dout_o);
 output csb1;
 output io_wbs_ack;
 input io_wbs_clk;
 input io_wbs_cyc;
 input io_wbs_rst;
 input io_wbs_stb;
 input io_wbs_we;
 output wfg_drive_spi_cs_no;
 output wfg_drive_spi_sclk_o;
 output wfg_drive_spi_sdo_o;
 output [9:0] addr1;
 input [31:0] dout1;
 output [10:0] io_oeb;
 input [31:0] io_wbs_adr;
 output [31:0] io_wbs_datrd;
 input [31:0] io_wbs_datwr;
 output [31:0] wfg_drive_pat_dout_o;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire net181;
 wire clknet_leaf_0_io_wbs_clk;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire \wfg_core_top.active_o ;
 wire \wfg_core_top.cfg_subcycle_q[10] ;
 wire \wfg_core_top.cfg_subcycle_q[11] ;
 wire \wfg_core_top.cfg_subcycle_q[12] ;
 wire \wfg_core_top.cfg_subcycle_q[13] ;
 wire \wfg_core_top.cfg_subcycle_q[14] ;
 wire \wfg_core_top.cfg_subcycle_q[15] ;
 wire \wfg_core_top.cfg_subcycle_q[16] ;
 wire \wfg_core_top.cfg_subcycle_q[17] ;
 wire \wfg_core_top.cfg_subcycle_q[18] ;
 wire \wfg_core_top.cfg_subcycle_q[19] ;
 wire \wfg_core_top.cfg_subcycle_q[20] ;
 wire \wfg_core_top.cfg_subcycle_q[21] ;
 wire \wfg_core_top.cfg_subcycle_q[22] ;
 wire \wfg_core_top.cfg_subcycle_q[23] ;
 wire \wfg_core_top.cfg_subcycle_q[8] ;
 wire \wfg_core_top.cfg_subcycle_q[9] ;
 wire \wfg_core_top.cfg_sync_q[0] ;
 wire \wfg_core_top.cfg_sync_q[1] ;
 wire \wfg_core_top.cfg_sync_q[2] ;
 wire \wfg_core_top.cfg_sync_q[3] ;
 wire \wfg_core_top.cfg_sync_q[4] ;
 wire \wfg_core_top.cfg_sync_q[5] ;
 wire \wfg_core_top.cfg_sync_q[6] ;
 wire \wfg_core_top.cfg_sync_q[7] ;
 wire \wfg_core_top.wbs_ack_o ;
 wire \wfg_core_top.wbs_dat_o[0] ;
 wire \wfg_core_top.wbs_dat_o[10] ;
 wire \wfg_core_top.wbs_dat_o[11] ;
 wire \wfg_core_top.wbs_dat_o[12] ;
 wire \wfg_core_top.wbs_dat_o[13] ;
 wire \wfg_core_top.wbs_dat_o[14] ;
 wire \wfg_core_top.wbs_dat_o[15] ;
 wire \wfg_core_top.wbs_dat_o[16] ;
 wire \wfg_core_top.wbs_dat_o[17] ;
 wire \wfg_core_top.wbs_dat_o[18] ;
 wire \wfg_core_top.wbs_dat_o[19] ;
 wire \wfg_core_top.wbs_dat_o[1] ;
 wire \wfg_core_top.wbs_dat_o[20] ;
 wire \wfg_core_top.wbs_dat_o[21] ;
 wire \wfg_core_top.wbs_dat_o[22] ;
 wire \wfg_core_top.wbs_dat_o[23] ;
 wire \wfg_core_top.wbs_dat_o[2] ;
 wire \wfg_core_top.wbs_dat_o[3] ;
 wire \wfg_core_top.wbs_dat_o[4] ;
 wire \wfg_core_top.wbs_dat_o[5] ;
 wire \wfg_core_top.wbs_dat_o[6] ;
 wire \wfg_core_top.wbs_dat_o[7] ;
 wire \wfg_core_top.wbs_dat_o[8] ;
 wire \wfg_core_top.wbs_dat_o[9] ;
 wire \wfg_core_top.wfg_core.subcycle_count[0] ;
 wire \wfg_core_top.wfg_core.subcycle_count[10] ;
 wire \wfg_core_top.wfg_core.subcycle_count[11] ;
 wire \wfg_core_top.wfg_core.subcycle_count[12] ;
 wire \wfg_core_top.wfg_core.subcycle_count[13] ;
 wire \wfg_core_top.wfg_core.subcycle_count[14] ;
 wire \wfg_core_top.wfg_core.subcycle_count[15] ;
 wire \wfg_core_top.wfg_core.subcycle_count[1] ;
 wire \wfg_core_top.wfg_core.subcycle_count[2] ;
 wire \wfg_core_top.wfg_core.subcycle_count[3] ;
 wire \wfg_core_top.wfg_core.subcycle_count[4] ;
 wire \wfg_core_top.wfg_core.subcycle_count[5] ;
 wire \wfg_core_top.wfg_core.subcycle_count[6] ;
 wire \wfg_core_top.wfg_core.subcycle_count[7] ;
 wire \wfg_core_top.wfg_core.subcycle_count[8] ;
 wire \wfg_core_top.wfg_core.subcycle_count[9] ;
 wire \wfg_core_top.wfg_core.subcycle_dly ;
 wire \wfg_core_top.wfg_core.subcycle_pls_cnt[0] ;
 wire \wfg_core_top.wfg_core.subcycle_pls_cnt[1] ;
 wire \wfg_core_top.wfg_core.subcycle_pls_cnt[2] ;
 wire \wfg_core_top.wfg_core.subcycle_pls_cnt[3] ;
 wire \wfg_core_top.wfg_core.subcycle_pls_cnt[4] ;
 wire \wfg_core_top.wfg_core.subcycle_pls_cnt[5] ;
 wire \wfg_core_top.wfg_core.subcycle_pls_cnt[6] ;
 wire \wfg_core_top.wfg_core.subcycle_pls_cnt[7] ;
 wire \wfg_core_top.wfg_core.sync_count[0] ;
 wire \wfg_core_top.wfg_core.sync_count[1] ;
 wire \wfg_core_top.wfg_core.sync_count[2] ;
 wire \wfg_core_top.wfg_core.sync_count[3] ;
 wire \wfg_core_top.wfg_core.sync_count[4] ;
 wire \wfg_core_top.wfg_core.sync_count[5] ;
 wire \wfg_core_top.wfg_core.sync_count[6] ;
 wire \wfg_core_top.wfg_core.sync_count[7] ;
 wire \wfg_core_top.wfg_core.sync_dly ;
 wire \wfg_core_top.wfg_core.temp_subcycle ;
 wire \wfg_core_top.wfg_core.temp_sync ;
 wire \wfg_drive_pat_top.cfg_begin_q[0] ;
 wire \wfg_drive_pat_top.cfg_begin_q[1] ;
 wire \wfg_drive_pat_top.cfg_begin_q[2] ;
 wire \wfg_drive_pat_top.cfg_begin_q[3] ;
 wire \wfg_drive_pat_top.cfg_begin_q[4] ;
 wire \wfg_drive_pat_top.cfg_begin_q[5] ;
 wire \wfg_drive_pat_top.cfg_begin_q[6] ;
 wire \wfg_drive_pat_top.cfg_begin_q[7] ;
 wire \wfg_drive_pat_top.cfg_core_sel_q ;
 wire \wfg_drive_pat_top.cfg_end_q[10] ;
 wire \wfg_drive_pat_top.cfg_end_q[11] ;
 wire \wfg_drive_pat_top.cfg_end_q[12] ;
 wire \wfg_drive_pat_top.cfg_end_q[13] ;
 wire \wfg_drive_pat_top.cfg_end_q[14] ;
 wire \wfg_drive_pat_top.cfg_end_q[15] ;
 wire \wfg_drive_pat_top.cfg_end_q[8] ;
 wire \wfg_drive_pat_top.cfg_end_q[9] ;
 wire \wfg_drive_pat_top.patsel0_low_q[0] ;
 wire \wfg_drive_pat_top.patsel0_low_q[10] ;
 wire \wfg_drive_pat_top.patsel0_low_q[11] ;
 wire \wfg_drive_pat_top.patsel0_low_q[12] ;
 wire \wfg_drive_pat_top.patsel0_low_q[13] ;
 wire \wfg_drive_pat_top.patsel0_low_q[14] ;
 wire \wfg_drive_pat_top.patsel0_low_q[15] ;
 wire \wfg_drive_pat_top.patsel0_low_q[16] ;
 wire \wfg_drive_pat_top.patsel0_low_q[17] ;
 wire \wfg_drive_pat_top.patsel0_low_q[18] ;
 wire \wfg_drive_pat_top.patsel0_low_q[19] ;
 wire \wfg_drive_pat_top.patsel0_low_q[1] ;
 wire \wfg_drive_pat_top.patsel0_low_q[20] ;
 wire \wfg_drive_pat_top.patsel0_low_q[21] ;
 wire \wfg_drive_pat_top.patsel0_low_q[22] ;
 wire \wfg_drive_pat_top.patsel0_low_q[23] ;
 wire \wfg_drive_pat_top.patsel0_low_q[24] ;
 wire \wfg_drive_pat_top.patsel0_low_q[25] ;
 wire \wfg_drive_pat_top.patsel0_low_q[26] ;
 wire \wfg_drive_pat_top.patsel0_low_q[27] ;
 wire \wfg_drive_pat_top.patsel0_low_q[28] ;
 wire \wfg_drive_pat_top.patsel0_low_q[29] ;
 wire \wfg_drive_pat_top.patsel0_low_q[2] ;
 wire \wfg_drive_pat_top.patsel0_low_q[30] ;
 wire \wfg_drive_pat_top.patsel0_low_q[31] ;
 wire \wfg_drive_pat_top.patsel0_low_q[3] ;
 wire \wfg_drive_pat_top.patsel0_low_q[4] ;
 wire \wfg_drive_pat_top.patsel0_low_q[5] ;
 wire \wfg_drive_pat_top.patsel0_low_q[6] ;
 wire \wfg_drive_pat_top.patsel0_low_q[7] ;
 wire \wfg_drive_pat_top.patsel0_low_q[8] ;
 wire \wfg_drive_pat_top.patsel0_low_q[9] ;
 wire \wfg_drive_pat_top.patsel1_high_q[0] ;
 wire \wfg_drive_pat_top.patsel1_high_q[10] ;
 wire \wfg_drive_pat_top.patsel1_high_q[11] ;
 wire \wfg_drive_pat_top.patsel1_high_q[12] ;
 wire \wfg_drive_pat_top.patsel1_high_q[13] ;
 wire \wfg_drive_pat_top.patsel1_high_q[14] ;
 wire \wfg_drive_pat_top.patsel1_high_q[15] ;
 wire \wfg_drive_pat_top.patsel1_high_q[16] ;
 wire \wfg_drive_pat_top.patsel1_high_q[17] ;
 wire \wfg_drive_pat_top.patsel1_high_q[18] ;
 wire \wfg_drive_pat_top.patsel1_high_q[19] ;
 wire \wfg_drive_pat_top.patsel1_high_q[1] ;
 wire \wfg_drive_pat_top.patsel1_high_q[20] ;
 wire \wfg_drive_pat_top.patsel1_high_q[21] ;
 wire \wfg_drive_pat_top.patsel1_high_q[22] ;
 wire \wfg_drive_pat_top.patsel1_high_q[23] ;
 wire \wfg_drive_pat_top.patsel1_high_q[24] ;
 wire \wfg_drive_pat_top.patsel1_high_q[25] ;
 wire \wfg_drive_pat_top.patsel1_high_q[26] ;
 wire \wfg_drive_pat_top.patsel1_high_q[27] ;
 wire \wfg_drive_pat_top.patsel1_high_q[28] ;
 wire \wfg_drive_pat_top.patsel1_high_q[29] ;
 wire \wfg_drive_pat_top.patsel1_high_q[2] ;
 wire \wfg_drive_pat_top.patsel1_high_q[30] ;
 wire \wfg_drive_pat_top.patsel1_high_q[31] ;
 wire \wfg_drive_pat_top.patsel1_high_q[3] ;
 wire \wfg_drive_pat_top.patsel1_high_q[4] ;
 wire \wfg_drive_pat_top.patsel1_high_q[5] ;
 wire \wfg_drive_pat_top.patsel1_high_q[6] ;
 wire \wfg_drive_pat_top.patsel1_high_q[7] ;
 wire \wfg_drive_pat_top.patsel1_high_q[8] ;
 wire \wfg_drive_pat_top.patsel1_high_q[9] ;
 wire \wfg_drive_pat_top.wbs_ack_o ;
 wire \wfg_drive_pat_top.wbs_dat_o[0] ;
 wire \wfg_drive_pat_top.wbs_dat_o[10] ;
 wire \wfg_drive_pat_top.wbs_dat_o[11] ;
 wire \wfg_drive_pat_top.wbs_dat_o[12] ;
 wire \wfg_drive_pat_top.wbs_dat_o[13] ;
 wire \wfg_drive_pat_top.wbs_dat_o[14] ;
 wire \wfg_drive_pat_top.wbs_dat_o[15] ;
 wire \wfg_drive_pat_top.wbs_dat_o[16] ;
 wire \wfg_drive_pat_top.wbs_dat_o[17] ;
 wire \wfg_drive_pat_top.wbs_dat_o[18] ;
 wire \wfg_drive_pat_top.wbs_dat_o[19] ;
 wire \wfg_drive_pat_top.wbs_dat_o[1] ;
 wire \wfg_drive_pat_top.wbs_dat_o[20] ;
 wire \wfg_drive_pat_top.wbs_dat_o[21] ;
 wire \wfg_drive_pat_top.wbs_dat_o[22] ;
 wire \wfg_drive_pat_top.wbs_dat_o[23] ;
 wire \wfg_drive_pat_top.wbs_dat_o[24] ;
 wire \wfg_drive_pat_top.wbs_dat_o[25] ;
 wire \wfg_drive_pat_top.wbs_dat_o[26] ;
 wire \wfg_drive_pat_top.wbs_dat_o[27] ;
 wire \wfg_drive_pat_top.wbs_dat_o[28] ;
 wire \wfg_drive_pat_top.wbs_dat_o[29] ;
 wire \wfg_drive_pat_top.wbs_dat_o[2] ;
 wire \wfg_drive_pat_top.wbs_dat_o[30] ;
 wire \wfg_drive_pat_top.wbs_dat_o[31] ;
 wire \wfg_drive_pat_top.wbs_dat_o[3] ;
 wire \wfg_drive_pat_top.wbs_dat_o[4] ;
 wire \wfg_drive_pat_top.wbs_dat_o[5] ;
 wire \wfg_drive_pat_top.wbs_dat_o[6] ;
 wire \wfg_drive_pat_top.wbs_dat_o[7] ;
 wire \wfg_drive_pat_top.wbs_dat_o[8] ;
 wire \wfg_drive_pat_top.wbs_dat_o[9] ;
 wire \wfg_drive_pat_top.wfg_axis_tready_o ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[0].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[0].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[10].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[10].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[11].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[11].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[12].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[12].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[13].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[13].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[14].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[14].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[15].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[15].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[16].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[16].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[17].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[17].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[18].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[18].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[19].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[19].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[1].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[1].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[20].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[20].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[21].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[21].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[22].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[22].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[23].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[23].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[24].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[24].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[25].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[25].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[26].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[26].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[27].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[27].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[28].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[28].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[29].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[29].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[2].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[2].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[30].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[30].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[31].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[31].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[3].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[3].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[4].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[4].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[5].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[5].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[6].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[6].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[7].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[7].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[8].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[8].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[9].drv.axis_data_ff ;
 wire \wfg_drive_pat_top.wfg_drive_pat.gen_channels[9].drv.ctrl_en_q_i ;
 wire \wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[0] ;
 wire \wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[1] ;
 wire \wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[2] ;
 wire \wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[3] ;
 wire \wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[4] ;
 wire \wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[5] ;
 wire \wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[6] ;
 wire \wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[7] ;
 wire \wfg_drive_pat_top.wfg_drive_pat.wfg_sync_i ;
 wire \wfg_drive_spi_top.cfg_core_sel_q ;
 wire \wfg_drive_spi_top.cfg_cpol_q ;
 wire \wfg_drive_spi_top.cfg_dff_q[2] ;
 wire \wfg_drive_spi_top.cfg_dff_q[3] ;
 wire \wfg_drive_spi_top.cfg_lsbfirst_q ;
 wire \wfg_drive_spi_top.cfg_sspol_q ;
 wire \wfg_drive_spi_top.clkcfg_div_q[0] ;
 wire \wfg_drive_spi_top.clkcfg_div_q[1] ;
 wire \wfg_drive_spi_top.clkcfg_div_q[2] ;
 wire \wfg_drive_spi_top.clkcfg_div_q[3] ;
 wire \wfg_drive_spi_top.clkcfg_div_q[4] ;
 wire \wfg_drive_spi_top.clkcfg_div_q[5] ;
 wire \wfg_drive_spi_top.clkcfg_div_q[6] ;
 wire \wfg_drive_spi_top.clkcfg_div_q[7] ;
 wire \wfg_drive_spi_top.ctrl_en_q ;
 wire \wfg_drive_spi_top.wbs_ack_o ;
 wire \wfg_drive_spi_top.wbs_dat_o[0] ;
 wire \wfg_drive_spi_top.wbs_dat_o[1] ;
 wire \wfg_drive_spi_top.wbs_dat_o[2] ;
 wire \wfg_drive_spi_top.wbs_dat_o[3] ;
 wire \wfg_drive_spi_top.wbs_dat_o[4] ;
 wire \wfg_drive_spi_top.wbs_dat_o[5] ;
 wire \wfg_drive_spi_top.wbs_dat_o[6] ;
 wire \wfg_drive_spi_top.wbs_dat_o[7] ;
 wire \wfg_drive_spi_top.wfg_axis_tready_o ;
 wire \wfg_drive_spi_top.wfg_drive_spi.byte_cnt[0] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.byte_cnt[1] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.clk_div[0] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.clk_div[1] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.clk_div[2] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.clk_div[3] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.clk_div[4] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.clk_div[5] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.clk_div[6] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.clk_div[7] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.counter[0] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.counter[1] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.counter[2] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.counter[3] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.counter[4] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.counter[5] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.counter[6] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.counter[7] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.cpol ;
 wire \wfg_drive_spi_top.wfg_drive_spi.cspol ;
 wire \wfg_drive_spi_top.wfg_drive_spi.cur_state[0] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.cur_state[1] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.current_bit[0] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.current_bit[1] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.current_bit[2] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.current_bit[3] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.current_bit[4] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.lsbfirst ;
 wire \wfg_drive_spi_top.wfg_drive_spi.next_state[0] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.next_state[1] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_clk ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_cs ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[0] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[10] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[11] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[12] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[13] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[14] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[15] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[16] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[17] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[18] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[19] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[1] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[20] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[21] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[22] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[23] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[24] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[25] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[26] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[27] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[28] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[29] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[2] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[30] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[31] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[3] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[4] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[5] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[6] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[7] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[8] ;
 wire \wfg_drive_spi_top.wfg_drive_spi.spi_data[9] ;
 wire \wfg_interconnect_top.ctrl_en_q ;
 wire \wfg_interconnect_top.driver0_select_q[0] ;
 wire \wfg_interconnect_top.driver0_select_q[1] ;
 wire \wfg_interconnect_top.driver1_select_q[0] ;
 wire \wfg_interconnect_top.driver1_select_q[1] ;
 wire \wfg_interconnect_top.stimulus_0[0] ;
 wire \wfg_interconnect_top.stimulus_0[10] ;
 wire \wfg_interconnect_top.stimulus_0[11] ;
 wire \wfg_interconnect_top.stimulus_0[12] ;
 wire \wfg_interconnect_top.stimulus_0[13] ;
 wire \wfg_interconnect_top.stimulus_0[14] ;
 wire \wfg_interconnect_top.stimulus_0[15] ;
 wire \wfg_interconnect_top.stimulus_0[16] ;
 wire \wfg_interconnect_top.stimulus_0[17] ;
 wire \wfg_interconnect_top.stimulus_0[1] ;
 wire \wfg_interconnect_top.stimulus_0[2] ;
 wire \wfg_interconnect_top.stimulus_0[32] ;
 wire \wfg_interconnect_top.stimulus_0[3] ;
 wire \wfg_interconnect_top.stimulus_0[4] ;
 wire \wfg_interconnect_top.stimulus_0[5] ;
 wire \wfg_interconnect_top.stimulus_0[6] ;
 wire \wfg_interconnect_top.stimulus_0[7] ;
 wire \wfg_interconnect_top.stimulus_0[8] ;
 wire \wfg_interconnect_top.stimulus_0[9] ;
 wire \wfg_interconnect_top.stimulus_1[0] ;
 wire \wfg_interconnect_top.stimulus_1[10] ;
 wire \wfg_interconnect_top.stimulus_1[11] ;
 wire \wfg_interconnect_top.stimulus_1[12] ;
 wire \wfg_interconnect_top.stimulus_1[13] ;
 wire \wfg_interconnect_top.stimulus_1[14] ;
 wire \wfg_interconnect_top.stimulus_1[15] ;
 wire \wfg_interconnect_top.stimulus_1[16] ;
 wire \wfg_interconnect_top.stimulus_1[17] ;
 wire \wfg_interconnect_top.stimulus_1[18] ;
 wire \wfg_interconnect_top.stimulus_1[19] ;
 wire \wfg_interconnect_top.stimulus_1[1] ;
 wire \wfg_interconnect_top.stimulus_1[20] ;
 wire \wfg_interconnect_top.stimulus_1[21] ;
 wire \wfg_interconnect_top.stimulus_1[22] ;
 wire \wfg_interconnect_top.stimulus_1[23] ;
 wire \wfg_interconnect_top.stimulus_1[24] ;
 wire \wfg_interconnect_top.stimulus_1[25] ;
 wire \wfg_interconnect_top.stimulus_1[26] ;
 wire \wfg_interconnect_top.stimulus_1[27] ;
 wire \wfg_interconnect_top.stimulus_1[28] ;
 wire \wfg_interconnect_top.stimulus_1[29] ;
 wire \wfg_interconnect_top.stimulus_1[2] ;
 wire \wfg_interconnect_top.stimulus_1[30] ;
 wire \wfg_interconnect_top.stimulus_1[31] ;
 wire \wfg_interconnect_top.stimulus_1[32] ;
 wire \wfg_interconnect_top.stimulus_1[3] ;
 wire \wfg_interconnect_top.stimulus_1[4] ;
 wire \wfg_interconnect_top.stimulus_1[5] ;
 wire \wfg_interconnect_top.stimulus_1[6] ;
 wire \wfg_interconnect_top.stimulus_1[7] ;
 wire \wfg_interconnect_top.stimulus_1[8] ;
 wire \wfg_interconnect_top.stimulus_1[9] ;
 wire \wfg_interconnect_top.wbs_ack_o ;
 wire \wfg_interconnect_top.wbs_dat_o[0] ;
 wire \wfg_interconnect_top.wbs_dat_o[1] ;
 wire \wfg_stim_mem_top.cfg_gain_q[10] ;
 wire \wfg_stim_mem_top.cfg_gain_q[11] ;
 wire \wfg_stim_mem_top.cfg_gain_q[12] ;
 wire \wfg_stim_mem_top.cfg_gain_q[13] ;
 wire \wfg_stim_mem_top.cfg_gain_q[14] ;
 wire \wfg_stim_mem_top.cfg_gain_q[15] ;
 wire \wfg_stim_mem_top.cfg_gain_q[16] ;
 wire \wfg_stim_mem_top.cfg_gain_q[17] ;
 wire \wfg_stim_mem_top.cfg_gain_q[18] ;
 wire \wfg_stim_mem_top.cfg_gain_q[19] ;
 wire \wfg_stim_mem_top.cfg_gain_q[20] ;
 wire \wfg_stim_mem_top.cfg_gain_q[21] ;
 wire \wfg_stim_mem_top.cfg_gain_q[22] ;
 wire \wfg_stim_mem_top.cfg_gain_q[23] ;
 wire \wfg_stim_mem_top.cfg_gain_q[8] ;
 wire \wfg_stim_mem_top.cfg_gain_q[9] ;
 wire \wfg_stim_mem_top.cfg_inc_q[0] ;
 wire \wfg_stim_mem_top.cfg_inc_q[1] ;
 wire \wfg_stim_mem_top.cfg_inc_q[2] ;
 wire \wfg_stim_mem_top.cfg_inc_q[3] ;
 wire \wfg_stim_mem_top.cfg_inc_q[4] ;
 wire \wfg_stim_mem_top.cfg_inc_q[5] ;
 wire \wfg_stim_mem_top.cfg_inc_q[6] ;
 wire \wfg_stim_mem_top.cfg_inc_q[7] ;
 wire \wfg_stim_mem_top.ctrl_en_q ;
 wire \wfg_stim_mem_top.end_val_q[0] ;
 wire \wfg_stim_mem_top.end_val_q[10] ;
 wire \wfg_stim_mem_top.end_val_q[11] ;
 wire \wfg_stim_mem_top.end_val_q[12] ;
 wire \wfg_stim_mem_top.end_val_q[13] ;
 wire \wfg_stim_mem_top.end_val_q[14] ;
 wire \wfg_stim_mem_top.end_val_q[15] ;
 wire \wfg_stim_mem_top.end_val_q[1] ;
 wire \wfg_stim_mem_top.end_val_q[2] ;
 wire \wfg_stim_mem_top.end_val_q[3] ;
 wire \wfg_stim_mem_top.end_val_q[4] ;
 wire \wfg_stim_mem_top.end_val_q[5] ;
 wire \wfg_stim_mem_top.end_val_q[6] ;
 wire \wfg_stim_mem_top.end_val_q[7] ;
 wire \wfg_stim_mem_top.end_val_q[8] ;
 wire \wfg_stim_mem_top.end_val_q[9] ;
 wire \wfg_stim_mem_top.start_val_q[0] ;
 wire \wfg_stim_mem_top.start_val_q[10] ;
 wire \wfg_stim_mem_top.start_val_q[11] ;
 wire \wfg_stim_mem_top.start_val_q[12] ;
 wire \wfg_stim_mem_top.start_val_q[13] ;
 wire \wfg_stim_mem_top.start_val_q[14] ;
 wire \wfg_stim_mem_top.start_val_q[15] ;
 wire \wfg_stim_mem_top.start_val_q[1] ;
 wire \wfg_stim_mem_top.start_val_q[2] ;
 wire \wfg_stim_mem_top.start_val_q[3] ;
 wire \wfg_stim_mem_top.start_val_q[4] ;
 wire \wfg_stim_mem_top.start_val_q[5] ;
 wire \wfg_stim_mem_top.start_val_q[6] ;
 wire \wfg_stim_mem_top.start_val_q[7] ;
 wire \wfg_stim_mem_top.start_val_q[8] ;
 wire \wfg_stim_mem_top.start_val_q[9] ;
 wire \wfg_stim_mem_top.wbs_ack_o ;
 wire \wfg_stim_mem_top.wbs_dat_o[0] ;
 wire \wfg_stim_mem_top.wbs_dat_o[10] ;
 wire \wfg_stim_mem_top.wbs_dat_o[11] ;
 wire \wfg_stim_mem_top.wbs_dat_o[12] ;
 wire \wfg_stim_mem_top.wbs_dat_o[13] ;
 wire \wfg_stim_mem_top.wbs_dat_o[14] ;
 wire \wfg_stim_mem_top.wbs_dat_o[15] ;
 wire \wfg_stim_mem_top.wbs_dat_o[16] ;
 wire \wfg_stim_mem_top.wbs_dat_o[17] ;
 wire \wfg_stim_mem_top.wbs_dat_o[18] ;
 wire \wfg_stim_mem_top.wbs_dat_o[19] ;
 wire \wfg_stim_mem_top.wbs_dat_o[1] ;
 wire \wfg_stim_mem_top.wbs_dat_o[20] ;
 wire \wfg_stim_mem_top.wbs_dat_o[21] ;
 wire \wfg_stim_mem_top.wbs_dat_o[22] ;
 wire \wfg_stim_mem_top.wbs_dat_o[23] ;
 wire \wfg_stim_mem_top.wbs_dat_o[2] ;
 wire \wfg_stim_mem_top.wbs_dat_o[3] ;
 wire \wfg_stim_mem_top.wbs_dat_o[4] ;
 wire \wfg_stim_mem_top.wbs_dat_o[5] ;
 wire \wfg_stim_mem_top.wbs_dat_o[6] ;
 wire \wfg_stim_mem_top.wbs_dat_o[7] ;
 wire \wfg_stim_mem_top.wbs_dat_o[8] ;
 wire \wfg_stim_mem_top.wbs_dat_o[9] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.cur_address[10] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.cur_address[11] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.cur_address[12] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.cur_address[13] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.cur_address[14] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.cur_address[15] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.cur_state[0] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.cur_state[1] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.cur_state[2] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.cur_state[3] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[0] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[10] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[11] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[12] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[13] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[14] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[15] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[16] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[17] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[18] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[19] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[1] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[20] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[21] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[22] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[23] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[24] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[25] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[26] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[27] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[28] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[29] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[2] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[30] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[31] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[3] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[4] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[5] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[6] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[7] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[8] ;
 wire \wfg_stim_mem_top.wfg_stim_mem.data_calc[9] ;
 wire \wfg_stim_sine_top.ctrl_en_q ;
 wire \wfg_stim_sine_top.gain_val_q[0] ;
 wire \wfg_stim_sine_top.gain_val_q[10] ;
 wire \wfg_stim_sine_top.gain_val_q[11] ;
 wire \wfg_stim_sine_top.gain_val_q[12] ;
 wire \wfg_stim_sine_top.gain_val_q[13] ;
 wire \wfg_stim_sine_top.gain_val_q[14] ;
 wire \wfg_stim_sine_top.gain_val_q[15] ;
 wire \wfg_stim_sine_top.gain_val_q[1] ;
 wire \wfg_stim_sine_top.gain_val_q[2] ;
 wire \wfg_stim_sine_top.gain_val_q[3] ;
 wire \wfg_stim_sine_top.gain_val_q[4] ;
 wire \wfg_stim_sine_top.gain_val_q[5] ;
 wire \wfg_stim_sine_top.gain_val_q[6] ;
 wire \wfg_stim_sine_top.gain_val_q[7] ;
 wire \wfg_stim_sine_top.gain_val_q[8] ;
 wire \wfg_stim_sine_top.gain_val_q[9] ;
 wire \wfg_stim_sine_top.inc_val_q[0] ;
 wire \wfg_stim_sine_top.inc_val_q[10] ;
 wire \wfg_stim_sine_top.inc_val_q[11] ;
 wire \wfg_stim_sine_top.inc_val_q[12] ;
 wire \wfg_stim_sine_top.inc_val_q[13] ;
 wire \wfg_stim_sine_top.inc_val_q[14] ;
 wire \wfg_stim_sine_top.inc_val_q[15] ;
 wire \wfg_stim_sine_top.inc_val_q[1] ;
 wire \wfg_stim_sine_top.inc_val_q[2] ;
 wire \wfg_stim_sine_top.inc_val_q[3] ;
 wire \wfg_stim_sine_top.inc_val_q[4] ;
 wire \wfg_stim_sine_top.inc_val_q[5] ;
 wire \wfg_stim_sine_top.inc_val_q[6] ;
 wire \wfg_stim_sine_top.inc_val_q[7] ;
 wire \wfg_stim_sine_top.inc_val_q[8] ;
 wire \wfg_stim_sine_top.inc_val_q[9] ;
 wire \wfg_stim_sine_top.offset_val_q[0] ;
 wire \wfg_stim_sine_top.offset_val_q[10] ;
 wire \wfg_stim_sine_top.offset_val_q[11] ;
 wire \wfg_stim_sine_top.offset_val_q[12] ;
 wire \wfg_stim_sine_top.offset_val_q[13] ;
 wire \wfg_stim_sine_top.offset_val_q[14] ;
 wire \wfg_stim_sine_top.offset_val_q[15] ;
 wire \wfg_stim_sine_top.offset_val_q[16] ;
 wire \wfg_stim_sine_top.offset_val_q[17] ;
 wire \wfg_stim_sine_top.offset_val_q[1] ;
 wire \wfg_stim_sine_top.offset_val_q[2] ;
 wire \wfg_stim_sine_top.offset_val_q[3] ;
 wire \wfg_stim_sine_top.offset_val_q[4] ;
 wire \wfg_stim_sine_top.offset_val_q[5] ;
 wire \wfg_stim_sine_top.offset_val_q[6] ;
 wire \wfg_stim_sine_top.offset_val_q[7] ;
 wire \wfg_stim_sine_top.offset_val_q[8] ;
 wire \wfg_stim_sine_top.offset_val_q[9] ;
 wire \wfg_stim_sine_top.wbs_ack_o ;
 wire \wfg_stim_sine_top.wbs_dat_o[0] ;
 wire \wfg_stim_sine_top.wbs_dat_o[10] ;
 wire \wfg_stim_sine_top.wbs_dat_o[11] ;
 wire \wfg_stim_sine_top.wbs_dat_o[12] ;
 wire \wfg_stim_sine_top.wbs_dat_o[13] ;
 wire \wfg_stim_sine_top.wbs_dat_o[14] ;
 wire \wfg_stim_sine_top.wbs_dat_o[15] ;
 wire \wfg_stim_sine_top.wbs_dat_o[16] ;
 wire \wfg_stim_sine_top.wbs_dat_o[17] ;
 wire \wfg_stim_sine_top.wbs_dat_o[1] ;
 wire \wfg_stim_sine_top.wbs_dat_o[2] ;
 wire \wfg_stim_sine_top.wbs_dat_o[3] ;
 wire \wfg_stim_sine_top.wbs_dat_o[4] ;
 wire \wfg_stim_sine_top.wbs_dat_o[5] ;
 wire \wfg_stim_sine_top.wbs_dat_o[6] ;
 wire \wfg_stim_sine_top.wbs_dat_o[7] ;
 wire \wfg_stim_sine_top.wbs_dat_o[8] ;
 wire \wfg_stim_sine_top.wbs_dat_o[9] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.cur_state[0] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.cur_state[1] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.cur_state[2] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.iteration[0] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.iteration[1] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.iteration[2] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.iteration[3] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.overflow_chk[0] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.overflow_chk[10] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.overflow_chk[11] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.overflow_chk[12] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.overflow_chk[13] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.overflow_chk[14] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.overflow_chk[15] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.overflow_chk[16] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.overflow_chk[17] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.overflow_chk[1] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.overflow_chk[2] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.overflow_chk[3] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.overflow_chk[4] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.overflow_chk[5] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.overflow_chk[6] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.overflow_chk[7] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.overflow_chk[8] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.overflow_chk[9] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.phase_in[0] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.phase_in[10] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.phase_in[11] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.phase_in[12] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.phase_in[13] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.phase_in[14] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.phase_in[15] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.phase_in[1] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.phase_in[2] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.phase_in[3] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.phase_in[4] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.phase_in[5] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.phase_in[6] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.phase_in[7] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.phase_in[8] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.phase_in[9] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.quadrant[0] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.quadrant[1] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.sin_17[0] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.sin_17[10] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.sin_17[11] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.sin_17[12] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.sin_17[13] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.sin_17[14] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.sin_17[15] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.sin_17[16] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.sin_17[1] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.sin_17[2] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.sin_17[3] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.sin_17[4] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.sin_17[5] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.sin_17[6] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.sin_17[7] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.sin_17[8] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.sin_17[9] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.temp[14] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.temp[15] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.temp[16] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.temp[17] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.temp[18] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.temp[19] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.temp[20] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.temp[21] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.temp[22] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.temp[23] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.temp[24] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.temp[25] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.temp[26] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.temp[27] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.temp[28] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.temp[29] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.temp[30] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.temp[31] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.x[0] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.x[10] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.x[11] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.x[12] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.x[13] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.x[14] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.x[15] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.x[16] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.x[1] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.x[2] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.x[3] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.x[4] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.x[5] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.x[6] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.x[7] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.x[8] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.x[9] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.y[0] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.y[10] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.y[11] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.y[12] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.y[13] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.y[14] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.y[15] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.y[16] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.y[1] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.y[2] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.y[3] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.y[4] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.y[5] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.y[6] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.y[7] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.y[8] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.y[9] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.z[0] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.z[10] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.z[11] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.z[12] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.z[13] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.z[14] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.z[15] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.z[16] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.z[1] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.z[2] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.z[3] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.z[4] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.z[5] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.z[6] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.z[7] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.z[8] ;
 wire \wfg_stim_sine_top.wfg_stim_sine.z[9] ;
 wire \wfg_subcore_top.active_o ;
 wire \wfg_subcore_top.cfg_subcycle_q[10] ;
 wire \wfg_subcore_top.cfg_subcycle_q[11] ;
 wire \wfg_subcore_top.cfg_subcycle_q[12] ;
 wire \wfg_subcore_top.cfg_subcycle_q[13] ;
 wire \wfg_subcore_top.cfg_subcycle_q[14] ;
 wire \wfg_subcore_top.cfg_subcycle_q[15] ;
 wire \wfg_subcore_top.cfg_subcycle_q[16] ;
 wire \wfg_subcore_top.cfg_subcycle_q[17] ;
 wire \wfg_subcore_top.cfg_subcycle_q[18] ;
 wire \wfg_subcore_top.cfg_subcycle_q[19] ;
 wire \wfg_subcore_top.cfg_subcycle_q[20] ;
 wire \wfg_subcore_top.cfg_subcycle_q[21] ;
 wire \wfg_subcore_top.cfg_subcycle_q[22] ;
 wire \wfg_subcore_top.cfg_subcycle_q[23] ;
 wire \wfg_subcore_top.cfg_subcycle_q[8] ;
 wire \wfg_subcore_top.cfg_subcycle_q[9] ;
 wire \wfg_subcore_top.cfg_sync_q[0] ;
 wire \wfg_subcore_top.cfg_sync_q[1] ;
 wire \wfg_subcore_top.cfg_sync_q[2] ;
 wire \wfg_subcore_top.cfg_sync_q[3] ;
 wire \wfg_subcore_top.cfg_sync_q[4] ;
 wire \wfg_subcore_top.cfg_sync_q[5] ;
 wire \wfg_subcore_top.cfg_sync_q[6] ;
 wire \wfg_subcore_top.cfg_sync_q[7] ;
 wire \wfg_subcore_top.wbs_ack_o ;
 wire \wfg_subcore_top.wbs_dat_o[0] ;
 wire \wfg_subcore_top.wbs_dat_o[10] ;
 wire \wfg_subcore_top.wbs_dat_o[11] ;
 wire \wfg_subcore_top.wbs_dat_o[12] ;
 wire \wfg_subcore_top.wbs_dat_o[13] ;
 wire \wfg_subcore_top.wbs_dat_o[14] ;
 wire \wfg_subcore_top.wbs_dat_o[15] ;
 wire \wfg_subcore_top.wbs_dat_o[16] ;
 wire \wfg_subcore_top.wbs_dat_o[17] ;
 wire \wfg_subcore_top.wbs_dat_o[18] ;
 wire \wfg_subcore_top.wbs_dat_o[19] ;
 wire \wfg_subcore_top.wbs_dat_o[1] ;
 wire \wfg_subcore_top.wbs_dat_o[20] ;
 wire \wfg_subcore_top.wbs_dat_o[21] ;
 wire \wfg_subcore_top.wbs_dat_o[22] ;
 wire \wfg_subcore_top.wbs_dat_o[23] ;
 wire \wfg_subcore_top.wbs_dat_o[2] ;
 wire \wfg_subcore_top.wbs_dat_o[3] ;
 wire \wfg_subcore_top.wbs_dat_o[4] ;
 wire \wfg_subcore_top.wbs_dat_o[5] ;
 wire \wfg_subcore_top.wbs_dat_o[6] ;
 wire \wfg_subcore_top.wbs_dat_o[7] ;
 wire \wfg_subcore_top.wbs_dat_o[8] ;
 wire \wfg_subcore_top.wbs_dat_o[9] ;
 wire \wfg_subcore_top.wfg_subcore.subcycle_count[0] ;
 wire \wfg_subcore_top.wfg_subcore.subcycle_count[10] ;
 wire \wfg_subcore_top.wfg_subcore.subcycle_count[11] ;
 wire \wfg_subcore_top.wfg_subcore.subcycle_count[12] ;
 wire \wfg_subcore_top.wfg_subcore.subcycle_count[13] ;
 wire \wfg_subcore_top.wfg_subcore.subcycle_count[14] ;
 wire \wfg_subcore_top.wfg_subcore.subcycle_count[15] ;
 wire \wfg_subcore_top.wfg_subcore.subcycle_count[1] ;
 wire \wfg_subcore_top.wfg_subcore.subcycle_count[2] ;
 wire \wfg_subcore_top.wfg_subcore.subcycle_count[3] ;
 wire \wfg_subcore_top.wfg_subcore.subcycle_count[4] ;
 wire \wfg_subcore_top.wfg_subcore.subcycle_count[5] ;
 wire \wfg_subcore_top.wfg_subcore.subcycle_count[6] ;
 wire \wfg_subcore_top.wfg_subcore.subcycle_count[7] ;
 wire \wfg_subcore_top.wfg_subcore.subcycle_count[8] ;
 wire \wfg_subcore_top.wfg_subcore.subcycle_count[9] ;
 wire \wfg_subcore_top.wfg_subcore.subcycle_dly ;
 wire \wfg_subcore_top.wfg_subcore.sync_count[0] ;
 wire \wfg_subcore_top.wfg_subcore.sync_count[1] ;
 wire \wfg_subcore_top.wfg_subcore.sync_count[2] ;
 wire \wfg_subcore_top.wfg_subcore.sync_count[3] ;
 wire \wfg_subcore_top.wfg_subcore.sync_count[4] ;
 wire \wfg_subcore_top.wfg_subcore.sync_count[5] ;
 wire \wfg_subcore_top.wfg_subcore.sync_count[6] ;
 wire \wfg_subcore_top.wfg_subcore.sync_count[7] ;
 wire \wfg_subcore_top.wfg_subcore.sync_dly ;
 wire \wfg_subcore_top.wfg_subcore.temp_subcycle ;
 wire \wfg_subcore_top.wfg_subcore.temp_sync ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire clknet_leaf_1_io_wbs_clk;
 wire clknet_leaf_2_io_wbs_clk;
 wire clknet_leaf_3_io_wbs_clk;
 wire clknet_leaf_4_io_wbs_clk;
 wire clknet_leaf_5_io_wbs_clk;
 wire clknet_leaf_6_io_wbs_clk;
 wire clknet_leaf_7_io_wbs_clk;
 wire clknet_leaf_8_io_wbs_clk;
 wire clknet_leaf_9_io_wbs_clk;
 wire clknet_leaf_10_io_wbs_clk;
 wire clknet_leaf_11_io_wbs_clk;
 wire clknet_leaf_12_io_wbs_clk;
 wire clknet_leaf_13_io_wbs_clk;
 wire clknet_leaf_14_io_wbs_clk;
 wire clknet_leaf_15_io_wbs_clk;
 wire clknet_leaf_16_io_wbs_clk;
 wire clknet_leaf_17_io_wbs_clk;
 wire clknet_leaf_18_io_wbs_clk;
 wire clknet_leaf_19_io_wbs_clk;
 wire clknet_leaf_20_io_wbs_clk;
 wire clknet_leaf_21_io_wbs_clk;
 wire clknet_leaf_22_io_wbs_clk;
 wire clknet_leaf_23_io_wbs_clk;
 wire clknet_leaf_24_io_wbs_clk;
 wire clknet_leaf_25_io_wbs_clk;
 wire clknet_leaf_26_io_wbs_clk;
 wire clknet_leaf_27_io_wbs_clk;
 wire clknet_leaf_28_io_wbs_clk;
 wire clknet_leaf_29_io_wbs_clk;
 wire clknet_leaf_31_io_wbs_clk;
 wire clknet_leaf_32_io_wbs_clk;
 wire clknet_leaf_33_io_wbs_clk;
 wire clknet_leaf_34_io_wbs_clk;
 wire clknet_leaf_35_io_wbs_clk;
 wire clknet_leaf_36_io_wbs_clk;
 wire clknet_leaf_37_io_wbs_clk;
 wire clknet_leaf_38_io_wbs_clk;
 wire clknet_leaf_39_io_wbs_clk;
 wire clknet_leaf_40_io_wbs_clk;
 wire clknet_leaf_41_io_wbs_clk;
 wire clknet_leaf_42_io_wbs_clk;
 wire clknet_leaf_43_io_wbs_clk;
 wire clknet_leaf_44_io_wbs_clk;
 wire clknet_leaf_45_io_wbs_clk;
 wire clknet_leaf_46_io_wbs_clk;
 wire clknet_leaf_47_io_wbs_clk;
 wire clknet_leaf_48_io_wbs_clk;
 wire clknet_leaf_49_io_wbs_clk;
 wire clknet_leaf_50_io_wbs_clk;
 wire clknet_leaf_51_io_wbs_clk;
 wire clknet_leaf_52_io_wbs_clk;
 wire clknet_leaf_53_io_wbs_clk;
 wire clknet_leaf_54_io_wbs_clk;
 wire clknet_leaf_55_io_wbs_clk;
 wire clknet_leaf_56_io_wbs_clk;
 wire clknet_leaf_57_io_wbs_clk;
 wire clknet_leaf_58_io_wbs_clk;
 wire clknet_leaf_59_io_wbs_clk;
 wire clknet_leaf_60_io_wbs_clk;
 wire clknet_leaf_61_io_wbs_clk;
 wire clknet_leaf_62_io_wbs_clk;
 wire clknet_leaf_63_io_wbs_clk;
 wire clknet_leaf_64_io_wbs_clk;
 wire clknet_leaf_65_io_wbs_clk;
 wire clknet_leaf_66_io_wbs_clk;
 wire clknet_leaf_67_io_wbs_clk;
 wire clknet_leaf_68_io_wbs_clk;
 wire clknet_leaf_69_io_wbs_clk;
 wire clknet_leaf_70_io_wbs_clk;
 wire clknet_leaf_71_io_wbs_clk;
 wire clknet_leaf_72_io_wbs_clk;
 wire clknet_leaf_73_io_wbs_clk;
 wire clknet_leaf_74_io_wbs_clk;
 wire clknet_leaf_75_io_wbs_clk;
 wire clknet_leaf_76_io_wbs_clk;
 wire clknet_leaf_77_io_wbs_clk;
 wire clknet_leaf_78_io_wbs_clk;
 wire clknet_leaf_79_io_wbs_clk;
 wire clknet_leaf_80_io_wbs_clk;
 wire clknet_leaf_81_io_wbs_clk;
 wire clknet_leaf_82_io_wbs_clk;
 wire clknet_leaf_83_io_wbs_clk;
 wire clknet_leaf_84_io_wbs_clk;
 wire clknet_leaf_85_io_wbs_clk;
 wire clknet_leaf_86_io_wbs_clk;
 wire clknet_leaf_87_io_wbs_clk;
 wire clknet_leaf_88_io_wbs_clk;
 wire clknet_leaf_89_io_wbs_clk;
 wire clknet_leaf_90_io_wbs_clk;
 wire clknet_leaf_91_io_wbs_clk;
 wire clknet_leaf_92_io_wbs_clk;
 wire clknet_leaf_93_io_wbs_clk;
 wire clknet_leaf_94_io_wbs_clk;
 wire clknet_leaf_95_io_wbs_clk;
 wire clknet_leaf_96_io_wbs_clk;
 wire clknet_leaf_97_io_wbs_clk;
 wire clknet_leaf_98_io_wbs_clk;
 wire clknet_leaf_99_io_wbs_clk;
 wire clknet_leaf_100_io_wbs_clk;
 wire clknet_leaf_101_io_wbs_clk;
 wire clknet_leaf_102_io_wbs_clk;
 wire clknet_leaf_103_io_wbs_clk;
 wire clknet_leaf_104_io_wbs_clk;
 wire clknet_leaf_105_io_wbs_clk;
 wire clknet_leaf_106_io_wbs_clk;
 wire clknet_leaf_107_io_wbs_clk;
 wire clknet_leaf_108_io_wbs_clk;
 wire clknet_leaf_109_io_wbs_clk;
 wire clknet_0_io_wbs_clk;
 wire clknet_1_0_0_io_wbs_clk;
 wire clknet_1_0_1_io_wbs_clk;
 wire clknet_1_1_0_io_wbs_clk;
 wire clknet_1_1_1_io_wbs_clk;
 wire clknet_2_0_0_io_wbs_clk;
 wire clknet_2_1_0_io_wbs_clk;
 wire clknet_2_2_0_io_wbs_clk;
 wire clknet_2_3_0_io_wbs_clk;
 wire clknet_3_0_0_io_wbs_clk;
 wire clknet_3_1_0_io_wbs_clk;
 wire clknet_3_2_0_io_wbs_clk;
 wire clknet_3_3_0_io_wbs_clk;
 wire clknet_3_4_0_io_wbs_clk;
 wire clknet_3_5_0_io_wbs_clk;
 wire clknet_3_6_0_io_wbs_clk;
 wire clknet_3_7_0_io_wbs_clk;
 wire clknet_opt_1_0_io_wbs_clk;
 wire clknet_opt_2_0_io_wbs_clk;
 wire clknet_opt_3_0_io_wbs_clk;
 wire clknet_opt_4_0_io_wbs_clk;

 sky130_fd_sc_hd__inv_2 _10050_ (.A(\wfg_drive_spi_top.wfg_drive_spi.cur_state[1] ),
    .Y(_02696_));
 sky130_fd_sc_hd__or2_1 _10051_ (.A(\wfg_drive_spi_top.wfg_drive_spi.counter[1] ),
    .B(\wfg_drive_spi_top.wfg_drive_spi.counter[0] ),
    .X(_02697_));
 sky130_fd_sc_hd__or3_1 _10052_ (.A(\wfg_drive_spi_top.wfg_drive_spi.counter[3] ),
    .B(\wfg_drive_spi_top.wfg_drive_spi.counter[2] ),
    .C(_02697_),
    .X(_02698_));
 sky130_fd_sc_hd__or3_1 _10053_ (.A(\wfg_drive_spi_top.wfg_drive_spi.counter[5] ),
    .B(\wfg_drive_spi_top.wfg_drive_spi.counter[4] ),
    .C(_02698_),
    .X(_02699_));
 sky130_fd_sc_hd__or3_4 _10054_ (.A(\wfg_drive_spi_top.wfg_drive_spi.counter[7] ),
    .B(\wfg_drive_spi_top.wfg_drive_spi.counter[6] ),
    .C(_02699_),
    .X(_02700_));
 sky130_fd_sc_hd__or3_1 _10055_ (.A(\wfg_drive_spi_top.wfg_drive_spi.current_bit[2] ),
    .B(\wfg_drive_spi_top.wfg_drive_spi.current_bit[1] ),
    .C(\wfg_drive_spi_top.wfg_drive_spi.current_bit[0] ),
    .X(_02701_));
 sky130_fd_sc_hd__or2_1 _10056_ (.A(\wfg_drive_spi_top.wfg_drive_spi.current_bit[3] ),
    .B(_02701_),
    .X(_02702_));
 sky130_fd_sc_hd__or4b_2 _10057_ (.A(\wfg_drive_spi_top.wfg_drive_spi.current_bit[4] ),
    .B(_02700_),
    .C(_02702_),
    .D_N(\wfg_drive_spi_top.wfg_drive_spi.spi_clk ),
    .X(_02703_));
 sky130_fd_sc_hd__clkinv_4 _10058_ (.A(\wfg_interconnect_top.driver0_select_q[0] ),
    .Y(_02704_));
 sky130_fd_sc_hd__nor2_2 _10059_ (.A(\wfg_drive_spi_top.wfg_drive_spi.cur_state[1] ),
    .B(\wfg_drive_spi_top.wfg_drive_spi.cur_state[0] ),
    .Y(_02705_));
 sky130_fd_sc_hd__clkinv_2 _10060_ (.A(\wfg_interconnect_top.driver0_select_q[1] ),
    .Y(_02706_));
 sky130_fd_sc_hd__o2111a_1 _10061_ (.A1(_02704_),
    .A2(\wfg_interconnect_top.stimulus_1[32] ),
    .B1(_02705_),
    .C1(_02706_),
    .D1(\wfg_drive_spi_top.ctrl_en_q ),
    .X(_02707_));
 sky130_fd_sc_hd__and2b_1 _10062_ (.A_N(\wfg_core_top.wfg_core.sync_dly ),
    .B(\wfg_core_top.wfg_core.temp_sync ),
    .X(_02708_));
 sky130_fd_sc_hd__and2b_1 _10063_ (.A_N(\wfg_subcore_top.wfg_subcore.sync_dly ),
    .B(\wfg_subcore_top.wfg_subcore.temp_sync ),
    .X(_02709_));
 sky130_fd_sc_hd__mux2_1 _10064_ (.A0(_02708_),
    .A1(_02709_),
    .S(\wfg_drive_spi_top.cfg_core_sel_q ),
    .X(_02710_));
 sky130_fd_sc_hd__o311a_4 _10065_ (.A1(\wfg_interconnect_top.driver0_select_q[1] ),
    .A2(\wfg_interconnect_top.driver0_select_q[0] ),
    .A3(\wfg_interconnect_top.stimulus_0[32] ),
    .B1(_02707_),
    .C1(_02710_),
    .X(_02711_));
 sky130_fd_sc_hd__a31oi_4 _10066_ (.A1(_02696_),
    .A2(\wfg_drive_spi_top.wfg_drive_spi.cur_state[0] ),
    .A3(_02703_),
    .B1(_02711_),
    .Y(_02712_));
 sky130_fd_sc_hd__inv_2 _10067_ (.A(_02712_),
    .Y(\wfg_drive_spi_top.wfg_drive_spi.next_state[0] ));
 sky130_fd_sc_hd__inv_2 _10068_ (.A(\wfg_drive_spi_top.wfg_drive_spi.cur_state[0] ),
    .Y(_02713_));
 sky130_fd_sc_hd__nand2_1 _10069_ (.A(_02696_),
    .B(\wfg_drive_spi_top.wfg_drive_spi.cur_state[0] ),
    .Y(_02714_));
 sky130_fd_sc_hd__nor2_1 _10070_ (.A(_02703_),
    .B(_02714_),
    .Y(_02715_));
 sky130_fd_sc_hd__a31o_1 _10071_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.cur_state[1] ),
    .A2(_02713_),
    .A3(_02700_),
    .B1(_02715_),
    .X(\wfg_drive_spi_top.wfg_drive_spi.next_state[1] ));
 sky130_fd_sc_hd__or2_2 _10072_ (.A(\wfg_drive_spi_top.wfg_drive_spi.next_state[0] ),
    .B(\wfg_drive_spi_top.wfg_drive_spi.next_state[1] ),
    .X(_02716_));
 sky130_fd_sc_hd__clkbuf_2 _10073_ (.A(_02716_),
    .X(_02717_));
 sky130_fd_sc_hd__buf_4 _10074_ (.A(_02717_),
    .X(_00003_));
 sky130_fd_sc_hd__mux2_1 _10075_ (.A0(\wfg_drive_spi_top.cfg_dff_q[3] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.byte_cnt[1] ),
    .S(_00003_),
    .X(_02718_));
 sky130_fd_sc_hd__clkbuf_1 _10076_ (.A(_02718_),
    .X(_01253_));
 sky130_fd_sc_hd__clkbuf_8 _10077_ (.A(_02717_),
    .X(_02719_));
 sky130_fd_sc_hd__mux2_1 _10078_ (.A0(\wfg_drive_spi_top.cfg_dff_q[2] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.byte_cnt[0] ),
    .S(_02719_),
    .X(_02720_));
 sky130_fd_sc_hd__clkbuf_1 _10079_ (.A(_02720_),
    .X(_01252_));
 sky130_fd_sc_hd__mux2_1 _10080_ (.A0(\wfg_drive_spi_top.cfg_sspol_q ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.cspol ),
    .S(_02719_),
    .X(_02721_));
 sky130_fd_sc_hd__clkbuf_1 _10081_ (.A(_02721_),
    .X(_01251_));
 sky130_fd_sc_hd__mux2_1 _10082_ (.A0(\wfg_drive_spi_top.cfg_cpol_q ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.cpol ),
    .S(_02719_),
    .X(_02722_));
 sky130_fd_sc_hd__clkbuf_1 _10083_ (.A(_02722_),
    .X(_01250_));
 sky130_fd_sc_hd__buf_4 _10084_ (.A(\wfg_drive_spi_top.wfg_drive_spi.lsbfirst ),
    .X(_02723_));
 sky130_fd_sc_hd__mux2_1 _10085_ (.A0(\wfg_drive_spi_top.cfg_lsbfirst_q ),
    .A1(_02723_),
    .S(_02719_),
    .X(_02724_));
 sky130_fd_sc_hd__clkbuf_1 _10086_ (.A(_02724_),
    .X(_01249_));
 sky130_fd_sc_hd__mux2_1 _10087_ (.A0(\wfg_drive_spi_top.wfg_axis_tready_o ),
    .A1(_02705_),
    .S(_02719_),
    .X(_02725_));
 sky130_fd_sc_hd__clkbuf_1 _10088_ (.A(_02725_),
    .X(_01248_));
 sky130_fd_sc_hd__nor2_1 _10089_ (.A(\wfg_drive_spi_top.wfg_drive_spi.spi_clk ),
    .B(_02714_),
    .Y(_02726_));
 sky130_fd_sc_hd__inv_2 _10090_ (.A(_02700_),
    .Y(_02727_));
 sky130_fd_sc_hd__a21oi_1 _10091_ (.A1(_02713_),
    .A2(_02700_),
    .B1(_02696_),
    .Y(_02728_));
 sky130_fd_sc_hd__or3_4 _10092_ (.A(_02711_),
    .B(_02715_),
    .C(_02728_),
    .X(_02729_));
 sky130_fd_sc_hd__nor2_4 _10093_ (.A(_02727_),
    .B(_02729_),
    .Y(_02730_));
 sky130_fd_sc_hd__a21oi_1 _10094_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.next_state[0] ),
    .A2(_02730_),
    .B1(_02711_),
    .Y(_02731_));
 sky130_fd_sc_hd__mux2_1 _10095_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_clk ),
    .A1(_02726_),
    .S(_02731_),
    .X(_02732_));
 sky130_fd_sc_hd__clkbuf_1 _10096_ (.A(_02732_),
    .X(_01247_));
 sky130_fd_sc_hd__nor3_2 _10097_ (.A(_02711_),
    .B(_02715_),
    .C(_02728_),
    .Y(_02733_));
 sky130_fd_sc_hd__a31o_1 _10098_ (.A1(_02700_),
    .A2(\wfg_drive_spi_top.wfg_drive_spi.next_state[0] ),
    .A3(_02733_),
    .B1(_02726_),
    .X(_02734_));
 sky130_fd_sc_hd__buf_4 _10099_ (.A(_02734_),
    .X(_02735_));
 sky130_fd_sc_hd__clkbuf_4 _10100_ (.A(_02735_),
    .X(_02736_));
 sky130_fd_sc_hd__nor2_4 _10101_ (.A(_02712_),
    .B(_02735_),
    .Y(_02737_));
 sky130_fd_sc_hd__clkbuf_4 _10102_ (.A(_02737_),
    .X(_02738_));
 sky130_fd_sc_hd__inv_2 _10103_ (.A(_02723_),
    .Y(_02739_));
 sky130_fd_sc_hd__buf_6 _10104_ (.A(_02733_),
    .X(_02740_));
 sky130_fd_sc_hd__o211a_4 _10105_ (.A1(\wfg_interconnect_top.stimulus_0[17] ),
    .A2(\wfg_interconnect_top.driver0_select_q[0] ),
    .B1(_02729_),
    .C1(_02706_),
    .X(_02741_));
 sky130_fd_sc_hd__buf_2 _10106_ (.A(_02741_),
    .X(_02742_));
 sky130_fd_sc_hd__clkbuf_8 _10107_ (.A(_02704_),
    .X(_02743_));
 sky130_fd_sc_hd__or2_1 _10108_ (.A(\wfg_interconnect_top.stimulus_1[31] ),
    .B(_02743_),
    .X(_02744_));
 sky130_fd_sc_hd__a32o_1 _10109_ (.A1(_02739_),
    .A2(\wfg_drive_spi_top.wfg_drive_spi.spi_data[30] ),
    .A3(_02740_),
    .B1(_02742_),
    .B2(_02744_),
    .X(_02745_));
 sky130_fd_sc_hd__a22o_1 _10110_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[31] ),
    .A2(_02736_),
    .B1(_02738_),
    .B2(_02745_),
    .X(_01246_));
 sky130_fd_sc_hd__or2_1 _10111_ (.A(\wfg_interconnect_top.stimulus_1[30] ),
    .B(_02743_),
    .X(_02746_));
 sky130_fd_sc_hd__mux2_1 _10112_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[29] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[31] ),
    .S(_02723_),
    .X(_02747_));
 sky130_fd_sc_hd__buf_2 _10113_ (.A(_02733_),
    .X(_02748_));
 sky130_fd_sc_hd__buf_6 _10114_ (.A(_02748_),
    .X(_02749_));
 sky130_fd_sc_hd__a22o_1 _10115_ (.A1(_02742_),
    .A2(_02746_),
    .B1(_02747_),
    .B2(_02749_),
    .X(_02750_));
 sky130_fd_sc_hd__a22o_1 _10116_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[30] ),
    .A2(_02736_),
    .B1(_02738_),
    .B2(_02750_),
    .X(_01245_));
 sky130_fd_sc_hd__or2_1 _10117_ (.A(\wfg_interconnect_top.stimulus_1[29] ),
    .B(_02743_),
    .X(_02751_));
 sky130_fd_sc_hd__mux2_1 _10118_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[28] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[30] ),
    .S(_02723_),
    .X(_02752_));
 sky130_fd_sc_hd__a22o_1 _10119_ (.A1(_02742_),
    .A2(_02751_),
    .B1(_02752_),
    .B2(_02749_),
    .X(_02753_));
 sky130_fd_sc_hd__a22o_1 _10120_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[29] ),
    .A2(_02736_),
    .B1(_02738_),
    .B2(_02753_),
    .X(_01244_));
 sky130_fd_sc_hd__or2_1 _10121_ (.A(\wfg_interconnect_top.stimulus_1[28] ),
    .B(_02743_),
    .X(_02754_));
 sky130_fd_sc_hd__mux2_1 _10122_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[27] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[29] ),
    .S(_02723_),
    .X(_02755_));
 sky130_fd_sc_hd__a22o_1 _10123_ (.A1(_02742_),
    .A2(_02754_),
    .B1(_02755_),
    .B2(_02749_),
    .X(_02756_));
 sky130_fd_sc_hd__a22o_1 _10124_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[28] ),
    .A2(_02736_),
    .B1(_02738_),
    .B2(_02756_),
    .X(_01243_));
 sky130_fd_sc_hd__or2_1 _10125_ (.A(\wfg_interconnect_top.stimulus_1[27] ),
    .B(_02743_),
    .X(_02757_));
 sky130_fd_sc_hd__mux2_1 _10126_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[26] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[28] ),
    .S(_02723_),
    .X(_02758_));
 sky130_fd_sc_hd__a22o_1 _10127_ (.A1(_02742_),
    .A2(_02757_),
    .B1(_02758_),
    .B2(_02749_),
    .X(_02759_));
 sky130_fd_sc_hd__a22o_1 _10128_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[27] ),
    .A2(_02736_),
    .B1(_02738_),
    .B2(_02759_),
    .X(_01242_));
 sky130_fd_sc_hd__or2_1 _10129_ (.A(\wfg_interconnect_top.stimulus_1[26] ),
    .B(_02743_),
    .X(_02760_));
 sky130_fd_sc_hd__mux2_1 _10130_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[25] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[27] ),
    .S(_02723_),
    .X(_02761_));
 sky130_fd_sc_hd__a22o_1 _10131_ (.A1(_02742_),
    .A2(_02760_),
    .B1(_02761_),
    .B2(_02749_),
    .X(_02762_));
 sky130_fd_sc_hd__a22o_1 _10132_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[26] ),
    .A2(_02736_),
    .B1(_02738_),
    .B2(_02762_),
    .X(_01241_));
 sky130_fd_sc_hd__or2_1 _10133_ (.A(\wfg_interconnect_top.stimulus_1[25] ),
    .B(_02743_),
    .X(_02763_));
 sky130_fd_sc_hd__mux2_1 _10134_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[24] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[26] ),
    .S(_02723_),
    .X(_02764_));
 sky130_fd_sc_hd__a22o_1 _10135_ (.A1(_02742_),
    .A2(_02763_),
    .B1(_02764_),
    .B2(_02749_),
    .X(_02765_));
 sky130_fd_sc_hd__a22o_1 _10136_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[25] ),
    .A2(_02736_),
    .B1(_02738_),
    .B2(_02765_),
    .X(_01240_));
 sky130_fd_sc_hd__or2_1 _10137_ (.A(\wfg_interconnect_top.stimulus_1[24] ),
    .B(_02743_),
    .X(_02766_));
 sky130_fd_sc_hd__mux2_1 _10138_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[23] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[25] ),
    .S(_02723_),
    .X(_02767_));
 sky130_fd_sc_hd__a22o_1 _10139_ (.A1(_02742_),
    .A2(_02766_),
    .B1(_02767_),
    .B2(_02740_),
    .X(_02768_));
 sky130_fd_sc_hd__a22o_1 _10140_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[24] ),
    .A2(_02736_),
    .B1(_02738_),
    .B2(_02768_),
    .X(_01239_));
 sky130_fd_sc_hd__or2_1 _10141_ (.A(\wfg_interconnect_top.stimulus_1[23] ),
    .B(_02743_),
    .X(_02769_));
 sky130_fd_sc_hd__buf_4 _10142_ (.A(\wfg_drive_spi_top.wfg_drive_spi.lsbfirst ),
    .X(_02770_));
 sky130_fd_sc_hd__mux2_1 _10143_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[22] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[24] ),
    .S(_02770_),
    .X(_02771_));
 sky130_fd_sc_hd__a22o_1 _10144_ (.A1(_02742_),
    .A2(_02769_),
    .B1(_02771_),
    .B2(_02740_),
    .X(_02772_));
 sky130_fd_sc_hd__a22o_1 _10145_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[23] ),
    .A2(_02736_),
    .B1(_02738_),
    .B2(_02772_),
    .X(_01238_));
 sky130_fd_sc_hd__or2_1 _10146_ (.A(\wfg_interconnect_top.stimulus_1[22] ),
    .B(_02704_),
    .X(_02773_));
 sky130_fd_sc_hd__mux2_1 _10147_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[21] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[23] ),
    .S(_02770_),
    .X(_02774_));
 sky130_fd_sc_hd__a22o_1 _10148_ (.A1(_02742_),
    .A2(_02773_),
    .B1(_02774_),
    .B2(_02740_),
    .X(_02775_));
 sky130_fd_sc_hd__a22o_1 _10149_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[22] ),
    .A2(_02736_),
    .B1(_02738_),
    .B2(_02775_),
    .X(_01237_));
 sky130_fd_sc_hd__clkbuf_4 _10150_ (.A(_02735_),
    .X(_02776_));
 sky130_fd_sc_hd__buf_4 _10151_ (.A(_02737_),
    .X(_02777_));
 sky130_fd_sc_hd__or2_1 _10152_ (.A(\wfg_interconnect_top.stimulus_1[21] ),
    .B(_02704_),
    .X(_02778_));
 sky130_fd_sc_hd__mux2_1 _10153_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[20] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[22] ),
    .S(_02770_),
    .X(_02779_));
 sky130_fd_sc_hd__a22o_1 _10154_ (.A1(_02741_),
    .A2(_02778_),
    .B1(_02779_),
    .B2(_02740_),
    .X(_02780_));
 sky130_fd_sc_hd__a22o_1 _10155_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[21] ),
    .A2(_02776_),
    .B1(_02777_),
    .B2(_02780_),
    .X(_01236_));
 sky130_fd_sc_hd__or2_1 _10156_ (.A(\wfg_interconnect_top.stimulus_1[20] ),
    .B(_02704_),
    .X(_02781_));
 sky130_fd_sc_hd__mux2_1 _10157_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[19] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[21] ),
    .S(_02770_),
    .X(_02782_));
 sky130_fd_sc_hd__a22o_1 _10158_ (.A1(_02741_),
    .A2(_02781_),
    .B1(_02782_),
    .B2(_02740_),
    .X(_02783_));
 sky130_fd_sc_hd__a22o_1 _10159_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[20] ),
    .A2(_02776_),
    .B1(_02777_),
    .B2(_02783_),
    .X(_01235_));
 sky130_fd_sc_hd__or2_1 _10160_ (.A(\wfg_interconnect_top.stimulus_1[19] ),
    .B(_02704_),
    .X(_02784_));
 sky130_fd_sc_hd__mux2_1 _10161_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[18] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[20] ),
    .S(_02770_),
    .X(_02785_));
 sky130_fd_sc_hd__a22o_1 _10162_ (.A1(_02741_),
    .A2(_02784_),
    .B1(_02785_),
    .B2(_02740_),
    .X(_02786_));
 sky130_fd_sc_hd__a22o_1 _10163_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[19] ),
    .A2(_02776_),
    .B1(_02777_),
    .B2(_02786_),
    .X(_01234_));
 sky130_fd_sc_hd__or2_1 _10164_ (.A(\wfg_interconnect_top.stimulus_1[18] ),
    .B(_02704_),
    .X(_02787_));
 sky130_fd_sc_hd__mux2_1 _10165_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[17] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[19] ),
    .S(_02770_),
    .X(_02788_));
 sky130_fd_sc_hd__a22o_1 _10166_ (.A1(_02741_),
    .A2(_02787_),
    .B1(_02788_),
    .B2(_02740_),
    .X(_02789_));
 sky130_fd_sc_hd__a22o_1 _10167_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[18] ),
    .A2(_02776_),
    .B1(_02777_),
    .B2(_02789_),
    .X(_01233_));
 sky130_fd_sc_hd__or2_1 _10168_ (.A(\wfg_interconnect_top.stimulus_1[17] ),
    .B(_02704_),
    .X(_02790_));
 sky130_fd_sc_hd__mux2_1 _10169_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[16] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[18] ),
    .S(_02770_),
    .X(_02791_));
 sky130_fd_sc_hd__a22o_1 _10170_ (.A1(_02741_),
    .A2(_02790_),
    .B1(_02791_),
    .B2(_02740_),
    .X(_02792_));
 sky130_fd_sc_hd__a22o_1 _10171_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[17] ),
    .A2(_02776_),
    .B1(_02777_),
    .B2(_02792_),
    .X(_01232_));
 sky130_fd_sc_hd__buf_4 _10172_ (.A(_02729_),
    .X(_02793_));
 sky130_fd_sc_hd__mux2_1 _10173_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[15] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[17] ),
    .S(_02770_),
    .X(_02794_));
 sky130_fd_sc_hd__or2_1 _10174_ (.A(_02793_),
    .B(_02794_),
    .X(_02795_));
 sky130_fd_sc_hd__nor2_8 _10175_ (.A(\wfg_interconnect_top.driver0_select_q[1] ),
    .B(\wfg_interconnect_top.driver0_select_q[0] ),
    .Y(_02796_));
 sky130_fd_sc_hd__buf_2 _10176_ (.A(_02796_),
    .X(_02797_));
 sky130_fd_sc_hd__nor2_4 _10177_ (.A(\wfg_interconnect_top.driver0_select_q[1] ),
    .B(_02704_),
    .Y(_02798_));
 sky130_fd_sc_hd__buf_2 _10178_ (.A(_02798_),
    .X(_02799_));
 sky130_fd_sc_hd__clkbuf_4 _10179_ (.A(_02733_),
    .X(_02800_));
 sky130_fd_sc_hd__a221o_1 _10180_ (.A1(\wfg_interconnect_top.stimulus_0[16] ),
    .A2(_02797_),
    .B1(_02799_),
    .B2(\wfg_interconnect_top.stimulus_1[16] ),
    .C1(_02800_),
    .X(_02801_));
 sky130_fd_sc_hd__a32o_1 _10181_ (.A1(_02777_),
    .A2(_02795_),
    .A3(_02801_),
    .B1(_02776_),
    .B2(\wfg_drive_spi_top.wfg_drive_spi.spi_data[16] ),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _10182_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[14] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[16] ),
    .S(_02770_),
    .X(_02802_));
 sky130_fd_sc_hd__or2_1 _10183_ (.A(_02793_),
    .B(_02802_),
    .X(_02803_));
 sky130_fd_sc_hd__a221o_1 _10184_ (.A1(\wfg_interconnect_top.stimulus_0[15] ),
    .A2(_02797_),
    .B1(_02799_),
    .B2(\wfg_interconnect_top.stimulus_1[15] ),
    .C1(_02800_),
    .X(_02804_));
 sky130_fd_sc_hd__a32o_1 _10185_ (.A1(_02777_),
    .A2(_02803_),
    .A3(_02804_),
    .B1(_02776_),
    .B2(\wfg_drive_spi_top.wfg_drive_spi.spi_data[15] ),
    .X(_01230_));
 sky130_fd_sc_hd__mux2_1 _10186_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[13] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[15] ),
    .S(_02770_),
    .X(_02805_));
 sky130_fd_sc_hd__or2_1 _10187_ (.A(_02793_),
    .B(_02805_),
    .X(_02806_));
 sky130_fd_sc_hd__a221o_1 _10188_ (.A1(\wfg_interconnect_top.stimulus_0[14] ),
    .A2(_02797_),
    .B1(_02799_),
    .B2(\wfg_interconnect_top.stimulus_1[14] ),
    .C1(_02800_),
    .X(_02807_));
 sky130_fd_sc_hd__a32o_1 _10189_ (.A1(_02777_),
    .A2(_02806_),
    .A3(_02807_),
    .B1(_02776_),
    .B2(\wfg_drive_spi_top.wfg_drive_spi.spi_data[14] ),
    .X(_01229_));
 sky130_fd_sc_hd__clkbuf_2 _10190_ (.A(_02729_),
    .X(_02808_));
 sky130_fd_sc_hd__clkbuf_4 _10191_ (.A(\wfg_drive_spi_top.wfg_drive_spi.lsbfirst ),
    .X(_02809_));
 sky130_fd_sc_hd__mux2_1 _10192_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[12] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[14] ),
    .S(_02809_),
    .X(_02810_));
 sky130_fd_sc_hd__or2_1 _10193_ (.A(_02808_),
    .B(_02810_),
    .X(_02811_));
 sky130_fd_sc_hd__a221o_1 _10194_ (.A1(\wfg_interconnect_top.stimulus_0[13] ),
    .A2(_02797_),
    .B1(_02799_),
    .B2(\wfg_interconnect_top.stimulus_1[13] ),
    .C1(_02800_),
    .X(_02812_));
 sky130_fd_sc_hd__a32o_1 _10195_ (.A1(_02777_),
    .A2(_02811_),
    .A3(_02812_),
    .B1(_02776_),
    .B2(\wfg_drive_spi_top.wfg_drive_spi.spi_data[13] ),
    .X(_01228_));
 sky130_fd_sc_hd__clkbuf_4 _10196_ (.A(_02737_),
    .X(_02813_));
 sky130_fd_sc_hd__mux2_1 _10197_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[11] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[13] ),
    .S(_02809_),
    .X(_02814_));
 sky130_fd_sc_hd__or2_1 _10198_ (.A(_02808_),
    .B(_02814_),
    .X(_02815_));
 sky130_fd_sc_hd__a221o_1 _10199_ (.A1(\wfg_interconnect_top.stimulus_0[12] ),
    .A2(_02797_),
    .B1(_02799_),
    .B2(\wfg_interconnect_top.stimulus_1[12] ),
    .C1(_02800_),
    .X(_02816_));
 sky130_fd_sc_hd__a32o_1 _10200_ (.A1(_02813_),
    .A2(_02815_),
    .A3(_02816_),
    .B1(_02776_),
    .B2(\wfg_drive_spi_top.wfg_drive_spi.spi_data[12] ),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _10201_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[10] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[12] ),
    .S(_02809_),
    .X(_02817_));
 sky130_fd_sc_hd__or2_1 _10202_ (.A(_02808_),
    .B(_02817_),
    .X(_02818_));
 sky130_fd_sc_hd__a221o_1 _10203_ (.A1(\wfg_interconnect_top.stimulus_0[11] ),
    .A2(_02797_),
    .B1(_02799_),
    .B2(\wfg_interconnect_top.stimulus_1[11] ),
    .C1(_02800_),
    .X(_02819_));
 sky130_fd_sc_hd__clkbuf_4 _10204_ (.A(_02735_),
    .X(_02820_));
 sky130_fd_sc_hd__a32o_1 _10205_ (.A1(_02813_),
    .A2(_02818_),
    .A3(_02819_),
    .B1(_02820_),
    .B2(\wfg_drive_spi_top.wfg_drive_spi.spi_data[11] ),
    .X(_01226_));
 sky130_fd_sc_hd__mux2_1 _10206_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[9] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[11] ),
    .S(_02809_),
    .X(_02821_));
 sky130_fd_sc_hd__or2_1 _10207_ (.A(_02808_),
    .B(_02821_),
    .X(_02822_));
 sky130_fd_sc_hd__a221o_1 _10208_ (.A1(\wfg_interconnect_top.stimulus_0[10] ),
    .A2(_02797_),
    .B1(_02799_),
    .B2(\wfg_interconnect_top.stimulus_1[10] ),
    .C1(_02800_),
    .X(_02823_));
 sky130_fd_sc_hd__a32o_1 _10209_ (.A1(_02813_),
    .A2(_02822_),
    .A3(_02823_),
    .B1(_02820_),
    .B2(\wfg_drive_spi_top.wfg_drive_spi.spi_data[10] ),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_1 _10210_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[8] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[10] ),
    .S(_02809_),
    .X(_02824_));
 sky130_fd_sc_hd__or2_1 _10211_ (.A(_02808_),
    .B(_02824_),
    .X(_02825_));
 sky130_fd_sc_hd__a221o_1 _10212_ (.A1(\wfg_interconnect_top.stimulus_0[9] ),
    .A2(_02797_),
    .B1(_02799_),
    .B2(\wfg_interconnect_top.stimulus_1[9] ),
    .C1(_02800_),
    .X(_02826_));
 sky130_fd_sc_hd__a32o_1 _10213_ (.A1(_02813_),
    .A2(_02825_),
    .A3(_02826_),
    .B1(_02820_),
    .B2(\wfg_drive_spi_top.wfg_drive_spi.spi_data[9] ),
    .X(_01224_));
 sky130_fd_sc_hd__mux2_1 _10214_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[7] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[9] ),
    .S(_02809_),
    .X(_02827_));
 sky130_fd_sc_hd__or2_1 _10215_ (.A(_02808_),
    .B(_02827_),
    .X(_02828_));
 sky130_fd_sc_hd__a221o_1 _10216_ (.A1(\wfg_interconnect_top.stimulus_0[8] ),
    .A2(_02797_),
    .B1(_02799_),
    .B2(\wfg_interconnect_top.stimulus_1[8] ),
    .C1(_02748_),
    .X(_02829_));
 sky130_fd_sc_hd__a32o_1 _10217_ (.A1(_02813_),
    .A2(_02828_),
    .A3(_02829_),
    .B1(_02820_),
    .B2(\wfg_drive_spi_top.wfg_drive_spi.spi_data[8] ),
    .X(_01223_));
 sky130_fd_sc_hd__mux2_1 _10218_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[6] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[8] ),
    .S(_02809_),
    .X(_02830_));
 sky130_fd_sc_hd__or2_1 _10219_ (.A(_02808_),
    .B(_02830_),
    .X(_02831_));
 sky130_fd_sc_hd__a221o_1 _10220_ (.A1(\wfg_interconnect_top.stimulus_0[7] ),
    .A2(_02797_),
    .B1(_02799_),
    .B2(\wfg_interconnect_top.stimulus_1[7] ),
    .C1(_02748_),
    .X(_02832_));
 sky130_fd_sc_hd__a32o_1 _10221_ (.A1(_02813_),
    .A2(_02831_),
    .A3(_02832_),
    .B1(_02820_),
    .B2(\wfg_drive_spi_top.wfg_drive_spi.spi_data[7] ),
    .X(_01222_));
 sky130_fd_sc_hd__mux2_1 _10222_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[5] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[7] ),
    .S(_02809_),
    .X(_02833_));
 sky130_fd_sc_hd__or2_1 _10223_ (.A(_02808_),
    .B(_02833_),
    .X(_02834_));
 sky130_fd_sc_hd__a221o_1 _10224_ (.A1(\wfg_interconnect_top.stimulus_0[6] ),
    .A2(_02796_),
    .B1(_02798_),
    .B2(\wfg_interconnect_top.stimulus_1[6] ),
    .C1(_02748_),
    .X(_02835_));
 sky130_fd_sc_hd__a32o_1 _10225_ (.A1(_02813_),
    .A2(_02834_),
    .A3(_02835_),
    .B1(_02820_),
    .B2(\wfg_drive_spi_top.wfg_drive_spi.spi_data[6] ),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_1 _10226_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[4] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[6] ),
    .S(_02809_),
    .X(_02836_));
 sky130_fd_sc_hd__or2_1 _10227_ (.A(_02808_),
    .B(_02836_),
    .X(_02837_));
 sky130_fd_sc_hd__a221o_1 _10228_ (.A1(\wfg_interconnect_top.stimulus_0[5] ),
    .A2(_02796_),
    .B1(_02798_),
    .B2(\wfg_interconnect_top.stimulus_1[5] ),
    .C1(_02748_),
    .X(_02838_));
 sky130_fd_sc_hd__a32o_1 _10229_ (.A1(_02813_),
    .A2(_02837_),
    .A3(_02838_),
    .B1(_02820_),
    .B2(\wfg_drive_spi_top.wfg_drive_spi.spi_data[5] ),
    .X(_01220_));
 sky130_fd_sc_hd__mux2_1 _10230_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[3] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[5] ),
    .S(_02809_),
    .X(_02839_));
 sky130_fd_sc_hd__or2_1 _10231_ (.A(_02808_),
    .B(_02839_),
    .X(_02840_));
 sky130_fd_sc_hd__a221o_1 _10232_ (.A1(\wfg_interconnect_top.stimulus_0[4] ),
    .A2(_02796_),
    .B1(_02798_),
    .B2(\wfg_interconnect_top.stimulus_1[4] ),
    .C1(_02748_),
    .X(_02841_));
 sky130_fd_sc_hd__a32o_1 _10233_ (.A1(_02813_),
    .A2(_02840_),
    .A3(_02841_),
    .B1(_02820_),
    .B2(\wfg_drive_spi_top.wfg_drive_spi.spi_data[4] ),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_1 _10234_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[2] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[4] ),
    .S(\wfg_drive_spi_top.wfg_drive_spi.lsbfirst ),
    .X(_02842_));
 sky130_fd_sc_hd__or2_1 _10235_ (.A(_02729_),
    .B(_02842_),
    .X(_02843_));
 sky130_fd_sc_hd__a221o_1 _10236_ (.A1(\wfg_interconnect_top.stimulus_0[3] ),
    .A2(_02796_),
    .B1(_02798_),
    .B2(\wfg_interconnect_top.stimulus_1[3] ),
    .C1(_02748_),
    .X(_02844_));
 sky130_fd_sc_hd__a32o_1 _10237_ (.A1(_02813_),
    .A2(_02843_),
    .A3(_02844_),
    .B1(_02820_),
    .B2(\wfg_drive_spi_top.wfg_drive_spi.spi_data[3] ),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_1 _10238_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[1] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[3] ),
    .S(\wfg_drive_spi_top.wfg_drive_spi.lsbfirst ),
    .X(_02845_));
 sky130_fd_sc_hd__or2_1 _10239_ (.A(_02729_),
    .B(_02845_),
    .X(_02846_));
 sky130_fd_sc_hd__a221o_1 _10240_ (.A1(\wfg_interconnect_top.stimulus_0[2] ),
    .A2(_02796_),
    .B1(_02798_),
    .B2(\wfg_interconnect_top.stimulus_1[2] ),
    .C1(_02748_),
    .X(_02847_));
 sky130_fd_sc_hd__a32o_1 _10241_ (.A1(_02737_),
    .A2(_02846_),
    .A3(_02847_),
    .B1(_02820_),
    .B2(\wfg_drive_spi_top.wfg_drive_spi.spi_data[2] ),
    .X(_01217_));
 sky130_fd_sc_hd__mux2_1 _10242_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[0] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[2] ),
    .S(\wfg_drive_spi_top.wfg_drive_spi.lsbfirst ),
    .X(_02848_));
 sky130_fd_sc_hd__or2_1 _10243_ (.A(_02729_),
    .B(_02848_),
    .X(_02849_));
 sky130_fd_sc_hd__a221o_1 _10244_ (.A1(\wfg_interconnect_top.stimulus_0[1] ),
    .A2(_02796_),
    .B1(_02798_),
    .B2(\wfg_interconnect_top.stimulus_1[1] ),
    .C1(_02748_),
    .X(_02850_));
 sky130_fd_sc_hd__a32o_1 _10245_ (.A1(_02737_),
    .A2(_02849_),
    .A3(_02850_),
    .B1(_02735_),
    .B2(\wfg_drive_spi_top.wfg_drive_spi.spi_data[1] ),
    .X(_01216_));
 sky130_fd_sc_hd__a221o_1 _10246_ (.A1(\wfg_interconnect_top.stimulus_0[0] ),
    .A2(_02796_),
    .B1(_02798_),
    .B2(\wfg_interconnect_top.stimulus_1[0] ),
    .C1(_02748_),
    .X(_02851_));
 sky130_fd_sc_hd__a21o_1 _10247_ (.A1(_02723_),
    .A2(\wfg_drive_spi_top.wfg_drive_spi.spi_data[1] ),
    .B1(_02793_),
    .X(_02852_));
 sky130_fd_sc_hd__a32o_1 _10248_ (.A1(_02737_),
    .A2(_02851_),
    .A3(_02852_),
    .B1(_02735_),
    .B2(\wfg_drive_spi_top.wfg_drive_spi.spi_data[0] ),
    .X(_01215_));
 sky130_fd_sc_hd__a211o_1 _10249_ (.A1(_02702_),
    .A2(_02800_),
    .B1(_02735_),
    .C1(_02712_),
    .X(_02853_));
 sky130_fd_sc_hd__a22o_1 _10250_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.byte_cnt[1] ),
    .A2(_02711_),
    .B1(_02853_),
    .B2(\wfg_drive_spi_top.wfg_drive_spi.current_bit[4] ),
    .X(_01214_));
 sky130_fd_sc_hd__nor2_1 _10251_ (.A(\wfg_drive_spi_top.wfg_drive_spi.byte_cnt[0] ),
    .B(_02749_),
    .Y(_02854_));
 sky130_fd_sc_hd__a211o_1 _10252_ (.A1(_02701_),
    .A2(_02800_),
    .B1(_02735_),
    .C1(_02712_),
    .X(_02855_));
 sky130_fd_sc_hd__a2bb2o_1 _10253_ (.A1_N(_02853_),
    .A2_N(_02854_),
    .B1(_02855_),
    .B2(\wfg_drive_spi_top.wfg_drive_spi.current_bit[3] ),
    .X(_01213_));
 sky130_fd_sc_hd__or4_1 _10254_ (.A(\wfg_drive_spi_top.wfg_drive_spi.current_bit[1] ),
    .B(\wfg_drive_spi_top.wfg_drive_spi.current_bit[0] ),
    .C(_02712_),
    .D(_02735_),
    .X(_02856_));
 sky130_fd_sc_hd__a21bo_1 _10255_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.current_bit[2] ),
    .A2(_02856_),
    .B1_N(_02855_),
    .X(_01212_));
 sky130_fd_sc_hd__or3_1 _10256_ (.A(\wfg_drive_spi_top.wfg_drive_spi.current_bit[0] ),
    .B(_02712_),
    .C(_02735_),
    .X(_02857_));
 sky130_fd_sc_hd__o21ai_1 _10257_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.current_bit[1] ),
    .A2(\wfg_drive_spi_top.wfg_drive_spi.current_bit[0] ),
    .B1(_02749_),
    .Y(_02858_));
 sky130_fd_sc_hd__a22o_1 _10258_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.current_bit[1] ),
    .A2(_02857_),
    .B1(_02858_),
    .B2(_02777_),
    .X(_01211_));
 sky130_fd_sc_hd__a21bo_1 _10259_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.cur_state[0] ),
    .A2(_02737_),
    .B1_N(\wfg_drive_spi_top.wfg_drive_spi.current_bit[0] ),
    .X(_02859_));
 sky130_fd_sc_hd__nand2_1 _10260_ (.A(_02857_),
    .B(_02859_),
    .Y(_01210_));
 sky130_fd_sc_hd__mux2_1 _10261_ (.A0(\wfg_drive_spi_top.clkcfg_div_q[7] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.clk_div[7] ),
    .S(_02719_),
    .X(_02860_));
 sky130_fd_sc_hd__clkbuf_1 _10262_ (.A(_02860_),
    .X(_01209_));
 sky130_fd_sc_hd__mux2_1 _10263_ (.A0(\wfg_drive_spi_top.clkcfg_div_q[6] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.clk_div[6] ),
    .S(_02719_),
    .X(_02861_));
 sky130_fd_sc_hd__clkbuf_1 _10264_ (.A(_02861_),
    .X(_01208_));
 sky130_fd_sc_hd__mux2_1 _10265_ (.A0(\wfg_drive_spi_top.clkcfg_div_q[5] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.clk_div[5] ),
    .S(_02719_),
    .X(_02862_));
 sky130_fd_sc_hd__clkbuf_1 _10266_ (.A(_02862_),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_1 _10267_ (.A0(\wfg_drive_spi_top.clkcfg_div_q[4] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.clk_div[4] ),
    .S(_02719_),
    .X(_02863_));
 sky130_fd_sc_hd__clkbuf_1 _10268_ (.A(_02863_),
    .X(_01206_));
 sky130_fd_sc_hd__mux2_1 _10269_ (.A0(\wfg_drive_spi_top.clkcfg_div_q[3] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.clk_div[3] ),
    .S(_02719_),
    .X(_02864_));
 sky130_fd_sc_hd__clkbuf_1 _10270_ (.A(_02864_),
    .X(_01205_));
 sky130_fd_sc_hd__mux2_1 _10271_ (.A0(\wfg_drive_spi_top.clkcfg_div_q[2] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.clk_div[2] ),
    .S(_02717_),
    .X(_02865_));
 sky130_fd_sc_hd__clkbuf_1 _10272_ (.A(_02865_),
    .X(_01204_));
 sky130_fd_sc_hd__mux2_1 _10273_ (.A0(\wfg_drive_spi_top.clkcfg_div_q[1] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.clk_div[1] ),
    .S(_02717_),
    .X(_02866_));
 sky130_fd_sc_hd__clkbuf_1 _10274_ (.A(_02866_),
    .X(_01203_));
 sky130_fd_sc_hd__mux2_1 _10275_ (.A0(\wfg_drive_spi_top.clkcfg_div_q[0] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.clk_div[0] ),
    .S(_02717_),
    .X(_02867_));
 sky130_fd_sc_hd__clkbuf_1 _10276_ (.A(_02867_),
    .X(_01202_));
 sky130_fd_sc_hd__o21a_1 _10277_ (.A1(_02727_),
    .A2(_02793_),
    .B1(\wfg_drive_spi_top.wfg_drive_spi.clk_div[7] ),
    .X(_02868_));
 sky130_fd_sc_hd__nor2_1 _10278_ (.A(\wfg_drive_spi_top.wfg_drive_spi.counter[6] ),
    .B(_02699_),
    .Y(_02869_));
 sky130_fd_sc_hd__and3b_1 _10279_ (.A_N(_02869_),
    .B(_02740_),
    .C(\wfg_drive_spi_top.wfg_drive_spi.counter[7] ),
    .X(_02870_));
 sky130_fd_sc_hd__o21a_1 _10280_ (.A1(_02868_),
    .A2(_02870_),
    .B1(_00003_),
    .X(_01201_));
 sky130_fd_sc_hd__o21a_1 _10281_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.clk_div[6] ),
    .A2(\wfg_drive_spi_top.wfg_drive_spi.counter[7] ),
    .B1(_02869_),
    .X(_02871_));
 sky130_fd_sc_hd__a211o_1 _10282_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.counter[6] ),
    .A2(_02699_),
    .B1(_02793_),
    .C1(_02871_),
    .X(_02872_));
 sky130_fd_sc_hd__o211a_1 _10283_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.clk_div[6] ),
    .A2(_02749_),
    .B1(_02872_),
    .C1(_00003_),
    .X(_01200_));
 sky130_fd_sc_hd__o21a_1 _10284_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.counter[4] ),
    .A2(_02698_),
    .B1(\wfg_drive_spi_top.wfg_drive_spi.counter[5] ),
    .X(_02873_));
 sky130_fd_sc_hd__or3b_1 _10285_ (.A(_02793_),
    .B(_02873_),
    .C_N(_02699_),
    .X(_02874_));
 sky130_fd_sc_hd__o211a_1 _10286_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.clk_div[5] ),
    .A2(_02730_),
    .B1(_02874_),
    .C1(_00003_),
    .X(_01199_));
 sky130_fd_sc_hd__nor2_1 _10287_ (.A(\wfg_drive_spi_top.wfg_drive_spi.counter[4] ),
    .B(_02698_),
    .Y(_02875_));
 sky130_fd_sc_hd__and2_1 _10288_ (.A(\wfg_drive_spi_top.wfg_drive_spi.counter[4] ),
    .B(_02698_),
    .X(_02876_));
 sky130_fd_sc_hd__or4_1 _10289_ (.A(\wfg_drive_spi_top.wfg_drive_spi.counter[7] ),
    .B(\wfg_drive_spi_top.wfg_drive_spi.counter[6] ),
    .C(\wfg_drive_spi_top.wfg_drive_spi.counter[5] ),
    .D(\wfg_drive_spi_top.wfg_drive_spi.counter[4] ),
    .X(_02877_));
 sky130_fd_sc_hd__a21o_1 _10290_ (.A1(_02749_),
    .A2(_02877_),
    .B1(\wfg_drive_spi_top.wfg_drive_spi.clk_div[4] ),
    .X(_02878_));
 sky130_fd_sc_hd__o311a_1 _10291_ (.A1(_02875_),
    .A2(_02793_),
    .A3(_02876_),
    .B1(_02878_),
    .C1(_00003_),
    .X(_01198_));
 sky130_fd_sc_hd__o21a_1 _10292_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.counter[2] ),
    .A2(_02697_),
    .B1(\wfg_drive_spi_top.wfg_drive_spi.counter[3] ),
    .X(_02879_));
 sky130_fd_sc_hd__or3b_1 _10293_ (.A(_02793_),
    .B(_02879_),
    .C_N(_02698_),
    .X(_02880_));
 sky130_fd_sc_hd__o211a_1 _10294_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.clk_div[3] ),
    .A2(_02730_),
    .B1(_02880_),
    .C1(_00003_),
    .X(_01197_));
 sky130_fd_sc_hd__nor2_1 _10295_ (.A(\wfg_drive_spi_top.wfg_drive_spi.counter[2] ),
    .B(_02697_),
    .Y(_02881_));
 sky130_fd_sc_hd__a211o_1 _10296_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.counter[2] ),
    .A2(_02697_),
    .B1(_02881_),
    .C1(_02793_),
    .X(_02882_));
 sky130_fd_sc_hd__o211a_1 _10297_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.clk_div[2] ),
    .A2(_02730_),
    .B1(_02882_),
    .C1(_00003_),
    .X(_01196_));
 sky130_fd_sc_hd__nand2_1 _10298_ (.A(\wfg_drive_spi_top.wfg_drive_spi.counter[1] ),
    .B(\wfg_drive_spi_top.wfg_drive_spi.counter[0] ),
    .Y(_02883_));
 sky130_fd_sc_hd__o21ai_1 _10299_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.clk_div[1] ),
    .A2(_02730_),
    .B1(_00003_),
    .Y(_02884_));
 sky130_fd_sc_hd__a31oi_1 _10300_ (.A1(_02697_),
    .A2(_02730_),
    .A3(_02883_),
    .B1(_02884_),
    .Y(_01195_));
 sky130_fd_sc_hd__nand2_1 _10301_ (.A(\wfg_drive_spi_top.wfg_drive_spi.counter[0] ),
    .B(_02730_),
    .Y(_02885_));
 sky130_fd_sc_hd__o211a_1 _10302_ (.A1(\wfg_drive_spi_top.wfg_drive_spi.clk_div[0] ),
    .A2(_02730_),
    .B1(_02885_),
    .C1(_00003_),
    .X(_01194_));
 sky130_fd_sc_hd__clkbuf_4 _10303_ (.A(\wfg_stim_mem_top.cfg_gain_q[8] ),
    .X(_02886_));
 sky130_fd_sc_hd__buf_4 _10304_ (.A(_02886_),
    .X(_02887_));
 sky130_fd_sc_hd__clkbuf_8 _10305_ (.A(net25),
    .X(_02888_));
 sky130_fd_sc_hd__buf_4 _10306_ (.A(_02888_),
    .X(_02889_));
 sky130_fd_sc_hd__and2_1 _10307_ (.A(_02887_),
    .B(_02889_),
    .X(_02890_));
 sky130_fd_sc_hd__buf_2 _10308_ (.A(_02890_),
    .X(_02891_));
 sky130_fd_sc_hd__buf_6 _10309_ (.A(\wfg_stim_mem_top.cfg_gain_q[9] ),
    .X(_02892_));
 sky130_fd_sc_hd__nand2_8 _10310_ (.A(_02892_),
    .B(_02888_),
    .Y(_02893_));
 sky130_fd_sc_hd__clkbuf_4 _10311_ (.A(\wfg_stim_mem_top.cfg_gain_q[13] ),
    .X(_02894_));
 sky130_fd_sc_hd__buf_6 _10312_ (.A(_02894_),
    .X(_02895_));
 sky130_fd_sc_hd__buf_4 _10313_ (.A(\wfg_stim_mem_top.cfg_gain_q[12] ),
    .X(_02896_));
 sky130_fd_sc_hd__buf_8 _10314_ (.A(_02896_),
    .X(_02897_));
 sky130_fd_sc_hd__o21ai_1 _10315_ (.A1(_02895_),
    .A2(_02897_),
    .B1(_02889_),
    .Y(_02898_));
 sky130_fd_sc_hd__clkbuf_4 _10316_ (.A(\wfg_stim_mem_top.cfg_gain_q[12] ),
    .X(_02899_));
 sky130_fd_sc_hd__clkbuf_4 _10317_ (.A(_02899_),
    .X(_02900_));
 sky130_fd_sc_hd__and2_1 _10318_ (.A(_02900_),
    .B(_02888_),
    .X(_02901_));
 sky130_fd_sc_hd__a2bb2o_1 _10319_ (.A1_N(_02893_),
    .A2_N(_02898_),
    .B1(_02895_),
    .B2(_02901_),
    .X(_02902_));
 sky130_fd_sc_hd__nand2_1 _10320_ (.A(_02891_),
    .B(_02902_),
    .Y(_02903_));
 sky130_fd_sc_hd__or2_1 _10321_ (.A(_02891_),
    .B(_02902_),
    .X(_02904_));
 sky130_fd_sc_hd__nand2_2 _10322_ (.A(_02903_),
    .B(_02904_),
    .Y(_02905_));
 sky130_fd_sc_hd__clkbuf_4 _10323_ (.A(\wfg_stim_mem_top.cfg_gain_q[11] ),
    .X(_02906_));
 sky130_fd_sc_hd__clkbuf_4 _10324_ (.A(_02906_),
    .X(_02907_));
 sky130_fd_sc_hd__buf_4 _10325_ (.A(_02907_),
    .X(_02908_));
 sky130_fd_sc_hd__buf_8 _10326_ (.A(_02908_),
    .X(_02909_));
 sky130_fd_sc_hd__buf_4 _10327_ (.A(_02889_),
    .X(_02910_));
 sky130_fd_sc_hd__nand2_4 _10328_ (.A(_02909_),
    .B(_02910_),
    .Y(_02911_));
 sky130_fd_sc_hd__xor2_4 _10329_ (.A(_02905_),
    .B(_02911_),
    .X(_02912_));
 sky130_fd_sc_hd__buf_4 _10330_ (.A(_02912_),
    .X(_02913_));
 sky130_fd_sc_hd__clkbuf_4 _10331_ (.A(_02913_),
    .X(_02914_));
 sky130_fd_sc_hd__a21oi_2 _10332_ (.A1(_02895_),
    .A2(_02901_),
    .B1(_02898_),
    .Y(_02915_));
 sky130_fd_sc_hd__xnor2_4 _10333_ (.A(_02893_),
    .B(_02915_),
    .Y(_02916_));
 sky130_fd_sc_hd__buf_4 _10334_ (.A(\wfg_stim_mem_top.cfg_gain_q[14] ),
    .X(_02917_));
 sky130_fd_sc_hd__buf_8 _10335_ (.A(_02917_),
    .X(_02918_));
 sky130_fd_sc_hd__buf_4 _10336_ (.A(\wfg_stim_mem_top.cfg_gain_q[16] ),
    .X(_02919_));
 sky130_fd_sc_hd__buf_4 _10337_ (.A(_02919_),
    .X(_02920_));
 sky130_fd_sc_hd__buf_8 _10338_ (.A(_02920_),
    .X(_02921_));
 sky130_fd_sc_hd__buf_4 _10339_ (.A(\wfg_stim_mem_top.cfg_gain_q[15] ),
    .X(_02922_));
 sky130_fd_sc_hd__buf_8 _10340_ (.A(_02922_),
    .X(_02923_));
 sky130_fd_sc_hd__and3_1 _10341_ (.A(_02921_),
    .B(_02923_),
    .C(_02888_),
    .X(_02924_));
 sky130_fd_sc_hd__and2_1 _10342_ (.A(_02918_),
    .B(_02924_),
    .X(_02925_));
 sky130_fd_sc_hd__buf_4 _10343_ (.A(\wfg_stim_mem_top.cfg_gain_q[14] ),
    .X(_02926_));
 sky130_fd_sc_hd__buf_4 _10344_ (.A(_02926_),
    .X(_02927_));
 sky130_fd_sc_hd__nand2_2 _10345_ (.A(_02927_),
    .B(_02889_),
    .Y(_02928_));
 sky130_fd_sc_hd__o21ai_1 _10346_ (.A1(_02921_),
    .A2(_02923_),
    .B1(_02889_),
    .Y(_02929_));
 sky130_fd_sc_hd__nand2_1 _10347_ (.A(_02928_),
    .B(_02929_),
    .Y(_02930_));
 sky130_fd_sc_hd__and2b_1 _10348_ (.A_N(_02925_),
    .B(_02930_),
    .X(_02931_));
 sky130_fd_sc_hd__xnor2_4 _10349_ (.A(_02916_),
    .B(_02931_),
    .Y(_02932_));
 sky130_fd_sc_hd__clkbuf_4 _10350_ (.A(_02932_),
    .X(_02933_));
 sky130_fd_sc_hd__buf_4 _10351_ (.A(\wfg_stim_mem_top.cfg_gain_q[17] ),
    .X(_02934_));
 sky130_fd_sc_hd__buf_8 _10352_ (.A(_02934_),
    .X(_02935_));
 sky130_fd_sc_hd__nand2_4 _10353_ (.A(_02935_),
    .B(_02888_),
    .Y(_02936_));
 sky130_fd_sc_hd__clkbuf_4 _10354_ (.A(\wfg_stim_mem_top.cfg_gain_q[18] ),
    .X(_02937_));
 sky130_fd_sc_hd__buf_4 _10355_ (.A(_02937_),
    .X(_02938_));
 sky130_fd_sc_hd__clkbuf_4 _10356_ (.A(_02938_),
    .X(_02939_));
 sky130_fd_sc_hd__clkbuf_4 _10357_ (.A(\wfg_stim_mem_top.cfg_gain_q[18] ),
    .X(_02940_));
 sky130_fd_sc_hd__buf_6 _10358_ (.A(_02940_),
    .X(_02941_));
 sky130_fd_sc_hd__nand2_1 _10359_ (.A(_02941_),
    .B(net25),
    .Y(_02942_));
 sky130_fd_sc_hd__buf_4 _10360_ (.A(\wfg_stim_mem_top.cfg_gain_q[19] ),
    .X(_02943_));
 sky130_fd_sc_hd__buf_6 _10361_ (.A(_02943_),
    .X(_02944_));
 sky130_fd_sc_hd__nand2_1 _10362_ (.A(_02944_),
    .B(net25),
    .Y(_02945_));
 sky130_fd_sc_hd__mux2_4 _10363_ (.A0(_02939_),
    .A1(_02942_),
    .S(_02945_),
    .X(_02946_));
 sky130_fd_sc_hd__xor2_4 _10364_ (.A(_02936_),
    .B(_02946_),
    .X(_02947_));
 sky130_fd_sc_hd__buf_4 _10365_ (.A(\wfg_stim_mem_top.cfg_gain_q[20] ),
    .X(_02948_));
 sky130_fd_sc_hd__buf_6 _10366_ (.A(_02948_),
    .X(_02949_));
 sky130_fd_sc_hd__buf_6 _10367_ (.A(_02949_),
    .X(_02950_));
 sky130_fd_sc_hd__buf_4 _10368_ (.A(net24),
    .X(_02951_));
 sky130_fd_sc_hd__clkbuf_4 _10369_ (.A(_02951_),
    .X(_02952_));
 sky130_fd_sc_hd__buf_6 _10370_ (.A(_02952_),
    .X(_02953_));
 sky130_fd_sc_hd__buf_4 _10371_ (.A(\wfg_stim_mem_top.cfg_gain_q[21] ),
    .X(_02954_));
 sky130_fd_sc_hd__buf_6 _10372_ (.A(_02954_),
    .X(_02955_));
 sky130_fd_sc_hd__clkbuf_4 _10373_ (.A(_02955_),
    .X(_02956_));
 sky130_fd_sc_hd__buf_4 _10374_ (.A(net22),
    .X(_02957_));
 sky130_fd_sc_hd__buf_4 _10375_ (.A(net21),
    .X(_02958_));
 sky130_fd_sc_hd__buf_4 _10376_ (.A(\wfg_stim_mem_top.cfg_gain_q[22] ),
    .X(_02959_));
 sky130_fd_sc_hd__clkbuf_8 _10377_ (.A(_02959_),
    .X(_02960_));
 sky130_fd_sc_hd__clkbuf_4 _10378_ (.A(_02960_),
    .X(_02961_));
 sky130_fd_sc_hd__a22o_1 _10379_ (.A1(_02956_),
    .A2(_02957_),
    .B1(_02958_),
    .B2(_02961_),
    .X(_02962_));
 sky130_fd_sc_hd__buf_4 _10380_ (.A(_02959_),
    .X(_02963_));
 sky130_fd_sc_hd__buf_4 _10381_ (.A(_02963_),
    .X(_02964_));
 sky130_fd_sc_hd__buf_4 _10382_ (.A(_02954_),
    .X(_02965_));
 sky130_fd_sc_hd__buf_4 _10383_ (.A(_02965_),
    .X(_02966_));
 sky130_fd_sc_hd__and4_1 _10384_ (.A(_02964_),
    .B(_02966_),
    .C(_02957_),
    .D(_02958_),
    .X(_02967_));
 sky130_fd_sc_hd__a31o_2 _10385_ (.A1(_02950_),
    .A2(_02953_),
    .A3(_02962_),
    .B1(_02967_),
    .X(_02968_));
 sky130_fd_sc_hd__buf_6 _10386_ (.A(_02944_),
    .X(_02969_));
 sky130_fd_sc_hd__inv_2 _10387_ (.A(_02969_),
    .Y(_02970_));
 sky130_fd_sc_hd__o22ai_4 _10388_ (.A1(_02970_),
    .A2(_02942_),
    .B1(_02946_),
    .B2(_02936_),
    .Y(_02971_));
 sky130_fd_sc_hd__xor2_1 _10389_ (.A(_02947_),
    .B(_02968_),
    .X(_02972_));
 sky130_fd_sc_hd__and2_1 _10390_ (.A(_02971_),
    .B(_02972_),
    .X(_02973_));
 sky130_fd_sc_hd__a21oi_1 _10391_ (.A1(_02947_),
    .A2(_02968_),
    .B1(_02973_),
    .Y(_02974_));
 sky130_fd_sc_hd__a21oi_4 _10392_ (.A1(_02916_),
    .A2(_02930_),
    .B1(_02925_),
    .Y(_02975_));
 sky130_fd_sc_hd__clkbuf_4 _10393_ (.A(_02975_),
    .X(_02976_));
 sky130_fd_sc_hd__xnor2_1 _10394_ (.A(_02933_),
    .B(_02974_),
    .Y(_02977_));
 sky130_fd_sc_hd__or2_1 _10395_ (.A(_02976_),
    .B(_02977_),
    .X(_02978_));
 sky130_fd_sc_hd__o21ai_1 _10396_ (.A1(_02933_),
    .A2(_02974_),
    .B1(_02978_),
    .Y(_02979_));
 sky130_fd_sc_hd__o21ai_2 _10397_ (.A1(_02905_),
    .A2(_02911_),
    .B1(_02903_),
    .Y(_02980_));
 sky130_fd_sc_hd__clkbuf_4 _10398_ (.A(_02980_),
    .X(_02981_));
 sky130_fd_sc_hd__clkbuf_4 _10399_ (.A(_02981_),
    .X(_02982_));
 sky130_fd_sc_hd__xor2_1 _10400_ (.A(_02913_),
    .B(_02979_),
    .X(_02983_));
 sky130_fd_sc_hd__nand2_1 _10401_ (.A(_02982_),
    .B(_02983_),
    .Y(_02984_));
 sky130_fd_sc_hd__a21bo_1 _10402_ (.A1(_02914_),
    .A2(_02979_),
    .B1_N(_02984_),
    .X(_02985_));
 sky130_fd_sc_hd__buf_6 _10403_ (.A(_02966_),
    .X(_02986_));
 sky130_fd_sc_hd__clkbuf_4 _10404_ (.A(_02957_),
    .X(_02987_));
 sky130_fd_sc_hd__buf_6 _10405_ (.A(_02964_),
    .X(_02988_));
 sky130_fd_sc_hd__a22o_1 _10406_ (.A1(_02986_),
    .A2(_02952_),
    .B1(_02987_),
    .B2(_02988_),
    .X(_02989_));
 sky130_fd_sc_hd__and4_1 _10407_ (.A(_02988_),
    .B(_02986_),
    .C(_02951_),
    .D(_02987_),
    .X(_02990_));
 sky130_fd_sc_hd__a31o_1 _10408_ (.A1(_02950_),
    .A2(_02910_),
    .A3(_02989_),
    .B1(_02990_),
    .X(_02991_));
 sky130_fd_sc_hd__xor2_1 _10409_ (.A(_02947_),
    .B(_02991_),
    .X(_02992_));
 sky130_fd_sc_hd__and2_1 _10410_ (.A(_02971_),
    .B(_02992_),
    .X(_02993_));
 sky130_fd_sc_hd__a21oi_1 _10411_ (.A1(_02947_),
    .A2(_02991_),
    .B1(_02993_),
    .Y(_02994_));
 sky130_fd_sc_hd__xnor2_1 _10412_ (.A(_02933_),
    .B(_02994_),
    .Y(_02995_));
 sky130_fd_sc_hd__or2_1 _10413_ (.A(_02976_),
    .B(_02995_),
    .X(_02996_));
 sky130_fd_sc_hd__o21ai_1 _10414_ (.A1(_02933_),
    .A2(_02994_),
    .B1(_02996_),
    .Y(_02997_));
 sky130_fd_sc_hd__xor2_1 _10415_ (.A(_02914_),
    .B(_02997_),
    .X(_02998_));
 sky130_fd_sc_hd__nand2_1 _10416_ (.A(_02982_),
    .B(_02998_),
    .Y(_02999_));
 sky130_fd_sc_hd__or2_1 _10417_ (.A(_02982_),
    .B(_02998_),
    .X(_03000_));
 sky130_fd_sc_hd__and2_1 _10418_ (.A(_02999_),
    .B(_03000_),
    .X(_03001_));
 sky130_fd_sc_hd__and3_1 _10419_ (.A(_02988_),
    .B(_02986_),
    .C(_02889_),
    .X(_03002_));
 sky130_fd_sc_hd__and2_1 _10420_ (.A(_02953_),
    .B(_03002_),
    .X(_03003_));
 sky130_fd_sc_hd__a22o_1 _10421_ (.A1(_02986_),
    .A2(_02889_),
    .B1(_02953_),
    .B2(_02988_),
    .X(_03004_));
 sky130_fd_sc_hd__and2b_1 _10422_ (.A_N(_03003_),
    .B(_03004_),
    .X(_03005_));
 sky130_fd_sc_hd__a31o_1 _10423_ (.A1(_02950_),
    .A2(_02910_),
    .A3(_03005_),
    .B1(_03003_),
    .X(_03006_));
 sky130_fd_sc_hd__xor2_1 _10424_ (.A(_02947_),
    .B(_03006_),
    .X(_03007_));
 sky130_fd_sc_hd__xnor2_1 _10425_ (.A(_02971_),
    .B(_03007_),
    .Y(_03008_));
 sky130_fd_sc_hd__nand2_2 _10426_ (.A(_02950_),
    .B(_02889_),
    .Y(_03009_));
 sky130_fd_sc_hd__or2_1 _10427_ (.A(_02988_),
    .B(_02986_),
    .X(_03010_));
 sky130_fd_sc_hd__and3b_1 _10428_ (.A_N(_03002_),
    .B(_03010_),
    .C(_02910_),
    .X(_03011_));
 sky130_fd_sc_hd__xor2_2 _10429_ (.A(_03009_),
    .B(_03011_),
    .X(_03012_));
 sky130_fd_sc_hd__clkbuf_4 _10430_ (.A(\wfg_stim_mem_top.cfg_gain_q[23] ),
    .X(_03013_));
 sky130_fd_sc_hd__clkbuf_8 _10431_ (.A(_03013_),
    .X(_03014_));
 sky130_fd_sc_hd__buf_6 _10432_ (.A(_03014_),
    .X(_03015_));
 sky130_fd_sc_hd__buf_6 _10433_ (.A(_03015_),
    .X(_03016_));
 sky130_fd_sc_hd__nand2_1 _10434_ (.A(_03016_),
    .B(_02953_),
    .Y(_03017_));
 sky130_fd_sc_hd__clkbuf_4 _10435_ (.A(\wfg_stim_mem_top.cfg_gain_q[10] ),
    .X(_03018_));
 sky130_fd_sc_hd__buf_6 _10436_ (.A(_03018_),
    .X(_03019_));
 sky130_fd_sc_hd__and2_2 _10437_ (.A(_03019_),
    .B(_02888_),
    .X(_03020_));
 sky130_fd_sc_hd__clkbuf_4 _10438_ (.A(_03020_),
    .X(_03021_));
 sky130_fd_sc_hd__buf_6 _10439_ (.A(_02987_),
    .X(_03022_));
 sky130_fd_sc_hd__nand2_1 _10440_ (.A(_03016_),
    .B(_03022_),
    .Y(_03023_));
 sky130_fd_sc_hd__nand2_1 _10441_ (.A(_03021_),
    .B(_03023_),
    .Y(_03024_));
 sky130_fd_sc_hd__xnor2_1 _10442_ (.A(_03017_),
    .B(_03024_),
    .Y(_03025_));
 sky130_fd_sc_hd__nor2_1 _10443_ (.A(_03012_),
    .B(_03025_),
    .Y(_03026_));
 sky130_fd_sc_hd__and2_1 _10444_ (.A(_03012_),
    .B(_03025_),
    .X(_03027_));
 sky130_fd_sc_hd__nor2_1 _10445_ (.A(_03026_),
    .B(_03027_),
    .Y(_03028_));
 sky130_fd_sc_hd__buf_4 _10446_ (.A(_02958_),
    .X(_03029_));
 sky130_fd_sc_hd__nand2_1 _10447_ (.A(_03016_),
    .B(_03029_),
    .Y(_03030_));
 sky130_fd_sc_hd__nand2_1 _10448_ (.A(_03021_),
    .B(_03030_),
    .Y(_03031_));
 sky130_fd_sc_hd__xor2_1 _10449_ (.A(_03023_),
    .B(_03031_),
    .X(_03032_));
 sky130_fd_sc_hd__xnor2_1 _10450_ (.A(_03009_),
    .B(_03005_),
    .Y(_03033_));
 sky130_fd_sc_hd__a2bb2o_1 _10451_ (.A1_N(_03024_),
    .A2_N(_03030_),
    .B1(_03032_),
    .B2(_03033_),
    .X(_03034_));
 sky130_fd_sc_hd__xor2_1 _10452_ (.A(_03028_),
    .B(_03034_),
    .X(_03035_));
 sky130_fd_sc_hd__xor2_1 _10453_ (.A(_03008_),
    .B(_03035_),
    .X(_03036_));
 sky130_fd_sc_hd__xor2_1 _10454_ (.A(_03033_),
    .B(_03032_),
    .X(_03037_));
 sky130_fd_sc_hd__buf_4 _10455_ (.A(net20),
    .X(_03038_));
 sky130_fd_sc_hd__clkbuf_4 _10456_ (.A(_03038_),
    .X(_03039_));
 sky130_fd_sc_hd__buf_4 _10457_ (.A(_03039_),
    .X(_03040_));
 sky130_fd_sc_hd__nand2_1 _10458_ (.A(_03016_),
    .B(_03040_),
    .Y(_03041_));
 sky130_fd_sc_hd__and2b_1 _10459_ (.A_N(_02990_),
    .B(_02989_),
    .X(_03042_));
 sky130_fd_sc_hd__xnor2_1 _10460_ (.A(_03009_),
    .B(_03042_),
    .Y(_03043_));
 sky130_fd_sc_hd__nand2_1 _10461_ (.A(_03021_),
    .B(_03041_),
    .Y(_03044_));
 sky130_fd_sc_hd__xor2_1 _10462_ (.A(_03030_),
    .B(_03044_),
    .X(_03045_));
 sky130_fd_sc_hd__nand2_1 _10463_ (.A(_03043_),
    .B(_03045_),
    .Y(_03046_));
 sky130_fd_sc_hd__o21ai_1 _10464_ (.A1(_03031_),
    .A2(_03041_),
    .B1(_03046_),
    .Y(_03047_));
 sky130_fd_sc_hd__nor2_1 _10465_ (.A(_02971_),
    .B(_02992_),
    .Y(_03048_));
 sky130_fd_sc_hd__nor2_1 _10466_ (.A(_02993_),
    .B(_03048_),
    .Y(_03049_));
 sky130_fd_sc_hd__xor2_1 _10467_ (.A(_03037_),
    .B(_03047_),
    .X(_03050_));
 sky130_fd_sc_hd__and2_1 _10468_ (.A(_03049_),
    .B(_03050_),
    .X(_03051_));
 sky130_fd_sc_hd__a21oi_1 _10469_ (.A1(_03037_),
    .A2(_03047_),
    .B1(_03051_),
    .Y(_03052_));
 sky130_fd_sc_hd__nor2_1 _10470_ (.A(_03036_),
    .B(_03052_),
    .Y(_03053_));
 sky130_fd_sc_hd__nand2_1 _10471_ (.A(_02976_),
    .B(_02995_),
    .Y(_03054_));
 sky130_fd_sc_hd__nand2_1 _10472_ (.A(_02996_),
    .B(_03054_),
    .Y(_03055_));
 sky130_fd_sc_hd__and2_1 _10473_ (.A(_03036_),
    .B(_03052_),
    .X(_03056_));
 sky130_fd_sc_hd__or2_1 _10474_ (.A(_03053_),
    .B(_03056_),
    .X(_03057_));
 sky130_fd_sc_hd__nor2_1 _10475_ (.A(_03055_),
    .B(_03057_),
    .Y(_03058_));
 sky130_fd_sc_hd__and2_1 _10476_ (.A(_02971_),
    .B(_03007_),
    .X(_03059_));
 sky130_fd_sc_hd__a21oi_1 _10477_ (.A1(_02947_),
    .A2(_03006_),
    .B1(_03059_),
    .Y(_03060_));
 sky130_fd_sc_hd__xnor2_1 _10478_ (.A(_02933_),
    .B(_03060_),
    .Y(_03061_));
 sky130_fd_sc_hd__xnor2_1 _10479_ (.A(_02976_),
    .B(_03061_),
    .Y(_03062_));
 sky130_fd_sc_hd__a31o_1 _10480_ (.A1(_02950_),
    .A2(_02910_),
    .A3(_03010_),
    .B1(_03002_),
    .X(_03063_));
 sky130_fd_sc_hd__and2_1 _10481_ (.A(_02947_),
    .B(_03063_),
    .X(_03064_));
 sky130_fd_sc_hd__nor2_1 _10482_ (.A(_02947_),
    .B(_03063_),
    .Y(_03065_));
 sky130_fd_sc_hd__nor2_1 _10483_ (.A(_03064_),
    .B(_03065_),
    .Y(_03066_));
 sky130_fd_sc_hd__xnor2_2 _10484_ (.A(_02971_),
    .B(_03066_),
    .Y(_03067_));
 sky130_fd_sc_hd__a41o_1 _10485_ (.A1(_03016_),
    .A2(_03022_),
    .A3(_03017_),
    .A4(_03021_),
    .B1(_03026_),
    .X(_03068_));
 sky130_fd_sc_hd__buf_6 _10486_ (.A(_03019_),
    .X(_03069_));
 sky130_fd_sc_hd__nand2_1 _10487_ (.A(_03069_),
    .B(_02888_),
    .Y(_03070_));
 sky130_fd_sc_hd__nand2_1 _10488_ (.A(_03016_),
    .B(_02889_),
    .Y(_03071_));
 sky130_fd_sc_hd__and2_2 _10489_ (.A(_03070_),
    .B(_03071_),
    .X(_03072_));
 sky130_fd_sc_hd__a31o_1 _10490_ (.A1(_03016_),
    .A2(_03017_),
    .A3(_03021_),
    .B1(_03072_),
    .X(_03073_));
 sky130_fd_sc_hd__xnor2_1 _10491_ (.A(_03012_),
    .B(_03073_),
    .Y(_03074_));
 sky130_fd_sc_hd__xnor2_1 _10492_ (.A(_03068_),
    .B(_03074_),
    .Y(_03075_));
 sky130_fd_sc_hd__xnor2_1 _10493_ (.A(_03067_),
    .B(_03075_),
    .Y(_03076_));
 sky130_fd_sc_hd__and2b_1 _10494_ (.A_N(_03008_),
    .B(_03035_),
    .X(_03077_));
 sky130_fd_sc_hd__a21oi_1 _10495_ (.A1(_03028_),
    .A2(_03034_),
    .B1(_03077_),
    .Y(_03078_));
 sky130_fd_sc_hd__xor2_1 _10496_ (.A(_03076_),
    .B(_03078_),
    .X(_03079_));
 sky130_fd_sc_hd__nor2_1 _10497_ (.A(_03062_),
    .B(_03079_),
    .Y(_03080_));
 sky130_fd_sc_hd__and2_1 _10498_ (.A(_03062_),
    .B(_03079_),
    .X(_03081_));
 sky130_fd_sc_hd__nor2_1 _10499_ (.A(_03080_),
    .B(_03081_),
    .Y(_03082_));
 sky130_fd_sc_hd__o21a_1 _10500_ (.A1(_03053_),
    .A2(_03058_),
    .B1(_03082_),
    .X(_03083_));
 sky130_fd_sc_hd__nor3_1 _10501_ (.A(_03082_),
    .B(_03053_),
    .C(_03058_),
    .Y(_03084_));
 sky130_fd_sc_hd__nor2_1 _10502_ (.A(_03083_),
    .B(_03084_),
    .Y(_03085_));
 sky130_fd_sc_hd__xnor2_1 _10503_ (.A(_03001_),
    .B(_03085_),
    .Y(_03086_));
 sky130_fd_sc_hd__or2_1 _10504_ (.A(_02982_),
    .B(_02983_),
    .X(_03087_));
 sky130_fd_sc_hd__and2_1 _10505_ (.A(_02984_),
    .B(_03087_),
    .X(_03088_));
 sky130_fd_sc_hd__and2_1 _10506_ (.A(_03055_),
    .B(_03057_),
    .X(_03089_));
 sky130_fd_sc_hd__nor2_1 _10507_ (.A(_03058_),
    .B(_03089_),
    .Y(_03090_));
 sky130_fd_sc_hd__or2_1 _10508_ (.A(_03043_),
    .B(_03045_),
    .X(_03091_));
 sky130_fd_sc_hd__and2_1 _10509_ (.A(_03046_),
    .B(_03091_),
    .X(_03092_));
 sky130_fd_sc_hd__buf_4 _10510_ (.A(net19),
    .X(_03093_));
 sky130_fd_sc_hd__clkbuf_4 _10511_ (.A(_03093_),
    .X(_03094_));
 sky130_fd_sc_hd__buf_4 _10512_ (.A(_03094_),
    .X(_03095_));
 sky130_fd_sc_hd__nand2_1 _10513_ (.A(_03015_),
    .B(_03095_),
    .Y(_03096_));
 sky130_fd_sc_hd__nand2_1 _10514_ (.A(_03021_),
    .B(_03096_),
    .Y(_03097_));
 sky130_fd_sc_hd__xor2_1 _10515_ (.A(_03041_),
    .B(_03097_),
    .X(_03098_));
 sky130_fd_sc_hd__and2b_1 _10516_ (.A_N(_02967_),
    .B(_02962_),
    .X(_03099_));
 sky130_fd_sc_hd__buf_4 _10517_ (.A(_02949_),
    .X(_03100_));
 sky130_fd_sc_hd__nand2_1 _10518_ (.A(_03100_),
    .B(_02952_),
    .Y(_03101_));
 sky130_fd_sc_hd__xnor2_2 _10519_ (.A(_03099_),
    .B(_03101_),
    .Y(_03102_));
 sky130_fd_sc_hd__a2bb2o_1 _10520_ (.A1_N(_03044_),
    .A2_N(_03096_),
    .B1(_03098_),
    .B2(_03102_),
    .X(_03103_));
 sky130_fd_sc_hd__nand2_1 _10521_ (.A(_03092_),
    .B(_03103_),
    .Y(_03104_));
 sky130_fd_sc_hd__nor2_1 _10522_ (.A(_02971_),
    .B(_02972_),
    .Y(_03105_));
 sky130_fd_sc_hd__nor2_1 _10523_ (.A(_02973_),
    .B(_03105_),
    .Y(_03106_));
 sky130_fd_sc_hd__xor2_1 _10524_ (.A(_03092_),
    .B(_03103_),
    .X(_03107_));
 sky130_fd_sc_hd__nand2_1 _10525_ (.A(_03106_),
    .B(_03107_),
    .Y(_03108_));
 sky130_fd_sc_hd__nor2_1 _10526_ (.A(_03049_),
    .B(_03050_),
    .Y(_03109_));
 sky130_fd_sc_hd__or2_1 _10527_ (.A(_03051_),
    .B(_03109_),
    .X(_03110_));
 sky130_fd_sc_hd__a21oi_1 _10528_ (.A1(_03104_),
    .A2(_03108_),
    .B1(_03110_),
    .Y(_03111_));
 sky130_fd_sc_hd__nand2_1 _10529_ (.A(_02976_),
    .B(_02977_),
    .Y(_03112_));
 sky130_fd_sc_hd__nand2_1 _10530_ (.A(_02978_),
    .B(_03112_),
    .Y(_03113_));
 sky130_fd_sc_hd__and3_1 _10531_ (.A(_03110_),
    .B(_03104_),
    .C(_03108_),
    .X(_03114_));
 sky130_fd_sc_hd__nor3_1 _10532_ (.A(_03111_),
    .B(_03113_),
    .C(_03114_),
    .Y(_03115_));
 sky130_fd_sc_hd__nor2_1 _10533_ (.A(_03111_),
    .B(_03115_),
    .Y(_03116_));
 sky130_fd_sc_hd__xnor2_1 _10534_ (.A(_03090_),
    .B(_03116_),
    .Y(_03117_));
 sky130_fd_sc_hd__and2b_1 _10535_ (.A_N(_03116_),
    .B(_03090_),
    .X(_03118_));
 sky130_fd_sc_hd__a21oi_1 _10536_ (.A1(_03088_),
    .A2(_03117_),
    .B1(_03118_),
    .Y(_03119_));
 sky130_fd_sc_hd__nor2_1 _10537_ (.A(_03086_),
    .B(_03119_),
    .Y(_03120_));
 sky130_fd_sc_hd__and2_1 _10538_ (.A(_03086_),
    .B(_03119_),
    .X(_03121_));
 sky130_fd_sc_hd__nor2_1 _10539_ (.A(_03120_),
    .B(_03121_),
    .Y(_03122_));
 sky130_fd_sc_hd__xnor2_1 _10540_ (.A(_02985_),
    .B(_03122_),
    .Y(_03123_));
 sky130_fd_sc_hd__xor2_1 _10541_ (.A(_03088_),
    .B(_03117_),
    .X(_03124_));
 sky130_fd_sc_hd__inv_2 _10542_ (.A(_03124_),
    .Y(_03125_));
 sky130_fd_sc_hd__xor2_1 _10543_ (.A(_03102_),
    .B(_03098_),
    .X(_03126_));
 sky130_fd_sc_hd__buf_4 _10544_ (.A(net18),
    .X(_03127_));
 sky130_fd_sc_hd__clkbuf_4 _10545_ (.A(_03127_),
    .X(_03128_));
 sky130_fd_sc_hd__buf_4 _10546_ (.A(_03128_),
    .X(_03129_));
 sky130_fd_sc_hd__nand2_1 _10547_ (.A(_03015_),
    .B(_03129_),
    .Y(_03130_));
 sky130_fd_sc_hd__nand2_1 _10548_ (.A(_03021_),
    .B(_03130_),
    .Y(_03131_));
 sky130_fd_sc_hd__xor2_1 _10549_ (.A(_03096_),
    .B(_03131_),
    .X(_03132_));
 sky130_fd_sc_hd__and4_1 _10550_ (.A(_02964_),
    .B(_02966_),
    .C(_02958_),
    .D(_03038_),
    .X(_03133_));
 sky130_fd_sc_hd__a22o_1 _10551_ (.A1(_02966_),
    .A2(_02958_),
    .B1(_03038_),
    .B2(_02964_),
    .X(_03134_));
 sky130_fd_sc_hd__and2b_1 _10552_ (.A_N(_03133_),
    .B(_03134_),
    .X(_03135_));
 sky130_fd_sc_hd__nand2_1 _10553_ (.A(_03100_),
    .B(_02987_),
    .Y(_03136_));
 sky130_fd_sc_hd__xnor2_2 _10554_ (.A(_03135_),
    .B(_03136_),
    .Y(_03137_));
 sky130_fd_sc_hd__a2bb2o_1 _10555_ (.A1_N(_03097_),
    .A2_N(_03130_),
    .B1(_03132_),
    .B2(_03137_),
    .X(_03138_));
 sky130_fd_sc_hd__nand2_1 _10556_ (.A(_03126_),
    .B(_03138_),
    .Y(_03139_));
 sky130_fd_sc_hd__a31o_2 _10557_ (.A1(_03100_),
    .A2(_03022_),
    .A3(_03134_),
    .B1(_03133_),
    .X(_03140_));
 sky130_fd_sc_hd__xor2_1 _10558_ (.A(_02947_),
    .B(_03140_),
    .X(_03141_));
 sky130_fd_sc_hd__buf_8 _10559_ (.A(_02935_),
    .X(_03142_));
 sky130_fd_sc_hd__clkbuf_4 _10560_ (.A(\wfg_stim_mem_top.cfg_gain_q[19] ),
    .X(_03143_));
 sky130_fd_sc_hd__buf_4 _10561_ (.A(_03143_),
    .X(_03144_));
 sky130_fd_sc_hd__clkbuf_4 _10562_ (.A(_03144_),
    .X(_03145_));
 sky130_fd_sc_hd__a22o_1 _10563_ (.A1(_02941_),
    .A2(_02888_),
    .B1(_02951_),
    .B2(_03145_),
    .X(_03146_));
 sky130_fd_sc_hd__and4_1 _10564_ (.A(_03145_),
    .B(_02941_),
    .C(_02888_),
    .D(_02951_),
    .X(_03147_));
 sky130_fd_sc_hd__a31o_1 _10565_ (.A1(_03142_),
    .A2(_02910_),
    .A3(_03146_),
    .B1(_03147_),
    .X(_03148_));
 sky130_fd_sc_hd__xor2_1 _10566_ (.A(_03141_),
    .B(_03148_),
    .X(_03149_));
 sky130_fd_sc_hd__xor2_1 _10567_ (.A(_03126_),
    .B(_03138_),
    .X(_03150_));
 sky130_fd_sc_hd__nand2_1 _10568_ (.A(_03149_),
    .B(_03150_),
    .Y(_03151_));
 sky130_fd_sc_hd__or2_1 _10569_ (.A(_03106_),
    .B(_03107_),
    .X(_03152_));
 sky130_fd_sc_hd__nand2_1 _10570_ (.A(_03108_),
    .B(_03152_),
    .Y(_03153_));
 sky130_fd_sc_hd__a21oi_1 _10571_ (.A1(_03139_),
    .A2(_03151_),
    .B1(_03153_),
    .Y(_03154_));
 sky130_fd_sc_hd__inv_2 _10572_ (.A(_03154_),
    .Y(_03155_));
 sky130_fd_sc_hd__and2_1 _10573_ (.A(_02947_),
    .B(_03140_),
    .X(_03156_));
 sky130_fd_sc_hd__a21oi_1 _10574_ (.A1(_03141_),
    .A2(_03148_),
    .B1(_03156_),
    .Y(_03157_));
 sky130_fd_sc_hd__xnor2_1 _10575_ (.A(_02933_),
    .B(_03157_),
    .Y(_03158_));
 sky130_fd_sc_hd__or2_1 _10576_ (.A(_02975_),
    .B(_03158_),
    .X(_03159_));
 sky130_fd_sc_hd__nand2_1 _10577_ (.A(_02976_),
    .B(_03158_),
    .Y(_03160_));
 sky130_fd_sc_hd__nand2_1 _10578_ (.A(_03159_),
    .B(_03160_),
    .Y(_03161_));
 sky130_fd_sc_hd__and3_1 _10579_ (.A(_03153_),
    .B(_03139_),
    .C(_03151_),
    .X(_03162_));
 sky130_fd_sc_hd__or3_1 _10580_ (.A(_03154_),
    .B(_03161_),
    .C(_03162_),
    .X(_03163_));
 sky130_fd_sc_hd__o21a_1 _10581_ (.A1(_03111_),
    .A2(_03114_),
    .B1(_03113_),
    .X(_03164_));
 sky130_fd_sc_hd__a211oi_1 _10582_ (.A1(_03155_),
    .A2(_03163_),
    .B1(_03115_),
    .C1(_03164_),
    .Y(_03165_));
 sky130_fd_sc_hd__o21ai_1 _10583_ (.A1(_02933_),
    .A2(_03157_),
    .B1(_03159_),
    .Y(_03166_));
 sky130_fd_sc_hd__xor2_1 _10584_ (.A(_02913_),
    .B(_03166_),
    .X(_03167_));
 sky130_fd_sc_hd__nand2_1 _10585_ (.A(_02981_),
    .B(_03167_),
    .Y(_03168_));
 sky130_fd_sc_hd__or2_1 _10586_ (.A(_02981_),
    .B(_03167_),
    .X(_03169_));
 sky130_fd_sc_hd__nand2_1 _10587_ (.A(_03168_),
    .B(_03169_),
    .Y(_03170_));
 sky130_fd_sc_hd__o211a_1 _10588_ (.A1(_03115_),
    .A2(_03164_),
    .B1(_03155_),
    .C1(_03163_),
    .X(_03171_));
 sky130_fd_sc_hd__or3_1 _10589_ (.A(_03165_),
    .B(_03170_),
    .C(_03171_),
    .X(_03172_));
 sky130_fd_sc_hd__and2b_1 _10590_ (.A_N(_03165_),
    .B(_03172_),
    .X(_03173_));
 sky130_fd_sc_hd__xor2_1 _10591_ (.A(_03124_),
    .B(_03173_),
    .X(_03174_));
 sky130_fd_sc_hd__a21bo_1 _10592_ (.A1(_02914_),
    .A2(_03166_),
    .B1_N(_03168_),
    .X(_03175_));
 sky130_fd_sc_hd__or2b_1 _10593_ (.A(_03174_),
    .B_N(_03175_),
    .X(_03176_));
 sky130_fd_sc_hd__o21a_1 _10594_ (.A1(_03125_),
    .A2(_03173_),
    .B1(_03176_),
    .X(_03177_));
 sky130_fd_sc_hd__xnor2_1 _10595_ (.A(_03123_),
    .B(_03177_),
    .Y(_03178_));
 sky130_fd_sc_hd__a21bo_1 _10596_ (.A1(_02914_),
    .A2(_02997_),
    .B1_N(_02999_),
    .X(_03179_));
 sky130_fd_sc_hd__and2b_1 _10597_ (.A_N(_03078_),
    .B(_03076_),
    .X(_03180_));
 sky130_fd_sc_hd__a21oi_1 _10598_ (.A1(_02971_),
    .A2(_03066_),
    .B1(_03064_),
    .Y(_03181_));
 sky130_fd_sc_hd__xnor2_2 _10599_ (.A(_02933_),
    .B(_03181_),
    .Y(_03182_));
 sky130_fd_sc_hd__xnor2_2 _10600_ (.A(_02976_),
    .B(_03182_),
    .Y(_03183_));
 sky130_fd_sc_hd__and2_1 _10601_ (.A(_03012_),
    .B(_03072_),
    .X(_03184_));
 sky130_fd_sc_hd__nand2_1 _10602_ (.A(_03067_),
    .B(_03184_),
    .Y(_03185_));
 sky130_fd_sc_hd__or3_1 _10603_ (.A(_03067_),
    .B(_03075_),
    .C(_03184_),
    .X(_03186_));
 sky130_fd_sc_hd__and2_1 _10604_ (.A(_03185_),
    .B(_03186_),
    .X(_03187_));
 sky130_fd_sc_hd__xnor2_1 _10605_ (.A(_03183_),
    .B(_03187_),
    .Y(_03188_));
 sky130_fd_sc_hd__o21a_1 _10606_ (.A1(_03180_),
    .A2(_03080_),
    .B1(_03188_),
    .X(_03189_));
 sky130_fd_sc_hd__nor3_1 _10607_ (.A(_03180_),
    .B(_03080_),
    .C(_03188_),
    .Y(_03190_));
 sky130_fd_sc_hd__nor2_1 _10608_ (.A(_03189_),
    .B(_03190_),
    .Y(_03191_));
 sky130_fd_sc_hd__or2_1 _10609_ (.A(_02933_),
    .B(_03060_),
    .X(_03192_));
 sky130_fd_sc_hd__or2_1 _10610_ (.A(_02976_),
    .B(_03061_),
    .X(_03193_));
 sky130_fd_sc_hd__nand3_1 _10611_ (.A(_02914_),
    .B(_03192_),
    .C(_03193_),
    .Y(_03194_));
 sky130_fd_sc_hd__a21o_1 _10612_ (.A1(_03192_),
    .A2(_03193_),
    .B1(_02914_),
    .X(_03195_));
 sky130_fd_sc_hd__nand2_1 _10613_ (.A(_03194_),
    .B(_03195_),
    .Y(_03196_));
 sky130_fd_sc_hd__xnor2_1 _10614_ (.A(_02982_),
    .B(_03196_),
    .Y(_03197_));
 sky130_fd_sc_hd__xor2_1 _10615_ (.A(_03191_),
    .B(_03197_),
    .X(_03198_));
 sky130_fd_sc_hd__a21oi_1 _10616_ (.A1(_03001_),
    .A2(_03085_),
    .B1(_03083_),
    .Y(_03199_));
 sky130_fd_sc_hd__nor2_1 _10617_ (.A(_03198_),
    .B(_03199_),
    .Y(_03200_));
 sky130_fd_sc_hd__and2_1 _10618_ (.A(_03198_),
    .B(_03199_),
    .X(_03201_));
 sky130_fd_sc_hd__nor2_1 _10619_ (.A(_03200_),
    .B(_03201_),
    .Y(_03202_));
 sky130_fd_sc_hd__xnor2_2 _10620_ (.A(_03179_),
    .B(_03202_),
    .Y(_03203_));
 sky130_fd_sc_hd__a21oi_1 _10621_ (.A1(_02985_),
    .A2(_03122_),
    .B1(_03120_),
    .Y(_03204_));
 sky130_fd_sc_hd__xor2_1 _10622_ (.A(_03203_),
    .B(_03204_),
    .X(_03205_));
 sky130_fd_sc_hd__and2b_1 _10623_ (.A_N(_03178_),
    .B(_03205_),
    .X(_03206_));
 sky130_fd_sc_hd__inv_2 _10624_ (.A(_03206_),
    .Y(_03207_));
 sky130_fd_sc_hd__buf_4 _10625_ (.A(_02919_),
    .X(_03208_));
 sky130_fd_sc_hd__clkbuf_4 _10626_ (.A(\wfg_stim_mem_top.cfg_gain_q[15] ),
    .X(_03209_));
 sky130_fd_sc_hd__buf_4 _10627_ (.A(_03209_),
    .X(_03210_));
 sky130_fd_sc_hd__and4_2 _10628_ (.A(_03208_),
    .B(_03210_),
    .C(net24),
    .D(_02957_),
    .X(_03211_));
 sky130_fd_sc_hd__buf_4 _10629_ (.A(\wfg_stim_mem_top.cfg_gain_q[15] ),
    .X(_03212_));
 sky130_fd_sc_hd__buf_4 _10630_ (.A(_03212_),
    .X(_03213_));
 sky130_fd_sc_hd__a22o_2 _10631_ (.A1(_03213_),
    .A2(_02951_),
    .B1(_02957_),
    .B2(_03208_),
    .X(_03214_));
 sky130_fd_sc_hd__and2b_1 _10632_ (.A_N(_03211_),
    .B(_03214_),
    .X(_03215_));
 sky130_fd_sc_hd__xnor2_1 _10633_ (.A(_02928_),
    .B(_03215_),
    .Y(_03216_));
 sky130_fd_sc_hd__buf_4 _10634_ (.A(\wfg_stim_mem_top.cfg_gain_q[16] ),
    .X(_03217_));
 sky130_fd_sc_hd__clkbuf_8 _10635_ (.A(_03217_),
    .X(_03218_));
 sky130_fd_sc_hd__and4_1 _10636_ (.A(_03218_),
    .B(_03213_),
    .C(_02957_),
    .D(_02958_),
    .X(_03219_));
 sky130_fd_sc_hd__clkbuf_4 _10637_ (.A(_02958_),
    .X(_03220_));
 sky130_fd_sc_hd__a22oi_1 _10638_ (.A1(_02923_),
    .A2(_02957_),
    .B1(_03220_),
    .B2(_02921_),
    .Y(_03221_));
 sky130_fd_sc_hd__and4bb_1 _10639_ (.A_N(_03219_),
    .B_N(_03221_),
    .C(_02927_),
    .D(_02951_),
    .X(_03222_));
 sky130_fd_sc_hd__nor2_1 _10640_ (.A(_03219_),
    .B(_03222_),
    .Y(_03223_));
 sky130_fd_sc_hd__xnor2_1 _10641_ (.A(_03216_),
    .B(_03223_),
    .Y(_03224_));
 sky130_fd_sc_hd__nand2_1 _10642_ (.A(_02916_),
    .B(_03224_),
    .Y(_03225_));
 sky130_fd_sc_hd__or2_1 _10643_ (.A(_02916_),
    .B(_03224_),
    .X(_03226_));
 sky130_fd_sc_hd__nand2_1 _10644_ (.A(_03225_),
    .B(_03226_),
    .Y(_03227_));
 sky130_fd_sc_hd__buf_4 _10645_ (.A(net15),
    .X(_03228_));
 sky130_fd_sc_hd__buf_4 _10646_ (.A(_03228_),
    .X(_03229_));
 sky130_fd_sc_hd__buf_4 _10647_ (.A(net14),
    .X(_03230_));
 sky130_fd_sc_hd__buf_4 _10648_ (.A(_03230_),
    .X(_03231_));
 sky130_fd_sc_hd__a22oi_1 _10649_ (.A1(_02956_),
    .A2(_03229_),
    .B1(_03231_),
    .B2(_02961_),
    .Y(_03232_));
 sky130_fd_sc_hd__buf_4 _10650_ (.A(net16),
    .X(_03233_));
 sky130_fd_sc_hd__buf_4 _10651_ (.A(_03233_),
    .X(_03234_));
 sky130_fd_sc_hd__nand2_1 _10652_ (.A(_02949_),
    .B(_03234_),
    .Y(_03235_));
 sky130_fd_sc_hd__buf_4 _10653_ (.A(_03230_),
    .X(_03236_));
 sky130_fd_sc_hd__and4_1 _10654_ (.A(_02961_),
    .B(_02956_),
    .C(_03229_),
    .D(_03236_),
    .X(_03237_));
 sky130_fd_sc_hd__o21ba_1 _10655_ (.A1(_03232_),
    .A2(_03235_),
    .B1_N(_03237_),
    .X(_03238_));
 sky130_fd_sc_hd__buf_4 _10656_ (.A(_02934_),
    .X(_03239_));
 sky130_fd_sc_hd__nand2_1 _10657_ (.A(_03239_),
    .B(_03039_),
    .Y(_03240_));
 sky130_fd_sc_hd__and4_1 _10658_ (.A(_02944_),
    .B(_02941_),
    .C(_03093_),
    .D(_03128_),
    .X(_03241_));
 sky130_fd_sc_hd__a22oi_1 _10659_ (.A1(_02939_),
    .A2(_03094_),
    .B1(_03128_),
    .B2(_03145_),
    .Y(_03242_));
 sky130_fd_sc_hd__nor2_1 _10660_ (.A(_03241_),
    .B(_03242_),
    .Y(_03243_));
 sky130_fd_sc_hd__xnor2_1 _10661_ (.A(_03240_),
    .B(_03243_),
    .Y(_03244_));
 sky130_fd_sc_hd__or2b_1 _10662_ (.A(_03238_),
    .B_N(_03244_),
    .X(_03245_));
 sky130_fd_sc_hd__nand2_1 _10663_ (.A(_03239_),
    .B(_03095_),
    .Y(_03246_));
 sky130_fd_sc_hd__buf_4 _10664_ (.A(net17),
    .X(_03247_));
 sky130_fd_sc_hd__buf_4 _10665_ (.A(_03247_),
    .X(_03248_));
 sky130_fd_sc_hd__a22oi_1 _10666_ (.A1(_02939_),
    .A2(_03128_),
    .B1(_03248_),
    .B2(_03145_),
    .Y(_03249_));
 sky130_fd_sc_hd__and4_1 _10667_ (.A(_02944_),
    .B(_02941_),
    .C(_03128_),
    .D(_03248_),
    .X(_03250_));
 sky130_fd_sc_hd__o21ba_1 _10668_ (.A1(_03246_),
    .A2(_03249_),
    .B1_N(_03250_),
    .X(_03251_));
 sky130_fd_sc_hd__xnor2_1 _10669_ (.A(_03238_),
    .B(_03244_),
    .Y(_03252_));
 sky130_fd_sc_hd__or2b_1 _10670_ (.A(_03251_),
    .B_N(_03252_),
    .X(_03253_));
 sky130_fd_sc_hd__nand2_1 _10671_ (.A(_03245_),
    .B(_03253_),
    .Y(_03254_));
 sky130_fd_sc_hd__or2b_1 _10672_ (.A(_03227_),
    .B_N(_03254_),
    .X(_03255_));
 sky130_fd_sc_hd__and4_1 _10673_ (.A(_03218_),
    .B(_03213_),
    .C(_02958_),
    .D(_03038_),
    .X(_03256_));
 sky130_fd_sc_hd__a22oi_1 _10674_ (.A1(_02923_),
    .A2(_03220_),
    .B1(_03039_),
    .B2(_02921_),
    .Y(_03257_));
 sky130_fd_sc_hd__and4bb_1 _10675_ (.A_N(_03256_),
    .B_N(_03257_),
    .C(_02927_),
    .D(_02987_),
    .X(_03258_));
 sky130_fd_sc_hd__nor2_1 _10676_ (.A(_03256_),
    .B(_03258_),
    .Y(_03259_));
 sky130_fd_sc_hd__o2bb2a_1 _10677_ (.A1_N(_02918_),
    .A2_N(_02952_),
    .B1(_03219_),
    .B2(_03221_),
    .X(_03260_));
 sky130_fd_sc_hd__nor2_1 _10678_ (.A(_03222_),
    .B(_03260_),
    .Y(_03261_));
 sky130_fd_sc_hd__and2b_1 _10679_ (.A_N(_03259_),
    .B(_03261_),
    .X(_03262_));
 sky130_fd_sc_hd__xnor2_1 _10680_ (.A(_03261_),
    .B(_03259_),
    .Y(_03263_));
 sky130_fd_sc_hd__and2_1 _10681_ (.A(_02916_),
    .B(_03263_),
    .X(_03264_));
 sky130_fd_sc_hd__xnor2_1 _10682_ (.A(_03254_),
    .B(_03227_),
    .Y(_03265_));
 sky130_fd_sc_hd__o21ai_1 _10683_ (.A1(_03262_),
    .A2(_03264_),
    .B1(_03265_),
    .Y(_03266_));
 sky130_fd_sc_hd__nand2_1 _10684_ (.A(_03255_),
    .B(_03266_),
    .Y(_03267_));
 sky130_fd_sc_hd__nand2_1 _10685_ (.A(_02914_),
    .B(_03267_),
    .Y(_03268_));
 sky130_fd_sc_hd__xor2_1 _10686_ (.A(_02912_),
    .B(_03267_),
    .X(_03269_));
 sky130_fd_sc_hd__nand2_1 _10687_ (.A(_02982_),
    .B(_03269_),
    .Y(_03270_));
 sky130_fd_sc_hd__buf_4 _10688_ (.A(_03233_),
    .X(_03271_));
 sky130_fd_sc_hd__and4_1 _10689_ (.A(_02964_),
    .B(_02966_),
    .C(_03271_),
    .D(_03228_),
    .X(_03272_));
 sky130_fd_sc_hd__a22oi_1 _10690_ (.A1(_02956_),
    .A2(_03271_),
    .B1(_03229_),
    .B2(_02961_),
    .Y(_03273_));
 sky130_fd_sc_hd__buf_4 _10691_ (.A(_03247_),
    .X(_03274_));
 sky130_fd_sc_hd__and4bb_1 _10692_ (.A_N(_03272_),
    .B_N(_03273_),
    .C(_02949_),
    .D(_03274_),
    .X(_03275_));
 sky130_fd_sc_hd__o2bb2a_1 _10693_ (.A1_N(_02949_),
    .A2_N(_03274_),
    .B1(_03272_),
    .B2(_03273_),
    .X(_03276_));
 sky130_fd_sc_hd__nor2_1 _10694_ (.A(_03275_),
    .B(_03276_),
    .Y(_03277_));
 sky130_fd_sc_hd__nand2_1 _10695_ (.A(_03015_),
    .B(_03231_),
    .Y(_03278_));
 sky130_fd_sc_hd__buf_4 _10696_ (.A(net13),
    .X(_03279_));
 sky130_fd_sc_hd__buf_4 _10697_ (.A(_03279_),
    .X(_03280_));
 sky130_fd_sc_hd__buf_6 _10698_ (.A(_03280_),
    .X(_03281_));
 sky130_fd_sc_hd__nand2_2 _10699_ (.A(_03015_),
    .B(_03281_),
    .Y(_03282_));
 sky130_fd_sc_hd__nand2_1 _10700_ (.A(_03020_),
    .B(_03282_),
    .Y(_03283_));
 sky130_fd_sc_hd__xor2_1 _10701_ (.A(_03278_),
    .B(_03283_),
    .X(_03284_));
 sky130_fd_sc_hd__xor2_1 _10702_ (.A(_03277_),
    .B(_03284_),
    .X(_03285_));
 sky130_fd_sc_hd__buf_4 _10703_ (.A(net11),
    .X(_03286_));
 sky130_fd_sc_hd__buf_4 _10704_ (.A(_03286_),
    .X(_03287_));
 sky130_fd_sc_hd__buf_4 _10705_ (.A(_03287_),
    .X(_03288_));
 sky130_fd_sc_hd__nand2_1 _10706_ (.A(_03015_),
    .B(_03288_),
    .Y(_03289_));
 sky130_fd_sc_hd__nand2_1 _10707_ (.A(_03020_),
    .B(_03289_),
    .Y(_03290_));
 sky130_fd_sc_hd__xor2_1 _10708_ (.A(_03282_),
    .B(_03290_),
    .X(_03291_));
 sky130_fd_sc_hd__nor2_1 _10709_ (.A(_03232_),
    .B(_03237_),
    .Y(_03292_));
 sky130_fd_sc_hd__xnor2_1 _10710_ (.A(_03292_),
    .B(_03235_),
    .Y(_03293_));
 sky130_fd_sc_hd__a2bb2o_1 _10711_ (.A1_N(_03283_),
    .A2_N(_03289_),
    .B1(_03291_),
    .B2(_03293_),
    .X(_03294_));
 sky130_fd_sc_hd__nand2_1 _10712_ (.A(_03285_),
    .B(_03294_),
    .Y(_03295_));
 sky130_fd_sc_hd__xnor2_1 _10713_ (.A(_03252_),
    .B(_03251_),
    .Y(_03296_));
 sky130_fd_sc_hd__xor2_1 _10714_ (.A(_03285_),
    .B(_03294_),
    .X(_03297_));
 sky130_fd_sc_hd__nand2_1 _10715_ (.A(_03296_),
    .B(_03297_),
    .Y(_03298_));
 sky130_fd_sc_hd__nor2_1 _10716_ (.A(_03272_),
    .B(_03275_),
    .Y(_03299_));
 sky130_fd_sc_hd__nand2_1 _10717_ (.A(_03142_),
    .B(_03029_),
    .Y(_03300_));
 sky130_fd_sc_hd__and4_1 _10718_ (.A(_02969_),
    .B(_02939_),
    .C(_03039_),
    .D(_03094_),
    .X(_03301_));
 sky130_fd_sc_hd__buf_6 _10719_ (.A(_02941_),
    .X(_03302_));
 sky130_fd_sc_hd__a22oi_1 _10720_ (.A1(_03302_),
    .A2(_03039_),
    .B1(_03095_),
    .B2(_02969_),
    .Y(_03303_));
 sky130_fd_sc_hd__nor2_1 _10721_ (.A(_03301_),
    .B(_03303_),
    .Y(_03304_));
 sky130_fd_sc_hd__xnor2_1 _10722_ (.A(_03300_),
    .B(_03304_),
    .Y(_03305_));
 sky130_fd_sc_hd__xnor2_1 _10723_ (.A(_03299_),
    .B(_03305_),
    .Y(_03306_));
 sky130_fd_sc_hd__o21ba_1 _10724_ (.A1(_03240_),
    .A2(_03242_),
    .B1_N(_03241_),
    .X(_03307_));
 sky130_fd_sc_hd__xnor2_1 _10725_ (.A(_03306_),
    .B(_03307_),
    .Y(_03308_));
 sky130_fd_sc_hd__and4_2 _10726_ (.A(_02960_),
    .B(_02955_),
    .C(_03247_),
    .D(_03233_),
    .X(_03309_));
 sky130_fd_sc_hd__a22o_1 _10727_ (.A1(_02966_),
    .A2(_03247_),
    .B1(_03271_),
    .B2(_02964_),
    .X(_03310_));
 sky130_fd_sc_hd__and2b_1 _10728_ (.A_N(_03309_),
    .B(_03310_),
    .X(_03311_));
 sky130_fd_sc_hd__nand2_1 _10729_ (.A(_03100_),
    .B(_03129_),
    .Y(_03312_));
 sky130_fd_sc_hd__xnor2_1 _10730_ (.A(_03311_),
    .B(_03312_),
    .Y(_03313_));
 sky130_fd_sc_hd__buf_4 _10731_ (.A(_03229_),
    .X(_03314_));
 sky130_fd_sc_hd__nand2_2 _10732_ (.A(_03015_),
    .B(_03314_),
    .Y(_03315_));
 sky130_fd_sc_hd__nand2_1 _10733_ (.A(_03020_),
    .B(_03278_),
    .Y(_03316_));
 sky130_fd_sc_hd__xor2_1 _10734_ (.A(_03315_),
    .B(_03316_),
    .X(_03317_));
 sky130_fd_sc_hd__xor2_1 _10735_ (.A(_03313_),
    .B(_03317_),
    .X(_03318_));
 sky130_fd_sc_hd__a2bb2o_1 _10736_ (.A1_N(_03316_),
    .A2_N(_03282_),
    .B1(_03284_),
    .B2(_03277_),
    .X(_03319_));
 sky130_fd_sc_hd__and2_1 _10737_ (.A(_03318_),
    .B(_03319_),
    .X(_03320_));
 sky130_fd_sc_hd__nor2_1 _10738_ (.A(_03318_),
    .B(_03319_),
    .Y(_03321_));
 sky130_fd_sc_hd__nor2_1 _10739_ (.A(_03320_),
    .B(_03321_),
    .Y(_03322_));
 sky130_fd_sc_hd__and2_1 _10740_ (.A(_03308_),
    .B(_03322_),
    .X(_03323_));
 sky130_fd_sc_hd__nor2_1 _10741_ (.A(_03308_),
    .B(_03322_),
    .Y(_03324_));
 sky130_fd_sc_hd__a211o_1 _10742_ (.A1(_03295_),
    .A2(_03298_),
    .B1(_03323_),
    .C1(_03324_),
    .X(_03325_));
 sky130_fd_sc_hd__or3_1 _10743_ (.A(_03265_),
    .B(_03262_),
    .C(_03264_),
    .X(_03326_));
 sky130_fd_sc_hd__o211ai_1 _10744_ (.A1(_03323_),
    .A2(_03324_),
    .B1(_03295_),
    .C1(_03298_),
    .Y(_03327_));
 sky130_fd_sc_hd__and4_1 _10745_ (.A(_03325_),
    .B(_03266_),
    .C(_03326_),
    .D(_03327_),
    .X(_03328_));
 sky130_fd_sc_hd__inv_2 _10746_ (.A(_03328_),
    .Y(_03329_));
 sky130_fd_sc_hd__or2b_1 _10747_ (.A(_03223_),
    .B_N(_03216_),
    .X(_03330_));
 sky130_fd_sc_hd__or2b_1 _10748_ (.A(_03299_),
    .B_N(_03305_),
    .X(_03331_));
 sky130_fd_sc_hd__or2b_1 _10749_ (.A(_03307_),
    .B_N(_03306_),
    .X(_03332_));
 sky130_fd_sc_hd__a31o_1 _10750_ (.A1(_02918_),
    .A2(_02889_),
    .A3(_03214_),
    .B1(_03211_),
    .X(_03333_));
 sky130_fd_sc_hd__a22o_1 _10751_ (.A1(_02923_),
    .A2(_02888_),
    .B1(_02951_),
    .B2(_02921_),
    .X(_03334_));
 sky130_fd_sc_hd__a21bo_1 _10752_ (.A1(_02952_),
    .A2(_02924_),
    .B1_N(_03334_),
    .X(_03335_));
 sky130_fd_sc_hd__xor2_1 _10753_ (.A(_02928_),
    .B(_03335_),
    .X(_03336_));
 sky130_fd_sc_hd__xor2_1 _10754_ (.A(_03333_),
    .B(_03336_),
    .X(_03337_));
 sky130_fd_sc_hd__xnor2_1 _10755_ (.A(_02916_),
    .B(_03337_),
    .Y(_03338_));
 sky130_fd_sc_hd__a21oi_1 _10756_ (.A1(_03331_),
    .A2(_03332_),
    .B1(_03338_),
    .Y(_03339_));
 sky130_fd_sc_hd__and3_1 _10757_ (.A(_03331_),
    .B(_03332_),
    .C(_03338_),
    .X(_03340_));
 sky130_fd_sc_hd__or2_1 _10758_ (.A(_03339_),
    .B(_03340_),
    .X(_03341_));
 sky130_fd_sc_hd__a21oi_2 _10759_ (.A1(_03330_),
    .A2(_03225_),
    .B1(_03341_),
    .Y(_03342_));
 sky130_fd_sc_hd__o21ba_1 _10760_ (.A1(_03300_),
    .A2(_03303_),
    .B1_N(_03301_),
    .X(_03343_));
 sky130_fd_sc_hd__a31o_1 _10761_ (.A1(_03100_),
    .A2(_03129_),
    .A3(_03310_),
    .B1(_03309_),
    .X(_03344_));
 sky130_fd_sc_hd__nand2_1 _10762_ (.A(_03142_),
    .B(_03022_),
    .Y(_03345_));
 sky130_fd_sc_hd__and4_1 _10763_ (.A(_03145_),
    .B(_02939_),
    .C(_03220_),
    .D(_03039_),
    .X(_03346_));
 sky130_fd_sc_hd__a22oi_1 _10764_ (.A1(_03302_),
    .A2(_03220_),
    .B1(_03039_),
    .B2(_02969_),
    .Y(_03347_));
 sky130_fd_sc_hd__nor2_1 _10765_ (.A(_03346_),
    .B(_03347_),
    .Y(_03348_));
 sky130_fd_sc_hd__xnor2_1 _10766_ (.A(_03345_),
    .B(_03348_),
    .Y(_03349_));
 sky130_fd_sc_hd__xor2_1 _10767_ (.A(_03344_),
    .B(_03349_),
    .X(_03350_));
 sky130_fd_sc_hd__and2b_1 _10768_ (.A_N(_03343_),
    .B(_03350_),
    .X(_03351_));
 sky130_fd_sc_hd__and2b_1 _10769_ (.A_N(_03350_),
    .B(_03343_),
    .X(_03352_));
 sky130_fd_sc_hd__or2_1 _10770_ (.A(_03351_),
    .B(_03352_),
    .X(_03353_));
 sky130_fd_sc_hd__and4_2 _10771_ (.A(_02964_),
    .B(_02966_),
    .C(_03127_),
    .D(_03247_),
    .X(_03354_));
 sky130_fd_sc_hd__a22o_1 _10772_ (.A1(_02956_),
    .A2(_03128_),
    .B1(_03248_),
    .B2(_02961_),
    .X(_03355_));
 sky130_fd_sc_hd__or2b_1 _10773_ (.A(_03354_),
    .B_N(_03355_),
    .X(_03356_));
 sky130_fd_sc_hd__nand2_1 _10774_ (.A(_03100_),
    .B(_03095_),
    .Y(_03357_));
 sky130_fd_sc_hd__xnor2_1 _10775_ (.A(_03356_),
    .B(_03357_),
    .Y(_03358_));
 sky130_fd_sc_hd__nand2_1 _10776_ (.A(_03016_),
    .B(_03234_),
    .Y(_03359_));
 sky130_fd_sc_hd__nand2_1 _10777_ (.A(_03021_),
    .B(_03315_),
    .Y(_03360_));
 sky130_fd_sc_hd__xnor2_1 _10778_ (.A(_03359_),
    .B(_03360_),
    .Y(_03361_));
 sky130_fd_sc_hd__xnor2_1 _10779_ (.A(_03358_),
    .B(_03361_),
    .Y(_03362_));
 sky130_fd_sc_hd__a2bb2o_1 _10780_ (.A1_N(_03360_),
    .A2_N(_03278_),
    .B1(_03317_),
    .B2(_03313_),
    .X(_03363_));
 sky130_fd_sc_hd__and2b_1 _10781_ (.A_N(_03362_),
    .B(_03363_),
    .X(_03364_));
 sky130_fd_sc_hd__and2b_1 _10782_ (.A_N(_03363_),
    .B(_03362_),
    .X(_03365_));
 sky130_fd_sc_hd__or2_1 _10783_ (.A(_03364_),
    .B(_03365_),
    .X(_03366_));
 sky130_fd_sc_hd__nor2_2 _10784_ (.A(_03353_),
    .B(_03366_),
    .Y(_03367_));
 sky130_fd_sc_hd__and2_1 _10785_ (.A(_03353_),
    .B(_03366_),
    .X(_03368_));
 sky130_fd_sc_hd__nor2_1 _10786_ (.A(_03367_),
    .B(_03368_),
    .Y(_03369_));
 sky130_fd_sc_hd__o21a_1 _10787_ (.A1(_03320_),
    .A2(_03323_),
    .B1(_03369_),
    .X(_03370_));
 sky130_fd_sc_hd__and3_1 _10788_ (.A(_03341_),
    .B(_03330_),
    .C(_03225_),
    .X(_03371_));
 sky130_fd_sc_hd__nor3_1 _10789_ (.A(_03369_),
    .B(_03320_),
    .C(_03323_),
    .Y(_03372_));
 sky130_fd_sc_hd__nor4_2 _10790_ (.A(_03342_),
    .B(_03370_),
    .C(_03371_),
    .D(_03372_),
    .Y(_03373_));
 sky130_fd_sc_hd__o22a_1 _10791_ (.A1(_03342_),
    .A2(_03371_),
    .B1(_03372_),
    .B2(_03370_),
    .X(_03374_));
 sky130_fd_sc_hd__a211oi_2 _10792_ (.A1(_03325_),
    .A2(_03329_),
    .B1(_03373_),
    .C1(_03374_),
    .Y(_03375_));
 sky130_fd_sc_hd__inv_2 _10793_ (.A(_03375_),
    .Y(_03376_));
 sky130_fd_sc_hd__xnor2_1 _10794_ (.A(_02980_),
    .B(_03269_),
    .Y(_03377_));
 sky130_fd_sc_hd__o211a_1 _10795_ (.A1(_03373_),
    .A2(_03374_),
    .B1(_03325_),
    .C1(_03329_),
    .X(_03378_));
 sky130_fd_sc_hd__or3_2 _10796_ (.A(_03375_),
    .B(_03377_),
    .C(_03378_),
    .X(_03379_));
 sky130_fd_sc_hd__a31o_1 _10797_ (.A1(_02950_),
    .A2(_03095_),
    .A3(_03355_),
    .B1(_03354_),
    .X(_03380_));
 sky130_fd_sc_hd__nand2_1 _10798_ (.A(_03142_),
    .B(_02952_),
    .Y(_03381_));
 sky130_fd_sc_hd__and4_1 _10799_ (.A(_02969_),
    .B(_03302_),
    .C(_02987_),
    .D(_03029_),
    .X(_03382_));
 sky130_fd_sc_hd__a22oi_1 _10800_ (.A1(_03302_),
    .A2(_02987_),
    .B1(_03029_),
    .B2(_02969_),
    .Y(_03383_));
 sky130_fd_sc_hd__nor2_1 _10801_ (.A(_03382_),
    .B(_03383_),
    .Y(_03384_));
 sky130_fd_sc_hd__xnor2_1 _10802_ (.A(_03381_),
    .B(_03384_),
    .Y(_03385_));
 sky130_fd_sc_hd__xor2_1 _10803_ (.A(_03380_),
    .B(_03385_),
    .X(_03386_));
 sky130_fd_sc_hd__o21ba_1 _10804_ (.A1(_03345_),
    .A2(_03347_),
    .B1_N(_03346_),
    .X(_03387_));
 sky130_fd_sc_hd__xnor2_1 _10805_ (.A(_03386_),
    .B(_03387_),
    .Y(_03388_));
 sky130_fd_sc_hd__and4_1 _10806_ (.A(_02988_),
    .B(_02986_),
    .C(_03094_),
    .D(_03128_),
    .X(_03389_));
 sky130_fd_sc_hd__a22o_1 _10807_ (.A1(_02986_),
    .A2(_03094_),
    .B1(_03129_),
    .B2(_02988_),
    .X(_03390_));
 sky130_fd_sc_hd__and2b_1 _10808_ (.A_N(_03389_),
    .B(_03390_),
    .X(_03391_));
 sky130_fd_sc_hd__nand2_1 _10809_ (.A(_02950_),
    .B(_03040_),
    .Y(_03392_));
 sky130_fd_sc_hd__xnor2_1 _10810_ (.A(_03391_),
    .B(_03392_),
    .Y(_03393_));
 sky130_fd_sc_hd__nand2_2 _10811_ (.A(_03015_),
    .B(_03274_),
    .Y(_03394_));
 sky130_fd_sc_hd__nand2_1 _10812_ (.A(_03021_),
    .B(_03359_),
    .Y(_03395_));
 sky130_fd_sc_hd__xor2_1 _10813_ (.A(_03394_),
    .B(_03395_),
    .X(_03396_));
 sky130_fd_sc_hd__xor2_1 _10814_ (.A(_03393_),
    .B(_03396_),
    .X(_03397_));
 sky130_fd_sc_hd__o22ai_1 _10815_ (.A1(_03395_),
    .A2(_03315_),
    .B1(_03361_),
    .B2(_03358_),
    .Y(_03398_));
 sky130_fd_sc_hd__nand2_1 _10816_ (.A(_03397_),
    .B(_03398_),
    .Y(_03399_));
 sky130_fd_sc_hd__or2_1 _10817_ (.A(_03397_),
    .B(_03398_),
    .X(_03400_));
 sky130_fd_sc_hd__and2_1 _10818_ (.A(_03399_),
    .B(_03400_),
    .X(_03401_));
 sky130_fd_sc_hd__nand2_2 _10819_ (.A(_03388_),
    .B(_03401_),
    .Y(_03402_));
 sky130_fd_sc_hd__or2_1 _10820_ (.A(_03388_),
    .B(_03401_),
    .X(_03403_));
 sky130_fd_sc_hd__o211ai_4 _10821_ (.A1(_03364_),
    .A2(_03367_),
    .B1(_03402_),
    .C1(_03403_),
    .Y(_03404_));
 sky130_fd_sc_hd__and2_1 _10822_ (.A(_03344_),
    .B(_03349_),
    .X(_03405_));
 sky130_fd_sc_hd__or2_1 _10823_ (.A(_02924_),
    .B(_02929_),
    .X(_03406_));
 sky130_fd_sc_hd__nand2_1 _10824_ (.A(_02953_),
    .B(_02924_),
    .Y(_03407_));
 sky130_fd_sc_hd__a22o_1 _10825_ (.A1(_02928_),
    .A2(_03407_),
    .B1(_03334_),
    .B2(_02918_),
    .X(_03408_));
 sky130_fd_sc_hd__xnor2_1 _10826_ (.A(_03406_),
    .B(_03408_),
    .Y(_03409_));
 sky130_fd_sc_hd__xnor2_1 _10827_ (.A(_02916_),
    .B(_03409_),
    .Y(_03410_));
 sky130_fd_sc_hd__o21ai_1 _10828_ (.A1(_03405_),
    .A2(_03351_),
    .B1(_03410_),
    .Y(_03411_));
 sky130_fd_sc_hd__or3_1 _10829_ (.A(_03405_),
    .B(_03351_),
    .C(_03410_),
    .X(_03412_));
 sky130_fd_sc_hd__and2_1 _10830_ (.A(_03411_),
    .B(_03412_),
    .X(_03413_));
 sky130_fd_sc_hd__and2_1 _10831_ (.A(_03333_),
    .B(_03336_),
    .X(_03414_));
 sky130_fd_sc_hd__a21oi_1 _10832_ (.A1(_02916_),
    .A2(_03337_),
    .B1(_03414_),
    .Y(_03415_));
 sky130_fd_sc_hd__xnor2_1 _10833_ (.A(_03413_),
    .B(_03415_),
    .Y(_03416_));
 sky130_fd_sc_hd__a211o_1 _10834_ (.A1(_03402_),
    .A2(_03403_),
    .B1(_03364_),
    .C1(_03367_),
    .X(_03417_));
 sky130_fd_sc_hd__nand3_1 _10835_ (.A(_03404_),
    .B(_03416_),
    .C(_03417_),
    .Y(_03418_));
 sky130_fd_sc_hd__a21o_1 _10836_ (.A1(_03404_),
    .A2(_03417_),
    .B1(_03416_),
    .X(_03419_));
 sky130_fd_sc_hd__and2_1 _10837_ (.A(_03418_),
    .B(_03419_),
    .X(_03420_));
 sky130_fd_sc_hd__o21a_2 _10838_ (.A1(_03370_),
    .A2(_03373_),
    .B1(_03420_),
    .X(_03421_));
 sky130_fd_sc_hd__o21a_1 _10839_ (.A1(_03339_),
    .A2(_03342_),
    .B1(_02913_),
    .X(_03422_));
 sky130_fd_sc_hd__nor3_1 _10840_ (.A(_02913_),
    .B(_03339_),
    .C(_03342_),
    .Y(_03423_));
 sky130_fd_sc_hd__nor2_1 _10841_ (.A(_03422_),
    .B(_03423_),
    .Y(_03424_));
 sky130_fd_sc_hd__xnor2_2 _10842_ (.A(_02981_),
    .B(_03424_),
    .Y(_03425_));
 sky130_fd_sc_hd__nor3_2 _10843_ (.A(_03420_),
    .B(_03370_),
    .C(_03373_),
    .Y(_03426_));
 sky130_fd_sc_hd__nor3_4 _10844_ (.A(_03421_),
    .B(_03425_),
    .C(_03426_),
    .Y(_03427_));
 sky130_fd_sc_hd__o21a_1 _10845_ (.A1(_03421_),
    .A2(_03426_),
    .B1(_03425_),
    .X(_03428_));
 sky130_fd_sc_hd__a211oi_4 _10846_ (.A1(_03376_),
    .A2(_03379_),
    .B1(_03427_),
    .C1(_03428_),
    .Y(_03429_));
 sky130_fd_sc_hd__o211a_1 _10847_ (.A1(_03427_),
    .A2(_03428_),
    .B1(_03376_),
    .C1(_03379_),
    .X(_03430_));
 sky130_fd_sc_hd__a211oi_4 _10848_ (.A1(_03268_),
    .A2(_03270_),
    .B1(_03429_),
    .C1(_03430_),
    .Y(_03431_));
 sky130_fd_sc_hd__o211a_1 _10849_ (.A1(_03429_),
    .A2(_03430_),
    .B1(_03268_),
    .C1(_03270_),
    .X(_03432_));
 sky130_fd_sc_hd__xor2_1 _10850_ (.A(_03293_),
    .B(_03291_),
    .X(_03433_));
 sky130_fd_sc_hd__clkbuf_4 _10851_ (.A(_03069_),
    .X(_03434_));
 sky130_fd_sc_hd__buf_8 _10852_ (.A(_03434_),
    .X(_03435_));
 sky130_fd_sc_hd__buf_4 _10853_ (.A(net10),
    .X(_03436_));
 sky130_fd_sc_hd__buf_4 _10854_ (.A(_03436_),
    .X(_03437_));
 sky130_fd_sc_hd__nor2_1 _10855_ (.A(_03288_),
    .B(_03071_),
    .Y(_03438_));
 sky130_fd_sc_hd__nand2_1 _10856_ (.A(_03015_),
    .B(_03437_),
    .Y(_03439_));
 sky130_fd_sc_hd__and2_1 _10857_ (.A(_03020_),
    .B(_03439_),
    .X(_03440_));
 sky130_fd_sc_hd__xnor2_1 _10858_ (.A(_03289_),
    .B(_03440_),
    .Y(_03441_));
 sky130_fd_sc_hd__and4_1 _10859_ (.A(_02964_),
    .B(_02966_),
    .C(_03236_),
    .D(_03280_),
    .X(_03442_));
 sky130_fd_sc_hd__a22o_1 _10860_ (.A1(_02966_),
    .A2(_03236_),
    .B1(_03280_),
    .B2(_02964_),
    .X(_03443_));
 sky130_fd_sc_hd__and2b_1 _10861_ (.A_N(_03442_),
    .B(_03443_),
    .X(_03444_));
 sky130_fd_sc_hd__nand2_1 _10862_ (.A(_03100_),
    .B(_03314_),
    .Y(_03445_));
 sky130_fd_sc_hd__xnor2_1 _10863_ (.A(_03444_),
    .B(_03445_),
    .Y(_03446_));
 sky130_fd_sc_hd__a32o_1 _10864_ (.A1(_03435_),
    .A2(_03437_),
    .A3(_03438_),
    .B1(_03441_),
    .B2(_03446_),
    .X(_03447_));
 sky130_fd_sc_hd__nand2_1 _10865_ (.A(_03433_),
    .B(_03447_),
    .Y(_03448_));
 sky130_fd_sc_hd__a31o_1 _10866_ (.A1(_03100_),
    .A2(_03314_),
    .A3(_03443_),
    .B1(_03442_),
    .X(_03449_));
 sky130_fd_sc_hd__nor2_1 _10867_ (.A(_03250_),
    .B(_03249_),
    .Y(_03450_));
 sky130_fd_sc_hd__xnor2_1 _10868_ (.A(_03246_),
    .B(_03450_),
    .Y(_03451_));
 sky130_fd_sc_hd__xor2_1 _10869_ (.A(_03449_),
    .B(_03451_),
    .X(_03452_));
 sky130_fd_sc_hd__nand2_1 _10870_ (.A(_03142_),
    .B(_03129_),
    .Y(_03453_));
 sky130_fd_sc_hd__a22oi_1 _10871_ (.A1(_02939_),
    .A2(_03274_),
    .B1(_03234_),
    .B2(_03145_),
    .Y(_03454_));
 sky130_fd_sc_hd__and4_1 _10872_ (.A(_03145_),
    .B(_02939_),
    .C(_03248_),
    .D(_03271_),
    .X(_03455_));
 sky130_fd_sc_hd__o21ba_1 _10873_ (.A1(_03453_),
    .A2(_03454_),
    .B1_N(_03455_),
    .X(_03456_));
 sky130_fd_sc_hd__xnor2_1 _10874_ (.A(_03452_),
    .B(_03456_),
    .Y(_03457_));
 sky130_fd_sc_hd__xor2_1 _10875_ (.A(_03433_),
    .B(_03447_),
    .X(_03458_));
 sky130_fd_sc_hd__nand2_1 _10876_ (.A(_03457_),
    .B(_03458_),
    .Y(_03459_));
 sky130_fd_sc_hd__xnor2_1 _10877_ (.A(_03296_),
    .B(_03297_),
    .Y(_03460_));
 sky130_fd_sc_hd__a21o_1 _10878_ (.A1(_03448_),
    .A2(_03459_),
    .B1(_03460_),
    .X(_03461_));
 sky130_fd_sc_hd__nand2_1 _10879_ (.A(_03449_),
    .B(_03451_),
    .Y(_03462_));
 sky130_fd_sc_hd__or2b_1 _10880_ (.A(_03456_),
    .B_N(_03452_),
    .X(_03463_));
 sky130_fd_sc_hd__xnor2_1 _10881_ (.A(_02916_),
    .B(_03263_),
    .Y(_03464_));
 sky130_fd_sc_hd__a21oi_1 _10882_ (.A1(_03462_),
    .A2(_03463_),
    .B1(_03464_),
    .Y(_03465_));
 sky130_fd_sc_hd__and3_1 _10883_ (.A(_03462_),
    .B(_03463_),
    .C(_03464_),
    .X(_03466_));
 sky130_fd_sc_hd__nor2_1 _10884_ (.A(_03465_),
    .B(_03466_),
    .Y(_03467_));
 sky130_fd_sc_hd__o2bb2a_1 _10885_ (.A1_N(_02918_),
    .A2_N(_02987_),
    .B1(_03256_),
    .B2(_03257_),
    .X(_03468_));
 sky130_fd_sc_hd__and4_1 _10886_ (.A(_03218_),
    .B(_03210_),
    .C(_03038_),
    .D(_03093_),
    .X(_03469_));
 sky130_fd_sc_hd__a22oi_1 _10887_ (.A1(_02923_),
    .A2(_03038_),
    .B1(_03094_),
    .B2(_02921_),
    .Y(_03470_));
 sky130_fd_sc_hd__and4bb_1 _10888_ (.A_N(_03469_),
    .B_N(_03470_),
    .C(_02927_),
    .D(_03220_),
    .X(_03471_));
 sky130_fd_sc_hd__nor2_1 _10889_ (.A(_03469_),
    .B(_03471_),
    .Y(_03472_));
 sky130_fd_sc_hd__nor2_1 _10890_ (.A(_03258_),
    .B(_03468_),
    .Y(_03473_));
 sky130_fd_sc_hd__xnor2_1 _10891_ (.A(_03473_),
    .B(_03472_),
    .Y(_03474_));
 sky130_fd_sc_hd__nand2_1 _10892_ (.A(_02895_),
    .B(_02952_),
    .Y(_03475_));
 sky130_fd_sc_hd__xnor2_1 _10893_ (.A(_02901_),
    .B(_03475_),
    .Y(_03476_));
 sky130_fd_sc_hd__xnor2_1 _10894_ (.A(_02893_),
    .B(_03476_),
    .Y(_03477_));
 sky130_fd_sc_hd__nand2_1 _10895_ (.A(_03474_),
    .B(_03477_),
    .Y(_03478_));
 sky130_fd_sc_hd__o31a_1 _10896_ (.A1(_03258_),
    .A2(_03468_),
    .A3(_03472_),
    .B1(_03478_),
    .X(_03479_));
 sky130_fd_sc_hd__xnor2_1 _10897_ (.A(_03467_),
    .B(_03479_),
    .Y(_03480_));
 sky130_fd_sc_hd__nand3_1 _10898_ (.A(_03448_),
    .B(_03459_),
    .C(_03460_),
    .Y(_03481_));
 sky130_fd_sc_hd__nand3_1 _10899_ (.A(_03461_),
    .B(_03480_),
    .C(_03481_),
    .Y(_03482_));
 sky130_fd_sc_hd__a22oi_2 _10900_ (.A1(_03266_),
    .A2(_03326_),
    .B1(_03327_),
    .B2(_03325_),
    .Y(_03483_));
 sky130_fd_sc_hd__a211oi_2 _10901_ (.A1(_03461_),
    .A2(_03482_),
    .B1(_03328_),
    .C1(_03483_),
    .Y(_03484_));
 sky130_fd_sc_hd__and2b_1 _10902_ (.A_N(_03479_),
    .B(_03467_),
    .X(_03485_));
 sky130_fd_sc_hd__o21ai_2 _10903_ (.A1(_03465_),
    .A2(_03485_),
    .B1(_02912_),
    .Y(_03486_));
 sky130_fd_sc_hd__or3_1 _10904_ (.A(_02912_),
    .B(_03465_),
    .C(_03485_),
    .X(_03487_));
 sky130_fd_sc_hd__and2_1 _10905_ (.A(_03486_),
    .B(_03487_),
    .X(_03488_));
 sky130_fd_sc_hd__and3_1 _10906_ (.A(_02895_),
    .B(_02953_),
    .C(_02901_),
    .X(_03489_));
 sky130_fd_sc_hd__buf_4 _10907_ (.A(\wfg_stim_mem_top.cfg_gain_q[9] ),
    .X(_03490_));
 sky130_fd_sc_hd__buf_4 _10908_ (.A(_03490_),
    .X(_03491_));
 sky130_fd_sc_hd__buf_8 _10909_ (.A(_03491_),
    .X(_03492_));
 sky130_fd_sc_hd__and3_1 _10910_ (.A(_03492_),
    .B(_02910_),
    .C(_03476_),
    .X(_03493_));
 sky130_fd_sc_hd__or3_1 _10911_ (.A(_02891_),
    .B(_03489_),
    .C(_03493_),
    .X(_03494_));
 sky130_fd_sc_hd__o21a_1 _10912_ (.A1(_03489_),
    .A2(_03493_),
    .B1(_02891_),
    .X(_03495_));
 sky130_fd_sc_hd__a31o_1 _10913_ (.A1(_02909_),
    .A2(_02910_),
    .A3(_03494_),
    .B1(_03495_),
    .X(_03496_));
 sky130_fd_sc_hd__xnor2_1 _10914_ (.A(_03488_),
    .B(_03496_),
    .Y(_03497_));
 sky130_fd_sc_hd__o211a_1 _10915_ (.A1(_03328_),
    .A2(_03483_),
    .B1(_03461_),
    .C1(_03482_),
    .X(_03498_));
 sky130_fd_sc_hd__nor2_1 _10916_ (.A(_03484_),
    .B(_03498_),
    .Y(_03499_));
 sky130_fd_sc_hd__and2b_1 _10917_ (.A_N(_03497_),
    .B(_03499_),
    .X(_03500_));
 sky130_fd_sc_hd__o21ai_1 _10918_ (.A1(_03375_),
    .A2(_03378_),
    .B1(_03377_),
    .Y(_03501_));
 sky130_fd_sc_hd__o211a_1 _10919_ (.A1(_03484_),
    .A2(_03500_),
    .B1(_03501_),
    .C1(_03379_),
    .X(_03502_));
 sky130_fd_sc_hd__inv_2 _10920_ (.A(_03502_),
    .Y(_03503_));
 sky130_fd_sc_hd__nand2_1 _10921_ (.A(_03488_),
    .B(_03496_),
    .Y(_03504_));
 sky130_fd_sc_hd__a211oi_2 _10922_ (.A1(_03379_),
    .A2(_03501_),
    .B1(_03500_),
    .C1(_03484_),
    .Y(_03505_));
 sky130_fd_sc_hd__a211o_1 _10923_ (.A1(_03486_),
    .A2(_03504_),
    .B1(_03502_),
    .C1(_03505_),
    .X(_03506_));
 sky130_fd_sc_hd__o211a_1 _10924_ (.A1(_03431_),
    .A2(_03432_),
    .B1(_03503_),
    .C1(_03506_),
    .X(_03507_));
 sky130_fd_sc_hd__nand2_1 _10925_ (.A(_03461_),
    .B(_03481_),
    .Y(_03508_));
 sky130_fd_sc_hd__xor2_1 _10926_ (.A(_03480_),
    .B(_03508_),
    .X(_03509_));
 sky130_fd_sc_hd__a22oi_1 _10927_ (.A1(_02986_),
    .A2(_03281_),
    .B1(_03288_),
    .B2(_02988_),
    .Y(_03510_));
 sky130_fd_sc_hd__nand2_1 _10928_ (.A(_02949_),
    .B(_03231_),
    .Y(_03511_));
 sky130_fd_sc_hd__and4_1 _10929_ (.A(_02961_),
    .B(_02956_),
    .C(_03280_),
    .D(_03287_),
    .X(_03512_));
 sky130_fd_sc_hd__o21ba_1 _10930_ (.A1(_03510_),
    .A2(_03511_),
    .B1_N(_03512_),
    .X(_03513_));
 sky130_fd_sc_hd__nor2_1 _10931_ (.A(_03455_),
    .B(_03454_),
    .Y(_03514_));
 sky130_fd_sc_hd__xnor2_1 _10932_ (.A(_03453_),
    .B(_03514_),
    .Y(_03515_));
 sky130_fd_sc_hd__or2b_1 _10933_ (.A(_03513_),
    .B_N(_03515_),
    .X(_03516_));
 sky130_fd_sc_hd__nand2_1 _10934_ (.A(_03239_),
    .B(_03274_),
    .Y(_03517_));
 sky130_fd_sc_hd__a22oi_1 _10935_ (.A1(_02939_),
    .A2(_03234_),
    .B1(_03314_),
    .B2(_03145_),
    .Y(_03518_));
 sky130_fd_sc_hd__and4_1 _10936_ (.A(_03145_),
    .B(_02939_),
    .C(_03271_),
    .D(_03229_),
    .X(_03519_));
 sky130_fd_sc_hd__o21ba_1 _10937_ (.A1(_03517_),
    .A2(_03518_),
    .B1_N(_03519_),
    .X(_03520_));
 sky130_fd_sc_hd__xnor2_1 _10938_ (.A(_03513_),
    .B(_03515_),
    .Y(_03521_));
 sky130_fd_sc_hd__or2b_1 _10939_ (.A(_03520_),
    .B_N(_03521_),
    .X(_03522_));
 sky130_fd_sc_hd__xnor2_1 _10940_ (.A(_03474_),
    .B(_03477_),
    .Y(_03523_));
 sky130_fd_sc_hd__a21oi_2 _10941_ (.A1(_03516_),
    .A2(_03522_),
    .B1(_03523_),
    .Y(_03524_));
 sky130_fd_sc_hd__and3_1 _10942_ (.A(_03516_),
    .B(_03522_),
    .C(_03523_),
    .X(_03525_));
 sky130_fd_sc_hd__o2bb2a_1 _10943_ (.A1_N(_02927_),
    .A2_N(_03220_),
    .B1(_03469_),
    .B2(_03470_),
    .X(_03526_));
 sky130_fd_sc_hd__nor2_1 _10944_ (.A(_03471_),
    .B(_03526_),
    .Y(_03527_));
 sky130_fd_sc_hd__and4_1 _10945_ (.A(_03217_),
    .B(_03212_),
    .C(_03093_),
    .D(_03127_),
    .X(_03528_));
 sky130_fd_sc_hd__buf_4 _10946_ (.A(\wfg_stim_mem_top.cfg_gain_q[14] ),
    .X(_03529_));
 sky130_fd_sc_hd__nand2_1 _10947_ (.A(_03529_),
    .B(_03038_),
    .Y(_03530_));
 sky130_fd_sc_hd__buf_4 _10948_ (.A(_03209_),
    .X(_03531_));
 sky130_fd_sc_hd__buf_4 _10949_ (.A(_02919_),
    .X(_03532_));
 sky130_fd_sc_hd__a22oi_1 _10950_ (.A1(_03531_),
    .A2(_03093_),
    .B1(_03127_),
    .B2(_03532_),
    .Y(_03533_));
 sky130_fd_sc_hd__or3_1 _10951_ (.A(_03530_),
    .B(_03528_),
    .C(_03533_),
    .X(_03534_));
 sky130_fd_sc_hd__or2b_1 _10952_ (.A(_03528_),
    .B_N(_03534_),
    .X(_03535_));
 sky130_fd_sc_hd__xor2_1 _10953_ (.A(_03527_),
    .B(_03535_),
    .X(_03536_));
 sky130_fd_sc_hd__nand2_1 _10954_ (.A(_02900_),
    .B(_02957_),
    .Y(_03537_));
 sky130_fd_sc_hd__a22o_1 _10955_ (.A1(_02897_),
    .A2(_02952_),
    .B1(_02987_),
    .B2(_02895_),
    .X(_03538_));
 sky130_fd_sc_hd__o21a_1 _10956_ (.A1(_03537_),
    .A2(_03475_),
    .B1(_03538_),
    .X(_03539_));
 sky130_fd_sc_hd__xnor2_1 _10957_ (.A(_02893_),
    .B(_03539_),
    .Y(_03540_));
 sky130_fd_sc_hd__and2_1 _10958_ (.A(_03536_),
    .B(_03540_),
    .X(_03541_));
 sky130_fd_sc_hd__a21oi_1 _10959_ (.A1(_03527_),
    .A2(_03535_),
    .B1(_03541_),
    .Y(_03542_));
 sky130_fd_sc_hd__nor3_1 _10960_ (.A(_03524_),
    .B(_03525_),
    .C(_03542_),
    .Y(_03543_));
 sky130_fd_sc_hd__o21a_1 _10961_ (.A1(_03524_),
    .A2(_03525_),
    .B1(_03542_),
    .X(_03544_));
 sky130_fd_sc_hd__or2_1 _10962_ (.A(_03543_),
    .B(_03544_),
    .X(_03545_));
 sky130_fd_sc_hd__xnor2_1 _10963_ (.A(_03457_),
    .B(_03458_),
    .Y(_03546_));
 sky130_fd_sc_hd__xnor2_1 _10964_ (.A(_03521_),
    .B(_03520_),
    .Y(_03547_));
 sky130_fd_sc_hd__xor2_1 _10965_ (.A(_03446_),
    .B(_03441_),
    .X(_03548_));
 sky130_fd_sc_hd__nor2_1 _10966_ (.A(_03512_),
    .B(_03510_),
    .Y(_03549_));
 sky130_fd_sc_hd__xnor2_2 _10967_ (.A(_03549_),
    .B(_03511_),
    .Y(_03550_));
 sky130_fd_sc_hd__clkbuf_8 _10968_ (.A(net9),
    .X(_03551_));
 sky130_fd_sc_hd__nand4_4 _10969_ (.A(_03014_),
    .B(_03019_),
    .C(_02951_),
    .D(_03551_),
    .Y(_03552_));
 sky130_fd_sc_hd__xnor2_2 _10970_ (.A(_03070_),
    .B(_03439_),
    .Y(_03553_));
 sky130_fd_sc_hd__xor2_2 _10971_ (.A(_03552_),
    .B(_03553_),
    .X(_03554_));
 sky130_fd_sc_hd__nor2_1 _10972_ (.A(_03552_),
    .B(_03553_),
    .Y(_03555_));
 sky130_fd_sc_hd__a21o_1 _10973_ (.A1(_03550_),
    .A2(_03554_),
    .B1(_03555_),
    .X(_03556_));
 sky130_fd_sc_hd__xor2_1 _10974_ (.A(_03548_),
    .B(_03556_),
    .X(_03557_));
 sky130_fd_sc_hd__and2_1 _10975_ (.A(_03548_),
    .B(_03556_),
    .X(_03558_));
 sky130_fd_sc_hd__a21oi_1 _10976_ (.A1(_03547_),
    .A2(_03557_),
    .B1(_03558_),
    .Y(_03559_));
 sky130_fd_sc_hd__nor2_1 _10977_ (.A(_03546_),
    .B(_03559_),
    .Y(_03560_));
 sky130_fd_sc_hd__and2_1 _10978_ (.A(_03546_),
    .B(_03559_),
    .X(_03561_));
 sky130_fd_sc_hd__or2_1 _10979_ (.A(_03560_),
    .B(_03561_),
    .X(_03562_));
 sky130_fd_sc_hd__o21ba_1 _10980_ (.A1(_03545_),
    .A2(_03562_),
    .B1_N(_03560_),
    .X(_03563_));
 sky130_fd_sc_hd__and2b_1 _10981_ (.A_N(_03495_),
    .B(_03494_),
    .X(_03564_));
 sky130_fd_sc_hd__xnor2_1 _10982_ (.A(_02911_),
    .B(_03564_),
    .Y(_03565_));
 sky130_fd_sc_hd__o21ai_1 _10983_ (.A1(_03524_),
    .A2(_03543_),
    .B1(_03565_),
    .Y(_03566_));
 sky130_fd_sc_hd__or3_1 _10984_ (.A(_03524_),
    .B(_03543_),
    .C(_03565_),
    .X(_03567_));
 sky130_fd_sc_hd__and2_1 _10985_ (.A(_03566_),
    .B(_03567_),
    .X(_03568_));
 sky130_fd_sc_hd__nor2_1 _10986_ (.A(_03537_),
    .B(_03475_),
    .Y(_03569_));
 sky130_fd_sc_hd__a31o_1 _10987_ (.A1(_03492_),
    .A2(_02910_),
    .A3(_03538_),
    .B1(_03569_),
    .X(_03570_));
 sky130_fd_sc_hd__nor2_1 _10988_ (.A(_02891_),
    .B(_03570_),
    .Y(_03571_));
 sky130_fd_sc_hd__and2_1 _10989_ (.A(_02891_),
    .B(_03570_),
    .X(_03572_));
 sky130_fd_sc_hd__o21ba_1 _10990_ (.A1(_02911_),
    .A2(_03571_),
    .B1_N(_03572_),
    .X(_03573_));
 sky130_fd_sc_hd__xor2_1 _10991_ (.A(_03568_),
    .B(_03573_),
    .X(_03574_));
 sky130_fd_sc_hd__xnor2_1 _10992_ (.A(_03509_),
    .B(_03563_),
    .Y(_03575_));
 sky130_fd_sc_hd__nor2_1 _10993_ (.A(_03574_),
    .B(_03575_),
    .Y(_03576_));
 sky130_fd_sc_hd__o21ba_1 _10994_ (.A1(_03509_),
    .A2(_03563_),
    .B1_N(_03576_),
    .X(_03577_));
 sky130_fd_sc_hd__xnor2_1 _10995_ (.A(_03497_),
    .B(_03499_),
    .Y(_03578_));
 sky130_fd_sc_hd__or2b_1 _10996_ (.A(_03577_),
    .B_N(_03578_),
    .X(_03579_));
 sky130_fd_sc_hd__xor2_1 _10997_ (.A(_03578_),
    .B(_03577_),
    .X(_03580_));
 sky130_fd_sc_hd__or2b_1 _10998_ (.A(_03573_),
    .B_N(_03568_),
    .X(_03581_));
 sky130_fd_sc_hd__nand2_1 _10999_ (.A(_03566_),
    .B(_03581_),
    .Y(_03582_));
 sky130_fd_sc_hd__or2b_1 _11000_ (.A(_03580_),
    .B_N(_03582_),
    .X(_03583_));
 sky130_fd_sc_hd__a211oi_2 _11001_ (.A1(_03486_),
    .A2(_03504_),
    .B1(_03502_),
    .C1(_03505_),
    .Y(_03584_));
 sky130_fd_sc_hd__o211a_1 _11002_ (.A1(_03502_),
    .A2(_03505_),
    .B1(_03486_),
    .C1(_03504_),
    .X(_03585_));
 sky130_fd_sc_hd__a211oi_2 _11003_ (.A1(_03579_),
    .A2(_03583_),
    .B1(_03584_),
    .C1(_03585_),
    .Y(_03586_));
 sky130_fd_sc_hd__inv_2 _11004_ (.A(_03586_),
    .Y(_03587_));
 sky130_fd_sc_hd__a211oi_2 _11005_ (.A1(_03503_),
    .A2(_03506_),
    .B1(_03431_),
    .C1(_03432_),
    .Y(_03588_));
 sky130_fd_sc_hd__o211a_1 _11006_ (.A1(_03584_),
    .A2(_03585_),
    .B1(_03579_),
    .C1(_03583_),
    .X(_03589_));
 sky130_fd_sc_hd__or2_1 _11007_ (.A(_03586_),
    .B(_03589_),
    .X(_03590_));
 sky130_fd_sc_hd__or3_1 _11008_ (.A(_03588_),
    .B(_03507_),
    .C(_03590_),
    .X(_03591_));
 sky130_fd_sc_hd__xor2_1 _11009_ (.A(_03582_),
    .B(_03580_),
    .X(_03592_));
 sky130_fd_sc_hd__and2_1 _11010_ (.A(_03574_),
    .B(_03575_),
    .X(_03593_));
 sky130_fd_sc_hd__xnor2_1 _11011_ (.A(_03545_),
    .B(_03562_),
    .Y(_03594_));
 sky130_fd_sc_hd__xnor2_2 _11012_ (.A(_03550_),
    .B(_03554_),
    .Y(_03595_));
 sky130_fd_sc_hd__buf_4 _11013_ (.A(\wfg_stim_mem_top.cfg_gain_q[10] ),
    .X(_03596_));
 sky130_fd_sc_hd__buf_4 _11014_ (.A(net8),
    .X(_03597_));
 sky130_fd_sc_hd__and4_1 _11015_ (.A(_03014_),
    .B(_03596_),
    .C(net22),
    .D(_03597_),
    .X(_03598_));
 sky130_fd_sc_hd__a22o_1 _11016_ (.A1(_03019_),
    .A2(_02951_),
    .B1(_03551_),
    .B2(_03014_),
    .X(_03599_));
 sky130_fd_sc_hd__and3_1 _11017_ (.A(_03598_),
    .B(_03552_),
    .C(_03599_),
    .X(_03600_));
 sky130_fd_sc_hd__a21oi_1 _11018_ (.A1(_03552_),
    .A2(_03599_),
    .B1(_03598_),
    .Y(_03601_));
 sky130_fd_sc_hd__nand2_1 _11019_ (.A(_02949_),
    .B(_03281_),
    .Y(_03602_));
 sky130_fd_sc_hd__nand4_2 _11020_ (.A(_02961_),
    .B(_02956_),
    .C(_03288_),
    .D(_03437_),
    .Y(_03603_));
 sky130_fd_sc_hd__a22o_1 _11021_ (.A1(_02956_),
    .A2(_03287_),
    .B1(_03437_),
    .B2(_02961_),
    .X(_03604_));
 sky130_fd_sc_hd__nand3b_2 _11022_ (.A_N(_03602_),
    .B(_03603_),
    .C(_03604_),
    .Y(_03605_));
 sky130_fd_sc_hd__a21bo_1 _11023_ (.A1(_03603_),
    .A2(_03604_),
    .B1_N(_03602_),
    .X(_03606_));
 sky130_fd_sc_hd__or4bb_1 _11024_ (.A(_03600_),
    .B(_03601_),
    .C_N(_03605_),
    .D_N(_03606_),
    .X(_03607_));
 sky130_fd_sc_hd__or2b_2 _11025_ (.A(_03600_),
    .B_N(_03607_),
    .X(_03608_));
 sky130_fd_sc_hd__or2b_1 _11026_ (.A(_03595_),
    .B_N(_03608_),
    .X(_03609_));
 sky130_fd_sc_hd__xor2_2 _11027_ (.A(_03595_),
    .B(_03608_),
    .X(_03610_));
 sky130_fd_sc_hd__nand4_2 _11028_ (.A(_03145_),
    .B(_02939_),
    .C(_03229_),
    .D(_03231_),
    .Y(_03611_));
 sky130_fd_sc_hd__nand2_1 _11029_ (.A(_02935_),
    .B(_03271_),
    .Y(_03612_));
 sky130_fd_sc_hd__a22o_1 _11030_ (.A1(_02941_),
    .A2(_03229_),
    .B1(_03236_),
    .B2(_02944_),
    .X(_03613_));
 sky130_fd_sc_hd__nand3b_2 _11031_ (.A_N(_03612_),
    .B(_03611_),
    .C(_03613_),
    .Y(_03614_));
 sky130_fd_sc_hd__nand2_1 _11032_ (.A(_03611_),
    .B(_03614_),
    .Y(_03615_));
 sky130_fd_sc_hd__nand2_1 _11033_ (.A(_03603_),
    .B(_03605_),
    .Y(_03616_));
 sky130_fd_sc_hd__nor2_1 _11034_ (.A(_03519_),
    .B(_03518_),
    .Y(_03617_));
 sky130_fd_sc_hd__xnor2_1 _11035_ (.A(_03517_),
    .B(_03617_),
    .Y(_03618_));
 sky130_fd_sc_hd__xor2_2 _11036_ (.A(_03616_),
    .B(_03618_),
    .X(_03619_));
 sky130_fd_sc_hd__xor2_2 _11037_ (.A(_03615_),
    .B(_03619_),
    .X(_03620_));
 sky130_fd_sc_hd__or2b_1 _11038_ (.A(_03610_),
    .B_N(_03620_),
    .X(_03621_));
 sky130_fd_sc_hd__xnor2_1 _11039_ (.A(_03547_),
    .B(_03557_),
    .Y(_03622_));
 sky130_fd_sc_hd__a21oi_1 _11040_ (.A1(_03609_),
    .A2(_03621_),
    .B1(_03622_),
    .Y(_03623_));
 sky130_fd_sc_hd__and3_1 _11041_ (.A(_03609_),
    .B(_03621_),
    .C(_03622_),
    .X(_03624_));
 sky130_fd_sc_hd__nor2_1 _11042_ (.A(_03623_),
    .B(_03624_),
    .Y(_03625_));
 sky130_fd_sc_hd__o21ai_1 _11043_ (.A1(_03528_),
    .A2(_03533_),
    .B1(_03530_),
    .Y(_03626_));
 sky130_fd_sc_hd__nand2_1 _11044_ (.A(_02917_),
    .B(_03093_),
    .Y(_03627_));
 sky130_fd_sc_hd__a22oi_2 _11045_ (.A1(_03213_),
    .A2(_03127_),
    .B1(_03248_),
    .B2(_03218_),
    .Y(_03628_));
 sky130_fd_sc_hd__and4_1 _11046_ (.A(_02920_),
    .B(_02922_),
    .C(_03127_),
    .D(_03247_),
    .X(_03629_));
 sky130_fd_sc_hd__o21bai_1 _11047_ (.A1(_03627_),
    .A2(_03628_),
    .B1_N(_03629_),
    .Y(_03630_));
 sky130_fd_sc_hd__and3_1 _11048_ (.A(_03534_),
    .B(_03626_),
    .C(_03630_),
    .X(_03631_));
 sky130_fd_sc_hd__a21oi_1 _11049_ (.A1(_03534_),
    .A2(_03626_),
    .B1(_03630_),
    .Y(_03632_));
 sky130_fd_sc_hd__clkbuf_4 _11050_ (.A(\wfg_stim_mem_top.cfg_gain_q[13] ),
    .X(_03633_));
 sky130_fd_sc_hd__clkbuf_4 _11051_ (.A(_03633_),
    .X(_03634_));
 sky130_fd_sc_hd__nand2_1 _11052_ (.A(_03634_),
    .B(_03220_),
    .Y(_03635_));
 sky130_fd_sc_hd__buf_4 _11053_ (.A(\wfg_stim_mem_top.cfg_gain_q[13] ),
    .X(_03636_));
 sky130_fd_sc_hd__clkbuf_4 _11054_ (.A(\wfg_stim_mem_top.cfg_gain_q[12] ),
    .X(_03637_));
 sky130_fd_sc_hd__and4_1 _11055_ (.A(_03636_),
    .B(_03637_),
    .C(_02957_),
    .D(_02958_),
    .X(_03638_));
 sky130_fd_sc_hd__a21o_1 _11056_ (.A1(_03635_),
    .A2(_03537_),
    .B1(_03638_),
    .X(_03639_));
 sky130_fd_sc_hd__xor2_1 _11057_ (.A(_02893_),
    .B(_03639_),
    .X(_03640_));
 sky130_fd_sc_hd__or3b_1 _11058_ (.A(_03631_),
    .B(_03632_),
    .C_N(_03640_),
    .X(_03641_));
 sky130_fd_sc_hd__or2b_1 _11059_ (.A(_03631_),
    .B_N(_03641_),
    .X(_03642_));
 sky130_fd_sc_hd__nand2_1 _11060_ (.A(_03616_),
    .B(_03618_),
    .Y(_03643_));
 sky130_fd_sc_hd__a21boi_1 _11061_ (.A1(_03615_),
    .A2(_03619_),
    .B1_N(_03643_),
    .Y(_03644_));
 sky130_fd_sc_hd__xnor2_1 _11062_ (.A(_03536_),
    .B(_03540_),
    .Y(_03645_));
 sky130_fd_sc_hd__xnor2_1 _11063_ (.A(_03644_),
    .B(_03645_),
    .Y(_03646_));
 sky130_fd_sc_hd__xnor2_1 _11064_ (.A(_03642_),
    .B(_03646_),
    .Y(_03647_));
 sky130_fd_sc_hd__a21o_1 _11065_ (.A1(_03625_),
    .A2(_03647_),
    .B1(_03623_),
    .X(_03648_));
 sky130_fd_sc_hd__xor2_1 _11066_ (.A(_03594_),
    .B(_03648_),
    .X(_03649_));
 sky130_fd_sc_hd__nor2_1 _11067_ (.A(_03644_),
    .B(_03645_),
    .Y(_03650_));
 sky130_fd_sc_hd__and2b_1 _11068_ (.A_N(_03646_),
    .B(_03642_),
    .X(_03651_));
 sky130_fd_sc_hd__nor2_1 _11069_ (.A(_03572_),
    .B(_03571_),
    .Y(_03652_));
 sky130_fd_sc_hd__xnor2_1 _11070_ (.A(_02911_),
    .B(_03652_),
    .Y(_03653_));
 sky130_fd_sc_hd__o21ai_1 _11071_ (.A1(_03650_),
    .A2(_03651_),
    .B1(_03653_),
    .Y(_03654_));
 sky130_fd_sc_hd__or3_1 _11072_ (.A(_03650_),
    .B(_03651_),
    .C(_03653_),
    .X(_03655_));
 sky130_fd_sc_hd__and2_1 _11073_ (.A(_03654_),
    .B(_03655_),
    .X(_03656_));
 sky130_fd_sc_hd__nor2_1 _11074_ (.A(_02893_),
    .B(_03639_),
    .Y(_03657_));
 sky130_fd_sc_hd__or3_1 _11075_ (.A(_02890_),
    .B(_03638_),
    .C(_03657_),
    .X(_03658_));
 sky130_fd_sc_hd__o21a_1 _11076_ (.A1(_03638_),
    .A2(_03657_),
    .B1(_02891_),
    .X(_03659_));
 sky130_fd_sc_hd__a31oi_2 _11077_ (.A1(_02909_),
    .A2(_02910_),
    .A3(_03658_),
    .B1(_03659_),
    .Y(_03660_));
 sky130_fd_sc_hd__xor2_1 _11078_ (.A(_03656_),
    .B(_03660_),
    .X(_03661_));
 sky130_fd_sc_hd__and2b_1 _11079_ (.A_N(_03594_),
    .B(_03648_),
    .X(_03662_));
 sky130_fd_sc_hd__o21ba_1 _11080_ (.A1(_03649_),
    .A2(_03661_),
    .B1_N(_03662_),
    .X(_03663_));
 sky130_fd_sc_hd__or3_1 _11081_ (.A(_03576_),
    .B(_03593_),
    .C(_03663_),
    .X(_03664_));
 sky130_fd_sc_hd__nor2_1 _11082_ (.A(_03576_),
    .B(_03593_),
    .Y(_03665_));
 sky130_fd_sc_hd__xor2_1 _11083_ (.A(_03665_),
    .B(_03663_),
    .X(_03666_));
 sky130_fd_sc_hd__or2b_1 _11084_ (.A(_03660_),
    .B_N(_03656_),
    .X(_03667_));
 sky130_fd_sc_hd__nand2_1 _11085_ (.A(_03654_),
    .B(_03667_),
    .Y(_03668_));
 sky130_fd_sc_hd__or2b_1 _11086_ (.A(_03666_),
    .B_N(_03668_),
    .X(_03669_));
 sky130_fd_sc_hd__nand3_1 _11087_ (.A(_03592_),
    .B(_03664_),
    .C(_03669_),
    .Y(_03670_));
 sky130_fd_sc_hd__xnor2_1 _11088_ (.A(_03625_),
    .B(_03647_),
    .Y(_03671_));
 sky130_fd_sc_hd__xnor2_2 _11089_ (.A(_03610_),
    .B(_03620_),
    .Y(_03672_));
 sky130_fd_sc_hd__a2bb2o_1 _11090_ (.A1_N(_03600_),
    .A2_N(_03601_),
    .B1(_03605_),
    .B2(_03606_),
    .X(_03673_));
 sky130_fd_sc_hd__clkbuf_4 _11091_ (.A(net8),
    .X(_03674_));
 sky130_fd_sc_hd__buf_4 _11092_ (.A(_03674_),
    .X(_03675_));
 sky130_fd_sc_hd__nand4_1 _11093_ (.A(_03015_),
    .B(_03069_),
    .C(_02957_),
    .D(_03675_),
    .Y(_03676_));
 sky130_fd_sc_hd__a22o_1 _11094_ (.A1(_03019_),
    .A2(net22),
    .B1(_03597_),
    .B2(_03014_),
    .X(_03677_));
 sky130_fd_sc_hd__clkbuf_4 _11095_ (.A(\wfg_stim_mem_top.cfg_gain_q[23] ),
    .X(_03678_));
 sky130_fd_sc_hd__clkbuf_4 _11096_ (.A(\wfg_stim_mem_top.cfg_gain_q[10] ),
    .X(_03679_));
 sky130_fd_sc_hd__clkbuf_4 _11097_ (.A(net7),
    .X(_03680_));
 sky130_fd_sc_hd__and4_1 _11098_ (.A(_03678_),
    .B(_03679_),
    .C(net21),
    .D(_03680_),
    .X(_03681_));
 sky130_fd_sc_hd__a21o_1 _11099_ (.A1(_03676_),
    .A2(_03677_),
    .B1(_03681_),
    .X(_03682_));
 sky130_fd_sc_hd__and2_1 _11100_ (.A(_02949_),
    .B(_03287_),
    .X(_03683_));
 sky130_fd_sc_hd__buf_4 _11101_ (.A(net10),
    .X(_03684_));
 sky130_fd_sc_hd__clkbuf_4 _11102_ (.A(_03551_),
    .X(_03685_));
 sky130_fd_sc_hd__nand4_1 _11103_ (.A(_02964_),
    .B(_02966_),
    .C(_03684_),
    .D(_03685_),
    .Y(_03686_));
 sky130_fd_sc_hd__a22o_1 _11104_ (.A1(_02955_),
    .A2(_03684_),
    .B1(_03551_),
    .B2(_02960_),
    .X(_03687_));
 sky130_fd_sc_hd__nand3_1 _11105_ (.A(_03683_),
    .B(_03686_),
    .C(_03687_),
    .Y(_03688_));
 sky130_fd_sc_hd__a21o_1 _11106_ (.A1(_03686_),
    .A2(_03687_),
    .B1(_03683_),
    .X(_03689_));
 sky130_fd_sc_hd__and3_1 _11107_ (.A(_03681_),
    .B(_03676_),
    .C(_03677_),
    .X(_03690_));
 sky130_fd_sc_hd__a31o_1 _11108_ (.A1(_03682_),
    .A2(_03688_),
    .A3(_03689_),
    .B1(_03690_),
    .X(_03691_));
 sky130_fd_sc_hd__and3_1 _11109_ (.A(_03607_),
    .B(_03673_),
    .C(_03691_),
    .X(_03692_));
 sky130_fd_sc_hd__a21oi_1 _11110_ (.A1(_03607_),
    .A2(_03673_),
    .B1(_03691_),
    .Y(_03693_));
 sky130_fd_sc_hd__nand4_1 _11111_ (.A(_02944_),
    .B(_02941_),
    .C(_03236_),
    .D(_03280_),
    .Y(_03694_));
 sky130_fd_sc_hd__a22o_1 _11112_ (.A1(_02941_),
    .A2(_03236_),
    .B1(_03280_),
    .B2(_02944_),
    .X(_03695_));
 sky130_fd_sc_hd__nand4_1 _11113_ (.A(_03239_),
    .B(_03314_),
    .C(_03694_),
    .D(_03695_),
    .Y(_03696_));
 sky130_fd_sc_hd__nand2_1 _11114_ (.A(_03694_),
    .B(_03696_),
    .Y(_03697_));
 sky130_fd_sc_hd__a21bo_1 _11115_ (.A1(_03683_),
    .A2(_03687_),
    .B1_N(_03686_),
    .X(_03698_));
 sky130_fd_sc_hd__a21bo_1 _11116_ (.A1(_03611_),
    .A2(_03613_),
    .B1_N(_03612_),
    .X(_03699_));
 sky130_fd_sc_hd__nand3_1 _11117_ (.A(_03698_),
    .B(_03614_),
    .C(_03699_),
    .Y(_03700_));
 sky130_fd_sc_hd__a21o_1 _11118_ (.A1(_03614_),
    .A2(_03699_),
    .B1(_03698_),
    .X(_03701_));
 sky130_fd_sc_hd__and3_1 _11119_ (.A(_03697_),
    .B(_03700_),
    .C(_03701_),
    .X(_03702_));
 sky130_fd_sc_hd__a21oi_1 _11120_ (.A1(_03700_),
    .A2(_03701_),
    .B1(_03697_),
    .Y(_03703_));
 sky130_fd_sc_hd__nor4_2 _11121_ (.A(_03692_),
    .B(_03693_),
    .C(_03702_),
    .D(_03703_),
    .Y(_03704_));
 sky130_fd_sc_hd__or2_2 _11122_ (.A(_03692_),
    .B(_03704_),
    .X(_03705_));
 sky130_fd_sc_hd__xor2_2 _11123_ (.A(_03672_),
    .B(_03705_),
    .X(_03706_));
 sky130_fd_sc_hd__or3_1 _11124_ (.A(_03627_),
    .B(_03629_),
    .C(_03628_),
    .X(_03707_));
 sky130_fd_sc_hd__o21ai_1 _11125_ (.A1(_03629_),
    .A2(_03628_),
    .B1(_03627_),
    .Y(_03708_));
 sky130_fd_sc_hd__and2_1 _11126_ (.A(_02926_),
    .B(_03127_),
    .X(_03709_));
 sky130_fd_sc_hd__a22o_1 _11127_ (.A1(_03210_),
    .A2(_03247_),
    .B1(_03233_),
    .B2(_03208_),
    .X(_03710_));
 sky130_fd_sc_hd__nand4_1 _11128_ (.A(_02921_),
    .B(_02923_),
    .C(_03248_),
    .D(_03271_),
    .Y(_03711_));
 sky130_fd_sc_hd__a21bo_1 _11129_ (.A1(_03709_),
    .A2(_03710_),
    .B1_N(_03711_),
    .X(_03712_));
 sky130_fd_sc_hd__nand3_1 _11130_ (.A(_03707_),
    .B(_03708_),
    .C(_03712_),
    .Y(_03713_));
 sky130_fd_sc_hd__a21o_1 _11131_ (.A1(_03707_),
    .A2(_03708_),
    .B1(_03712_),
    .X(_03714_));
 sky130_fd_sc_hd__a22oi_1 _11132_ (.A1(_02897_),
    .A2(_03220_),
    .B1(_03040_),
    .B2(_02895_),
    .Y(_03715_));
 sky130_fd_sc_hd__and4_1 _11133_ (.A(_03634_),
    .B(_02897_),
    .C(_03220_),
    .D(_03039_),
    .X(_03716_));
 sky130_fd_sc_hd__or2_1 _11134_ (.A(_03715_),
    .B(_03716_),
    .X(_03717_));
 sky130_fd_sc_hd__xor2_1 _11135_ (.A(_02893_),
    .B(_03717_),
    .X(_03718_));
 sky130_fd_sc_hd__nand3_1 _11136_ (.A(_03713_),
    .B(_03714_),
    .C(_03718_),
    .Y(_03719_));
 sky130_fd_sc_hd__nand2_1 _11137_ (.A(_03713_),
    .B(_03719_),
    .Y(_03720_));
 sky130_fd_sc_hd__a21bo_1 _11138_ (.A1(_03697_),
    .A2(_03701_),
    .B1_N(_03700_),
    .X(_03721_));
 sky130_fd_sc_hd__o21bai_1 _11139_ (.A1(_03631_),
    .A2(_03632_),
    .B1_N(_03640_),
    .Y(_03722_));
 sky130_fd_sc_hd__and3_1 _11140_ (.A(_03721_),
    .B(_03641_),
    .C(_03722_),
    .X(_03723_));
 sky130_fd_sc_hd__a21oi_1 _11141_ (.A1(_03641_),
    .A2(_03722_),
    .B1(_03721_),
    .Y(_03724_));
 sky130_fd_sc_hd__or2_1 _11142_ (.A(_03723_),
    .B(_03724_),
    .X(_03725_));
 sky130_fd_sc_hd__xnor2_1 _11143_ (.A(_03720_),
    .B(_03725_),
    .Y(_03726_));
 sky130_fd_sc_hd__and2_1 _11144_ (.A(_03672_),
    .B(_03705_),
    .X(_03727_));
 sky130_fd_sc_hd__a21oi_1 _11145_ (.A1(_03706_),
    .A2(_03726_),
    .B1(_03727_),
    .Y(_03728_));
 sky130_fd_sc_hd__nor2_1 _11146_ (.A(_03671_),
    .B(_03728_),
    .Y(_03729_));
 sky130_fd_sc_hd__xor2_1 _11147_ (.A(_03671_),
    .B(_03728_),
    .X(_03730_));
 sky130_fd_sc_hd__and2b_1 _11148_ (.A_N(_03725_),
    .B(_03720_),
    .X(_03731_));
 sky130_fd_sc_hd__and2b_1 _11149_ (.A_N(_03659_),
    .B(_03658_),
    .X(_03732_));
 sky130_fd_sc_hd__xnor2_1 _11150_ (.A(_02911_),
    .B(_03732_),
    .Y(_03733_));
 sky130_fd_sc_hd__o21ai_1 _11151_ (.A1(_03723_),
    .A2(_03731_),
    .B1(_03733_),
    .Y(_03734_));
 sky130_fd_sc_hd__or3_1 _11152_ (.A(_03723_),
    .B(_03731_),
    .C(_03733_),
    .X(_03735_));
 sky130_fd_sc_hd__and2_1 _11153_ (.A(_03734_),
    .B(_03735_),
    .X(_03736_));
 sky130_fd_sc_hd__nor2_1 _11154_ (.A(_02893_),
    .B(_03717_),
    .Y(_03737_));
 sky130_fd_sc_hd__or3_1 _11155_ (.A(_02890_),
    .B(_03716_),
    .C(_03737_),
    .X(_03738_));
 sky130_fd_sc_hd__o21a_1 _11156_ (.A1(_03716_),
    .A2(_03737_),
    .B1(_02891_),
    .X(_03739_));
 sky130_fd_sc_hd__a31oi_2 _11157_ (.A1(_02909_),
    .A2(_02953_),
    .A3(_03738_),
    .B1(_03739_),
    .Y(_03740_));
 sky130_fd_sc_hd__xnor2_1 _11158_ (.A(_03736_),
    .B(_03740_),
    .Y(_03741_));
 sky130_fd_sc_hd__and2_1 _11159_ (.A(_03730_),
    .B(_03741_),
    .X(_03742_));
 sky130_fd_sc_hd__xor2_1 _11160_ (.A(_03649_),
    .B(_03661_),
    .X(_03743_));
 sky130_fd_sc_hd__o21ai_1 _11161_ (.A1(_03729_),
    .A2(_03742_),
    .B1(_03743_),
    .Y(_03744_));
 sky130_fd_sc_hd__or3_1 _11162_ (.A(_03743_),
    .B(_03729_),
    .C(_03742_),
    .X(_03745_));
 sky130_fd_sc_hd__nand2_1 _11163_ (.A(_03744_),
    .B(_03745_),
    .Y(_03746_));
 sky130_fd_sc_hd__or2b_1 _11164_ (.A(_03740_),
    .B_N(_03736_),
    .X(_03747_));
 sky130_fd_sc_hd__nand2_1 _11165_ (.A(_03734_),
    .B(_03747_),
    .Y(_03748_));
 sky130_fd_sc_hd__or2b_1 _11166_ (.A(_03746_),
    .B_N(_03748_),
    .X(_03749_));
 sky130_fd_sc_hd__xor2_1 _11167_ (.A(_03668_),
    .B(_03666_),
    .X(_03750_));
 sky130_fd_sc_hd__a21oi_2 _11168_ (.A1(_03744_),
    .A2(_03749_),
    .B1(_03750_),
    .Y(_03751_));
 sky130_fd_sc_hd__a21oi_1 _11169_ (.A1(_03664_),
    .A2(_03669_),
    .B1(_03592_),
    .Y(_03752_));
 sky130_fd_sc_hd__a21oi_1 _11170_ (.A1(_03670_),
    .A2(_03751_),
    .B1(_03752_),
    .Y(_03753_));
 sky130_fd_sc_hd__inv_2 _11171_ (.A(_03588_),
    .Y(_03754_));
 sky130_fd_sc_hd__o221a_1 _11172_ (.A1(_03507_),
    .A2(_03587_),
    .B1(_03591_),
    .B2(_03753_),
    .C1(_03754_),
    .X(_03755_));
 sky130_fd_sc_hd__buf_2 _11173_ (.A(\wfg_stim_mem_top.cfg_gain_q[23] ),
    .X(_03756_));
 sky130_fd_sc_hd__buf_2 _11174_ (.A(\wfg_stim_mem_top.cfg_gain_q[10] ),
    .X(_03757_));
 sky130_fd_sc_hd__and4_1 _11175_ (.A(_03756_),
    .B(_03757_),
    .C(net18),
    .D(net4),
    .X(_03758_));
 sky130_fd_sc_hd__clkbuf_4 _11176_ (.A(_03756_),
    .X(_03759_));
 sky130_fd_sc_hd__clkbuf_4 _11177_ (.A(net3),
    .X(_03760_));
 sky130_fd_sc_hd__nand4_1 _11178_ (.A(_03759_),
    .B(_03679_),
    .C(_03247_),
    .D(_03760_),
    .Y(_03761_));
 sky130_fd_sc_hd__clkbuf_4 _11179_ (.A(net4),
    .X(_03762_));
 sky130_fd_sc_hd__a22o_1 _11180_ (.A1(_03018_),
    .A2(net18),
    .B1(_03762_),
    .B2(_03013_),
    .X(_03763_));
 sky130_fd_sc_hd__or3b_1 _11181_ (.A(_03758_),
    .B(_03761_),
    .C_N(_03763_),
    .X(_03764_));
 sky130_fd_sc_hd__nand4_1 _11182_ (.A(_03759_),
    .B(_03596_),
    .C(_03127_),
    .D(_03762_),
    .Y(_03765_));
 sky130_fd_sc_hd__and4_1 _11183_ (.A(_03756_),
    .B(_03757_),
    .C(net17),
    .D(net3),
    .X(_03766_));
 sky130_fd_sc_hd__a21o_1 _11184_ (.A1(_03765_),
    .A2(_03763_),
    .B1(_03766_),
    .X(_03767_));
 sky130_fd_sc_hd__and2_1 _11185_ (.A(_02948_),
    .B(_03680_),
    .X(_03768_));
 sky130_fd_sc_hd__buf_4 _11186_ (.A(net6),
    .X(_03769_));
 sky130_fd_sc_hd__clkbuf_4 _11187_ (.A(net5),
    .X(_03770_));
 sky130_fd_sc_hd__buf_4 _11188_ (.A(_03770_),
    .X(_03771_));
 sky130_fd_sc_hd__nand4_1 _11189_ (.A(_02960_),
    .B(_02965_),
    .C(_03769_),
    .D(_03771_),
    .Y(_03772_));
 sky130_fd_sc_hd__clkbuf_4 _11190_ (.A(\wfg_stim_mem_top.cfg_gain_q[21] ),
    .X(_03773_));
 sky130_fd_sc_hd__clkbuf_4 _11191_ (.A(\wfg_stim_mem_top.cfg_gain_q[22] ),
    .X(_03774_));
 sky130_fd_sc_hd__a22o_1 _11192_ (.A1(_03773_),
    .A2(_03769_),
    .B1(_03770_),
    .B2(_03774_),
    .X(_03775_));
 sky130_fd_sc_hd__nand3_1 _11193_ (.A(_03768_),
    .B(_03772_),
    .C(_03775_),
    .Y(_03776_));
 sky130_fd_sc_hd__a21o_1 _11194_ (.A1(_03772_),
    .A2(_03775_),
    .B1(_03768_),
    .X(_03777_));
 sky130_fd_sc_hd__nand4_2 _11195_ (.A(_03764_),
    .B(_03767_),
    .C(_03776_),
    .D(_03777_),
    .Y(_03778_));
 sky130_fd_sc_hd__a22o_1 _11196_ (.A1(_03757_),
    .A2(net17),
    .B1(_03760_),
    .B2(_03756_),
    .X(_03779_));
 sky130_fd_sc_hd__and4_1 _11197_ (.A(_03756_),
    .B(_03757_),
    .C(net16),
    .D(net2),
    .X(_03780_));
 sky130_fd_sc_hd__a21o_1 _11198_ (.A1(_03761_),
    .A2(_03779_),
    .B1(_03780_),
    .X(_03781_));
 sky130_fd_sc_hd__nand2_1 _11199_ (.A(\wfg_stim_mem_top.cfg_gain_q[20] ),
    .B(_03769_),
    .Y(_03782_));
 sky130_fd_sc_hd__a22oi_2 _11200_ (.A1(_02954_),
    .A2(_03770_),
    .B1(_03762_),
    .B2(_02959_),
    .Y(_03783_));
 sky130_fd_sc_hd__and4_1 _11201_ (.A(_02959_),
    .B(_02954_),
    .C(net5),
    .D(net4),
    .X(_03784_));
 sky130_fd_sc_hd__or3_1 _11202_ (.A(_03782_),
    .B(_03783_),
    .C(_03784_),
    .X(_03785_));
 sky130_fd_sc_hd__o21ai_1 _11203_ (.A1(_03783_),
    .A2(_03784_),
    .B1(_03782_),
    .Y(_03786_));
 sky130_fd_sc_hd__and3_1 _11204_ (.A(_03761_),
    .B(_03780_),
    .C(_03779_),
    .X(_03787_));
 sky130_fd_sc_hd__a31o_1 _11205_ (.A1(_03781_),
    .A2(_03785_),
    .A3(_03786_),
    .B1(_03787_),
    .X(_03788_));
 sky130_fd_sc_hd__a22o_1 _11206_ (.A1(_03764_),
    .A2(_03767_),
    .B1(_03776_),
    .B2(_03777_),
    .X(_03789_));
 sky130_fd_sc_hd__nand3_4 _11207_ (.A(_03778_),
    .B(_03788_),
    .C(_03789_),
    .Y(_03790_));
 sky130_fd_sc_hd__a21o_1 _11208_ (.A1(_03778_),
    .A2(_03789_),
    .B1(_03788_),
    .X(_03791_));
 sky130_fd_sc_hd__and4_1 _11209_ (.A(_03143_),
    .B(\wfg_stim_mem_top.cfg_gain_q[18] ),
    .C(net8),
    .D(net7),
    .X(_03792_));
 sky130_fd_sc_hd__clkbuf_4 _11210_ (.A(net9),
    .X(_03793_));
 sky130_fd_sc_hd__nand2_1 _11211_ (.A(\wfg_stim_mem_top.cfg_gain_q[17] ),
    .B(_03793_),
    .Y(_03794_));
 sky130_fd_sc_hd__a22oi_1 _11212_ (.A1(_02937_),
    .A2(_03674_),
    .B1(_03680_),
    .B2(_03143_),
    .Y(_03795_));
 sky130_fd_sc_hd__or3_1 _11213_ (.A(_03792_),
    .B(_03794_),
    .C(_03795_),
    .X(_03796_));
 sky130_fd_sc_hd__or2b_1 _11214_ (.A(_03792_),
    .B_N(_03796_),
    .X(_03797_));
 sky130_fd_sc_hd__buf_4 _11215_ (.A(_02934_),
    .X(_03798_));
 sky130_fd_sc_hd__buf_4 _11216_ (.A(_03143_),
    .X(_03799_));
 sky130_fd_sc_hd__nand4_1 _11217_ (.A(_03799_),
    .B(_02940_),
    .C(_03793_),
    .D(_03674_),
    .Y(_03800_));
 sky130_fd_sc_hd__a22o_1 _11218_ (.A1(_02940_),
    .A2(_03793_),
    .B1(_03674_),
    .B2(_02943_),
    .X(_03801_));
 sky130_fd_sc_hd__nand4_1 _11219_ (.A(_03798_),
    .B(_03684_),
    .C(_03800_),
    .D(_03801_),
    .Y(_03802_));
 sky130_fd_sc_hd__o21bai_1 _11220_ (.A1(_03782_),
    .A2(_03783_),
    .B1_N(_03784_),
    .Y(_03803_));
 sky130_fd_sc_hd__a22o_1 _11221_ (.A1(_02934_),
    .A2(_03684_),
    .B1(_03800_),
    .B2(_03801_),
    .X(_03804_));
 sky130_fd_sc_hd__nand3_1 _11222_ (.A(_03802_),
    .B(_03803_),
    .C(_03804_),
    .Y(_03805_));
 sky130_fd_sc_hd__a21o_1 _11223_ (.A1(_03802_),
    .A2(_03804_),
    .B1(_03803_),
    .X(_03806_));
 sky130_fd_sc_hd__nand3_1 _11224_ (.A(_03797_),
    .B(_03805_),
    .C(_03806_),
    .Y(_03807_));
 sky130_fd_sc_hd__a21o_1 _11225_ (.A1(_03805_),
    .A2(_03806_),
    .B1(_03797_),
    .X(_03808_));
 sky130_fd_sc_hd__nand4_4 _11226_ (.A(_03790_),
    .B(_03791_),
    .C(_03807_),
    .D(_03808_),
    .Y(_03809_));
 sky130_fd_sc_hd__and4_1 _11227_ (.A(_03774_),
    .B(_03773_),
    .C(net7),
    .D(_03769_),
    .X(_03810_));
 sky130_fd_sc_hd__nand2_1 _11228_ (.A(_02948_),
    .B(_03597_),
    .Y(_03811_));
 sky130_fd_sc_hd__buf_4 _11229_ (.A(net6),
    .X(_03812_));
 sky130_fd_sc_hd__a22oi_2 _11230_ (.A1(_02965_),
    .A2(_03680_),
    .B1(_03812_),
    .B2(_02963_),
    .Y(_03813_));
 sky130_fd_sc_hd__or3_1 _11231_ (.A(_03810_),
    .B(_03811_),
    .C(_03813_),
    .X(_03814_));
 sky130_fd_sc_hd__and4_1 _11232_ (.A(_03678_),
    .B(_03679_),
    .C(net19),
    .D(_03770_),
    .X(_03815_));
 sky130_fd_sc_hd__a22o_1 _11233_ (.A1(_03596_),
    .A2(net19),
    .B1(_03770_),
    .B2(_03678_),
    .X(_03816_));
 sky130_fd_sc_hd__or3b_1 _11234_ (.A(_03765_),
    .B(_03815_),
    .C_N(_03816_),
    .X(_03817_));
 sky130_fd_sc_hd__nand4_2 _11235_ (.A(_03014_),
    .B(_03019_),
    .C(_03093_),
    .D(_03771_),
    .Y(_03818_));
 sky130_fd_sc_hd__a21o_1 _11236_ (.A1(_03818_),
    .A2(_03816_),
    .B1(_03758_),
    .X(_03819_));
 sky130_fd_sc_hd__o21ai_1 _11237_ (.A1(_03810_),
    .A2(_03813_),
    .B1(_03811_),
    .Y(_03820_));
 sky130_fd_sc_hd__nand4_1 _11238_ (.A(_03814_),
    .B(_03817_),
    .C(_03819_),
    .D(_03820_),
    .Y(_03821_));
 sky130_fd_sc_hd__and3_1 _11239_ (.A(_03765_),
    .B(_03766_),
    .C(_03763_),
    .X(_03822_));
 sky130_fd_sc_hd__a31o_1 _11240_ (.A1(_03767_),
    .A2(_03776_),
    .A3(_03777_),
    .B1(_03822_),
    .X(_03823_));
 sky130_fd_sc_hd__a22o_1 _11241_ (.A1(_03817_),
    .A2(_03819_),
    .B1(_03820_),
    .B2(_03814_),
    .X(_03824_));
 sky130_fd_sc_hd__nand3_1 _11242_ (.A(_03821_),
    .B(_03823_),
    .C(_03824_),
    .Y(_03825_));
 sky130_fd_sc_hd__a21o_1 _11243_ (.A1(_03821_),
    .A2(_03824_),
    .B1(_03823_),
    .X(_03826_));
 sky130_fd_sc_hd__nand2_1 _11244_ (.A(_03800_),
    .B(_03802_),
    .Y(_03827_));
 sky130_fd_sc_hd__and4_1 _11245_ (.A(_02943_),
    .B(_02940_),
    .C(_03436_),
    .D(net9),
    .X(_03828_));
 sky130_fd_sc_hd__nand2_1 _11246_ (.A(_02934_),
    .B(_03286_),
    .Y(_03829_));
 sky130_fd_sc_hd__buf_4 _11247_ (.A(_02937_),
    .X(_03830_));
 sky130_fd_sc_hd__a22oi_2 _11248_ (.A1(_03830_),
    .A2(_03436_),
    .B1(_03551_),
    .B2(_03799_),
    .Y(_03831_));
 sky130_fd_sc_hd__or3_1 _11249_ (.A(_03828_),
    .B(_03829_),
    .C(_03831_),
    .X(_03832_));
 sky130_fd_sc_hd__a21bo_1 _11250_ (.A1(_03768_),
    .A2(_03775_),
    .B1_N(_03772_),
    .X(_03833_));
 sky130_fd_sc_hd__o21ai_1 _11251_ (.A1(_03828_),
    .A2(_03831_),
    .B1(_03829_),
    .Y(_03834_));
 sky130_fd_sc_hd__nand3_1 _11252_ (.A(_03832_),
    .B(_03833_),
    .C(_03834_),
    .Y(_03835_));
 sky130_fd_sc_hd__a21o_1 _11253_ (.A1(_03832_),
    .A2(_03834_),
    .B1(_03833_),
    .X(_03836_));
 sky130_fd_sc_hd__nand3_1 _11254_ (.A(_03827_),
    .B(_03835_),
    .C(_03836_),
    .Y(_03837_));
 sky130_fd_sc_hd__a21o_1 _11255_ (.A1(_03835_),
    .A2(_03836_),
    .B1(_03827_),
    .X(_03838_));
 sky130_fd_sc_hd__a22oi_4 _11256_ (.A1(_03825_),
    .A2(_03826_),
    .B1(_03837_),
    .B2(_03838_),
    .Y(_03839_));
 sky130_fd_sc_hd__and4_2 _11257_ (.A(_03825_),
    .B(_03826_),
    .C(_03837_),
    .D(_03838_),
    .X(_03840_));
 sky130_fd_sc_hd__a211oi_4 _11258_ (.A1(_03790_),
    .A2(_03809_),
    .B1(_03839_),
    .C1(_03840_),
    .Y(_03841_));
 sky130_fd_sc_hd__o211a_1 _11259_ (.A1(_03840_),
    .A2(_03839_),
    .B1(_03809_),
    .C1(_03790_),
    .X(_03842_));
 sky130_fd_sc_hd__nand4_1 _11260_ (.A(_02920_),
    .B(_03212_),
    .C(_03279_),
    .D(_03286_),
    .Y(_03843_));
 sky130_fd_sc_hd__and2_1 _11261_ (.A(\wfg_stim_mem_top.cfg_gain_q[14] ),
    .B(_03230_),
    .X(_03844_));
 sky130_fd_sc_hd__a22o_1 _11262_ (.A1(_03209_),
    .A2(_03279_),
    .B1(_03286_),
    .B2(_02919_),
    .X(_03845_));
 sky130_fd_sc_hd__nand3_1 _11263_ (.A(_03843_),
    .B(_03844_),
    .C(_03845_),
    .Y(_03846_));
 sky130_fd_sc_hd__nand2_1 _11264_ (.A(\wfg_stim_mem_top.cfg_gain_q[14] ),
    .B(_03279_),
    .Y(_03847_));
 sky130_fd_sc_hd__a22oi_2 _11265_ (.A1(_03212_),
    .A2(_03286_),
    .B1(_03436_),
    .B2(_03217_),
    .Y(_03848_));
 sky130_fd_sc_hd__and4_1 _11266_ (.A(_02919_),
    .B(_03209_),
    .C(net11),
    .D(net10),
    .X(_03849_));
 sky130_fd_sc_hd__o21bai_1 _11267_ (.A1(_03847_),
    .A2(_03848_),
    .B1_N(_03849_),
    .Y(_03850_));
 sky130_fd_sc_hd__a22o_1 _11268_ (.A1(_02926_),
    .A2(_03236_),
    .B1(_03843_),
    .B2(_03845_),
    .X(_03851_));
 sky130_fd_sc_hd__nand3_1 _11269_ (.A(_03846_),
    .B(_03850_),
    .C(_03851_),
    .Y(_03852_));
 sky130_fd_sc_hd__a21o_1 _11270_ (.A1(_03846_),
    .A2(_03851_),
    .B1(_03850_),
    .X(_03853_));
 sky130_fd_sc_hd__nand2_1 _11271_ (.A(_02892_),
    .B(_03094_),
    .Y(_03854_));
 sky130_fd_sc_hd__a22oi_1 _11272_ (.A1(_03637_),
    .A2(_03233_),
    .B1(_03228_),
    .B2(_03636_),
    .Y(_03855_));
 sky130_fd_sc_hd__and4_1 _11273_ (.A(\wfg_stim_mem_top.cfg_gain_q[13] ),
    .B(\wfg_stim_mem_top.cfg_gain_q[12] ),
    .C(_03233_),
    .D(_03228_),
    .X(_03856_));
 sky130_fd_sc_hd__nor2_1 _11274_ (.A(_03855_),
    .B(_03856_),
    .Y(_03857_));
 sky130_fd_sc_hd__xnor2_2 _11275_ (.A(_03854_),
    .B(_03857_),
    .Y(_03858_));
 sky130_fd_sc_hd__nand3_1 _11276_ (.A(_03852_),
    .B(_03853_),
    .C(_03858_),
    .Y(_03859_));
 sky130_fd_sc_hd__nand2_1 _11277_ (.A(_03852_),
    .B(_03859_),
    .Y(_03860_));
 sky130_fd_sc_hd__and4_1 _11278_ (.A(_03532_),
    .B(_02922_),
    .C(_03230_),
    .D(_03279_),
    .X(_03861_));
 sky130_fd_sc_hd__nand2_1 _11279_ (.A(_02926_),
    .B(_03228_),
    .Y(_03862_));
 sky130_fd_sc_hd__a22oi_2 _11280_ (.A1(_03210_),
    .A2(_03230_),
    .B1(_03280_),
    .B2(_03208_),
    .Y(_03863_));
 sky130_fd_sc_hd__or3_1 _11281_ (.A(_03861_),
    .B(_03862_),
    .C(_03863_),
    .X(_03864_));
 sky130_fd_sc_hd__a21bo_1 _11282_ (.A1(_03844_),
    .A2(_03845_),
    .B1_N(_03843_),
    .X(_03865_));
 sky130_fd_sc_hd__o21ai_1 _11283_ (.A1(_03861_),
    .A2(_03863_),
    .B1(_03862_),
    .Y(_03866_));
 sky130_fd_sc_hd__nand3_1 _11284_ (.A(_03864_),
    .B(_03865_),
    .C(_03866_),
    .Y(_03867_));
 sky130_fd_sc_hd__a21o_1 _11285_ (.A1(_03864_),
    .A2(_03866_),
    .B1(_03865_),
    .X(_03868_));
 sky130_fd_sc_hd__buf_4 _11286_ (.A(_02892_),
    .X(_03869_));
 sky130_fd_sc_hd__nand2_1 _11287_ (.A(_03869_),
    .B(_03040_),
    .Y(_03870_));
 sky130_fd_sc_hd__a22oi_1 _11288_ (.A1(_02897_),
    .A2(_03248_),
    .B1(_03234_),
    .B2(_03634_),
    .Y(_03871_));
 sky130_fd_sc_hd__buf_4 _11289_ (.A(\wfg_stim_mem_top.cfg_gain_q[13] ),
    .X(_03872_));
 sky130_fd_sc_hd__buf_4 _11290_ (.A(\wfg_stim_mem_top.cfg_gain_q[12] ),
    .X(_03873_));
 sky130_fd_sc_hd__and4_1 _11291_ (.A(_03872_),
    .B(_03873_),
    .C(_03247_),
    .D(_03271_),
    .X(_03874_));
 sky130_fd_sc_hd__nor2_1 _11292_ (.A(_03871_),
    .B(_03874_),
    .Y(_03875_));
 sky130_fd_sc_hd__xnor2_2 _11293_ (.A(_03870_),
    .B(_03875_),
    .Y(_03876_));
 sky130_fd_sc_hd__nand3_1 _11294_ (.A(_03867_),
    .B(_03868_),
    .C(_03876_),
    .Y(_03877_));
 sky130_fd_sc_hd__a21bo_1 _11295_ (.A1(_03797_),
    .A2(_03806_),
    .B1_N(_03805_),
    .X(_03878_));
 sky130_fd_sc_hd__a21o_1 _11296_ (.A1(_03867_),
    .A2(_03868_),
    .B1(_03876_),
    .X(_03879_));
 sky130_fd_sc_hd__nand3_1 _11297_ (.A(_03877_),
    .B(_03878_),
    .C(_03879_),
    .Y(_03880_));
 sky130_fd_sc_hd__a21o_1 _11298_ (.A1(_03877_),
    .A2(_03879_),
    .B1(_03878_),
    .X(_03881_));
 sky130_fd_sc_hd__and3_1 _11299_ (.A(_03860_),
    .B(_03880_),
    .C(_03881_),
    .X(_03882_));
 sky130_fd_sc_hd__a21oi_2 _11300_ (.A1(_03880_),
    .A2(_03881_),
    .B1(_03860_),
    .Y(_03883_));
 sky130_fd_sc_hd__nor4_4 _11301_ (.A(_03841_),
    .B(_03842_),
    .C(_03882_),
    .D(_03883_),
    .Y(_03884_));
 sky130_fd_sc_hd__and3_2 _11302_ (.A(_03821_),
    .B(_03823_),
    .C(_03824_),
    .X(_03885_));
 sky130_fd_sc_hd__and3_1 _11303_ (.A(_03758_),
    .B(_03818_),
    .C(_03816_),
    .X(_03886_));
 sky130_fd_sc_hd__a31o_1 _11304_ (.A1(_03814_),
    .A2(_03819_),
    .A3(_03820_),
    .B1(_03886_),
    .X(_03887_));
 sky130_fd_sc_hd__and4_1 _11305_ (.A(_03759_),
    .B(_03596_),
    .C(net20),
    .D(_03769_),
    .X(_03888_));
 sky130_fd_sc_hd__a22o_1 _11306_ (.A1(_03596_),
    .A2(net20),
    .B1(_03812_),
    .B2(_03759_),
    .X(_03889_));
 sky130_fd_sc_hd__or3b_1 _11307_ (.A(_03818_),
    .B(_03888_),
    .C_N(_03889_),
    .X(_03890_));
 sky130_fd_sc_hd__nand4_1 _11308_ (.A(_03014_),
    .B(_03019_),
    .C(_03038_),
    .D(_03812_),
    .Y(_03891_));
 sky130_fd_sc_hd__a21o_1 _11309_ (.A1(_03891_),
    .A2(_03889_),
    .B1(_03815_),
    .X(_03892_));
 sky130_fd_sc_hd__and2_1 _11310_ (.A(_02948_),
    .B(_03551_),
    .X(_03893_));
 sky130_fd_sc_hd__buf_4 _11311_ (.A(net7),
    .X(_03894_));
 sky130_fd_sc_hd__a22o_1 _11312_ (.A1(_02955_),
    .A2(_03597_),
    .B1(_03894_),
    .B2(_02960_),
    .X(_03895_));
 sky130_fd_sc_hd__nand4_1 _11313_ (.A(_02960_),
    .B(_02955_),
    .C(_03597_),
    .D(_03894_),
    .Y(_03896_));
 sky130_fd_sc_hd__nand3_1 _11314_ (.A(_03893_),
    .B(_03895_),
    .C(_03896_),
    .Y(_03897_));
 sky130_fd_sc_hd__a21o_1 _11315_ (.A1(_03895_),
    .A2(_03896_),
    .B1(_03893_),
    .X(_03898_));
 sky130_fd_sc_hd__nand4_2 _11316_ (.A(_03890_),
    .B(_03892_),
    .C(_03897_),
    .D(_03898_),
    .Y(_03899_));
 sky130_fd_sc_hd__a22o_1 _11317_ (.A1(_03890_),
    .A2(_03892_),
    .B1(_03897_),
    .B2(_03898_),
    .X(_03900_));
 sky130_fd_sc_hd__nand3_4 _11318_ (.A(_03887_),
    .B(_03899_),
    .C(_03900_),
    .Y(_03901_));
 sky130_fd_sc_hd__a21o_1 _11319_ (.A1(_03899_),
    .A2(_03900_),
    .B1(_03887_),
    .X(_03902_));
 sky130_fd_sc_hd__o21bai_1 _11320_ (.A1(_03811_),
    .A2(_03813_),
    .B1_N(_03810_),
    .Y(_03903_));
 sky130_fd_sc_hd__nand4_2 _11321_ (.A(_02944_),
    .B(_02941_),
    .C(_03287_),
    .D(_03684_),
    .Y(_03904_));
 sky130_fd_sc_hd__a22o_1 _11322_ (.A1(_02938_),
    .A2(_03286_),
    .B1(_03684_),
    .B2(_03144_),
    .X(_03905_));
 sky130_fd_sc_hd__nand4_2 _11323_ (.A(_02935_),
    .B(_03281_),
    .C(_03904_),
    .D(_03905_),
    .Y(_03906_));
 sky130_fd_sc_hd__a22o_1 _11324_ (.A1(_02935_),
    .A2(_03280_),
    .B1(_03904_),
    .B2(_03905_),
    .X(_03907_));
 sky130_fd_sc_hd__nand3_1 _11325_ (.A(_03903_),
    .B(_03906_),
    .C(_03907_),
    .Y(_03908_));
 sky130_fd_sc_hd__a21o_1 _11326_ (.A1(_03906_),
    .A2(_03907_),
    .B1(_03903_),
    .X(_03909_));
 sky130_fd_sc_hd__or2b_1 _11327_ (.A(_03828_),
    .B_N(_03832_),
    .X(_03910_));
 sky130_fd_sc_hd__a21o_1 _11328_ (.A1(_03908_),
    .A2(_03909_),
    .B1(_03910_),
    .X(_03911_));
 sky130_fd_sc_hd__nand3_1 _11329_ (.A(_03908_),
    .B(_03910_),
    .C(_03909_),
    .Y(_03912_));
 sky130_fd_sc_hd__a22o_1 _11330_ (.A1(_03901_),
    .A2(_03902_),
    .B1(_03911_),
    .B2(_03912_),
    .X(_03913_));
 sky130_fd_sc_hd__nand4_4 _11331_ (.A(_03912_),
    .B(_03901_),
    .C(_03902_),
    .D(_03911_),
    .Y(_03914_));
 sky130_fd_sc_hd__o211a_1 _11332_ (.A1(_03885_),
    .A2(_03840_),
    .B1(_03913_),
    .C1(_03914_),
    .X(_03915_));
 sky130_fd_sc_hd__a211oi_2 _11333_ (.A1(_03914_),
    .A2(_03913_),
    .B1(_03840_),
    .C1(_03885_),
    .Y(_03916_));
 sky130_fd_sc_hd__and2_1 _11334_ (.A(_03867_),
    .B(_03877_),
    .X(_03917_));
 sky130_fd_sc_hd__nand4_1 _11335_ (.A(_03218_),
    .B(_03210_),
    .C(_03228_),
    .D(_03236_),
    .Y(_03918_));
 sky130_fd_sc_hd__and2_1 _11336_ (.A(_02926_),
    .B(_03233_),
    .X(_03919_));
 sky130_fd_sc_hd__a22o_1 _11337_ (.A1(_03531_),
    .A2(_03228_),
    .B1(_03230_),
    .B2(_03532_),
    .X(_03920_));
 sky130_fd_sc_hd__nand3_1 _11338_ (.A(_03918_),
    .B(_03919_),
    .C(_03920_),
    .Y(_03921_));
 sky130_fd_sc_hd__a22o_1 _11339_ (.A1(_02917_),
    .A2(_03271_),
    .B1(_03918_),
    .B2(_03920_),
    .X(_03922_));
 sky130_fd_sc_hd__o21bai_1 _11340_ (.A1(_03862_),
    .A2(_03863_),
    .B1_N(_03861_),
    .Y(_03923_));
 sky130_fd_sc_hd__nand3_1 _11341_ (.A(_03921_),
    .B(_03922_),
    .C(_03923_),
    .Y(_03924_));
 sky130_fd_sc_hd__a21o_1 _11342_ (.A1(_03921_),
    .A2(_03922_),
    .B1(_03923_),
    .X(_03925_));
 sky130_fd_sc_hd__nand2_2 _11343_ (.A(_03490_),
    .B(_03220_),
    .Y(_03926_));
 sky130_fd_sc_hd__a22oi_1 _11344_ (.A1(_02900_),
    .A2(_03128_),
    .B1(_03248_),
    .B2(_03872_),
    .Y(_03927_));
 sky130_fd_sc_hd__and4_1 _11345_ (.A(_02894_),
    .B(_02896_),
    .C(_03127_),
    .D(_03247_),
    .X(_03928_));
 sky130_fd_sc_hd__nor2_2 _11346_ (.A(_03927_),
    .B(_03928_),
    .Y(_03929_));
 sky130_fd_sc_hd__xnor2_4 _11347_ (.A(_03926_),
    .B(_03929_),
    .Y(_03930_));
 sky130_fd_sc_hd__nand3_1 _11348_ (.A(_03924_),
    .B(_03925_),
    .C(_03930_),
    .Y(_03931_));
 sky130_fd_sc_hd__a21bo_1 _11349_ (.A1(_03827_),
    .A2(_03836_),
    .B1_N(_03835_),
    .X(_03932_));
 sky130_fd_sc_hd__a21o_1 _11350_ (.A1(_03924_),
    .A2(_03925_),
    .B1(_03930_),
    .X(_03933_));
 sky130_fd_sc_hd__and3_1 _11351_ (.A(_03931_),
    .B(_03932_),
    .C(_03933_),
    .X(_03934_));
 sky130_fd_sc_hd__a21oi_1 _11352_ (.A1(_03931_),
    .A2(_03933_),
    .B1(_03932_),
    .Y(_03935_));
 sky130_fd_sc_hd__nor3_2 _11353_ (.A(_03917_),
    .B(_03934_),
    .C(_03935_),
    .Y(_03936_));
 sky130_fd_sc_hd__o21a_1 _11354_ (.A1(_03934_),
    .A2(_03935_),
    .B1(_03917_),
    .X(_03937_));
 sky130_fd_sc_hd__o22ai_4 _11355_ (.A1(_03915_),
    .A2(_03916_),
    .B1(_03936_),
    .B2(_03937_),
    .Y(_03938_));
 sky130_fd_sc_hd__or4_4 _11356_ (.A(_03915_),
    .B(_03916_),
    .C(_03936_),
    .D(_03937_),
    .X(_03939_));
 sky130_fd_sc_hd__o211a_2 _11357_ (.A1(_03841_),
    .A2(_03884_),
    .B1(_03938_),
    .C1(_03939_),
    .X(_03940_));
 sky130_fd_sc_hd__a211oi_4 _11358_ (.A1(_03939_),
    .A2(_03938_),
    .B1(_03884_),
    .C1(_03841_),
    .Y(_03941_));
 sky130_fd_sc_hd__buf_6 _11359_ (.A(_02887_),
    .X(_03942_));
 sky130_fd_sc_hd__clkbuf_8 _11360_ (.A(_03942_),
    .X(_03943_));
 sky130_fd_sc_hd__buf_4 _11361_ (.A(_03943_),
    .X(_03944_));
 sky130_fd_sc_hd__buf_4 _11362_ (.A(_03869_),
    .X(_03945_));
 sky130_fd_sc_hd__a31o_1 _11363_ (.A1(_03945_),
    .A2(_03095_),
    .A3(_03857_),
    .B1(_03856_),
    .X(_03946_));
 sky130_fd_sc_hd__buf_4 _11364_ (.A(_02906_),
    .X(_03947_));
 sky130_fd_sc_hd__buf_4 _11365_ (.A(_02886_),
    .X(_03948_));
 sky130_fd_sc_hd__nand2_1 _11366_ (.A(_03948_),
    .B(_03029_),
    .Y(_03949_));
 sky130_fd_sc_hd__xnor2_1 _11367_ (.A(_03946_),
    .B(_03949_),
    .Y(_03950_));
 sky130_fd_sc_hd__and3_1 _11368_ (.A(_03947_),
    .B(_03129_),
    .C(_03950_),
    .X(_03951_));
 sky130_fd_sc_hd__a31o_1 _11369_ (.A1(_03944_),
    .A2(_03029_),
    .A3(_03946_),
    .B1(_03951_),
    .X(_03952_));
 sky130_fd_sc_hd__a21boi_2 _11370_ (.A1(_03860_),
    .A2(_03881_),
    .B1_N(_03880_),
    .Y(_03953_));
 sky130_fd_sc_hd__buf_4 _11371_ (.A(_02907_),
    .X(_03954_));
 sky130_fd_sc_hd__a31o_1 _11372_ (.A1(_03945_),
    .A2(_03040_),
    .A3(_03875_),
    .B1(_03874_),
    .X(_03955_));
 sky130_fd_sc_hd__nand2_1 _11373_ (.A(_03948_),
    .B(_03022_),
    .Y(_03956_));
 sky130_fd_sc_hd__xnor2_1 _11374_ (.A(_03955_),
    .B(_03956_),
    .Y(_03957_));
 sky130_fd_sc_hd__and3_1 _11375_ (.A(_03954_),
    .B(_03095_),
    .C(_03957_),
    .X(_03958_));
 sky130_fd_sc_hd__buf_6 _11376_ (.A(_02907_),
    .X(_03959_));
 sky130_fd_sc_hd__a21oi_1 _11377_ (.A1(_03959_),
    .A2(_03095_),
    .B1(_03957_),
    .Y(_03960_));
 sky130_fd_sc_hd__nor2_1 _11378_ (.A(_03958_),
    .B(_03960_),
    .Y(_03961_));
 sky130_fd_sc_hd__xnor2_1 _11379_ (.A(_03953_),
    .B(_03961_),
    .Y(_03962_));
 sky130_fd_sc_hd__xnor2_2 _11380_ (.A(_03952_),
    .B(_03962_),
    .Y(_03963_));
 sky130_fd_sc_hd__nor3_1 _11381_ (.A(_03940_),
    .B(_03941_),
    .C(_03963_),
    .Y(_03964_));
 sky130_fd_sc_hd__o211ai_4 _11382_ (.A1(_03885_),
    .A2(_03840_),
    .B1(_03913_),
    .C1(_03914_),
    .Y(_03965_));
 sky130_fd_sc_hd__a22o_1 _11383_ (.A1(_03596_),
    .A2(net21),
    .B1(_03894_),
    .B2(_03759_),
    .X(_03966_));
 sky130_fd_sc_hd__or3b_1 _11384_ (.A(_03891_),
    .B(_03681_),
    .C_N(_03966_),
    .X(_03967_));
 sky130_fd_sc_hd__nand4_2 _11385_ (.A(_03014_),
    .B(_03019_),
    .C(_02958_),
    .D(_03894_),
    .Y(_03968_));
 sky130_fd_sc_hd__a21o_1 _11386_ (.A1(_03968_),
    .A2(_03966_),
    .B1(_03888_),
    .X(_03969_));
 sky130_fd_sc_hd__nand2_1 _11387_ (.A(_02948_),
    .B(_03436_),
    .Y(_03970_));
 sky130_fd_sc_hd__a22oi_2 _11388_ (.A1(_02965_),
    .A2(_03793_),
    .B1(_03597_),
    .B2(_02960_),
    .Y(_03971_));
 sky130_fd_sc_hd__and4_1 _11389_ (.A(_02963_),
    .B(_02965_),
    .C(_03793_),
    .D(_03674_),
    .X(_03972_));
 sky130_fd_sc_hd__or3_1 _11390_ (.A(_03970_),
    .B(_03971_),
    .C(_03972_),
    .X(_03973_));
 sky130_fd_sc_hd__o21ai_1 _11391_ (.A1(_03971_),
    .A2(_03972_),
    .B1(_03970_),
    .Y(_03974_));
 sky130_fd_sc_hd__nand4_1 _11392_ (.A(_03967_),
    .B(_03969_),
    .C(_03973_),
    .D(_03974_),
    .Y(_03975_));
 sky130_fd_sc_hd__a22o_1 _11393_ (.A1(_03967_),
    .A2(_03969_),
    .B1(_03973_),
    .B2(_03974_),
    .X(_03976_));
 sky130_fd_sc_hd__and3_1 _11394_ (.A(_03815_),
    .B(_03891_),
    .C(_03889_),
    .X(_03977_));
 sky130_fd_sc_hd__a31o_1 _11395_ (.A1(_03892_),
    .A2(_03897_),
    .A3(_03898_),
    .B1(_03977_),
    .X(_03978_));
 sky130_fd_sc_hd__and3_2 _11396_ (.A(_03975_),
    .B(_03976_),
    .C(_03978_),
    .X(_03979_));
 sky130_fd_sc_hd__a21oi_2 _11397_ (.A1(_03975_),
    .A2(_03976_),
    .B1(_03978_),
    .Y(_03980_));
 sky130_fd_sc_hd__nand2_1 _11398_ (.A(_03904_),
    .B(_03906_),
    .Y(_03981_));
 sky130_fd_sc_hd__a21bo_1 _11399_ (.A1(_03893_),
    .A2(_03895_),
    .B1_N(_03896_),
    .X(_03982_));
 sky130_fd_sc_hd__nand2_1 _11400_ (.A(_03798_),
    .B(_03236_),
    .Y(_03983_));
 sky130_fd_sc_hd__nand4_1 _11401_ (.A(_02944_),
    .B(_02938_),
    .C(_03280_),
    .D(_03287_),
    .Y(_03984_));
 sky130_fd_sc_hd__a22o_1 _11402_ (.A1(_02938_),
    .A2(_03279_),
    .B1(_03287_),
    .B2(_03144_),
    .X(_03985_));
 sky130_fd_sc_hd__nand3b_1 _11403_ (.A_N(_03983_),
    .B(_03984_),
    .C(_03985_),
    .Y(_03986_));
 sky130_fd_sc_hd__a21bo_1 _11404_ (.A1(_03984_),
    .A2(_03985_),
    .B1_N(_03983_),
    .X(_03987_));
 sky130_fd_sc_hd__nand3_1 _11405_ (.A(_03982_),
    .B(_03986_),
    .C(_03987_),
    .Y(_03988_));
 sky130_fd_sc_hd__a21o_1 _11406_ (.A1(_03986_),
    .A2(_03987_),
    .B1(_03982_),
    .X(_03989_));
 sky130_fd_sc_hd__and3_1 _11407_ (.A(_03981_),
    .B(_03988_),
    .C(_03989_),
    .X(_03990_));
 sky130_fd_sc_hd__a21oi_2 _11408_ (.A1(_03988_),
    .A2(_03989_),
    .B1(_03981_),
    .Y(_03991_));
 sky130_fd_sc_hd__nor4_4 _11409_ (.A(_03979_),
    .B(_03980_),
    .C(_03990_),
    .D(_03991_),
    .Y(_03992_));
 sky130_fd_sc_hd__o22a_1 _11410_ (.A1(_03979_),
    .A2(_03980_),
    .B1(_03990_),
    .B2(_03991_),
    .X(_03993_));
 sky130_fd_sc_hd__a211oi_4 _11411_ (.A1(_03901_),
    .A2(_03914_),
    .B1(_03992_),
    .C1(_03993_),
    .Y(_03994_));
 sky130_fd_sc_hd__o211a_1 _11412_ (.A1(_03992_),
    .A2(_03993_),
    .B1(_03901_),
    .C1(_03914_),
    .X(_03995_));
 sky130_fd_sc_hd__a21bo_1 _11413_ (.A1(_03910_),
    .A2(_03909_),
    .B1_N(_03908_),
    .X(_03996_));
 sky130_fd_sc_hd__nand2_1 _11414_ (.A(_02917_),
    .B(_03248_),
    .Y(_03997_));
 sky130_fd_sc_hd__and4_1 _11415_ (.A(_03208_),
    .B(_03210_),
    .C(_03233_),
    .D(_03228_),
    .X(_03998_));
 sky130_fd_sc_hd__a22oi_2 _11416_ (.A1(_03213_),
    .A2(_03233_),
    .B1(_03229_),
    .B2(_03218_),
    .Y(_03999_));
 sky130_fd_sc_hd__or3_1 _11417_ (.A(_03997_),
    .B(_03998_),
    .C(_03999_),
    .X(_04000_));
 sky130_fd_sc_hd__o21ai_1 _11418_ (.A1(_03998_),
    .A2(_03999_),
    .B1(_03997_),
    .Y(_04001_));
 sky130_fd_sc_hd__a21bo_1 _11419_ (.A1(_03919_),
    .A2(_03920_),
    .B1_N(_03918_),
    .X(_04002_));
 sky130_fd_sc_hd__nand3_2 _11420_ (.A(_04000_),
    .B(_04001_),
    .C(_04002_),
    .Y(_04003_));
 sky130_fd_sc_hd__a21o_1 _11421_ (.A1(_04000_),
    .A2(_04001_),
    .B1(_04002_),
    .X(_04004_));
 sky130_fd_sc_hd__nand2_2 _11422_ (.A(_03869_),
    .B(_02987_),
    .Y(_04005_));
 sky130_fd_sc_hd__a22oi_1 _11423_ (.A1(_02900_),
    .A2(_03094_),
    .B1(_03128_),
    .B2(_03634_),
    .Y(_04006_));
 sky130_fd_sc_hd__and4_1 _11424_ (.A(_02894_),
    .B(_02896_),
    .C(_03093_),
    .D(_03127_),
    .X(_04007_));
 sky130_fd_sc_hd__or2_2 _11425_ (.A(_04006_),
    .B(_04007_),
    .X(_04008_));
 sky130_fd_sc_hd__xor2_4 _11426_ (.A(_04005_),
    .B(_04008_),
    .X(_04009_));
 sky130_fd_sc_hd__nand3_2 _11427_ (.A(_04003_),
    .B(_04004_),
    .C(_04009_),
    .Y(_04010_));
 sky130_fd_sc_hd__a21o_1 _11428_ (.A1(_04003_),
    .A2(_04004_),
    .B1(_04009_),
    .X(_04011_));
 sky130_fd_sc_hd__nand3_1 _11429_ (.A(_03996_),
    .B(_04010_),
    .C(_04011_),
    .Y(_04012_));
 sky130_fd_sc_hd__a21o_1 _11430_ (.A1(_04010_),
    .A2(_04011_),
    .B1(_03996_),
    .X(_04013_));
 sky130_fd_sc_hd__nand2_1 _11431_ (.A(_03924_),
    .B(_03931_),
    .Y(_04014_));
 sky130_fd_sc_hd__a21oi_2 _11432_ (.A1(_04012_),
    .A2(_04013_),
    .B1(_04014_),
    .Y(_04015_));
 sky130_fd_sc_hd__and3_1 _11433_ (.A(_04012_),
    .B(_04014_),
    .C(_04013_),
    .X(_04016_));
 sky130_fd_sc_hd__o22a_1 _11434_ (.A1(_03994_),
    .A2(_03995_),
    .B1(_04015_),
    .B2(_04016_),
    .X(_04017_));
 sky130_fd_sc_hd__nor4_4 _11435_ (.A(_04016_),
    .B(_03994_),
    .C(_03995_),
    .D(_04015_),
    .Y(_04018_));
 sky130_fd_sc_hd__a211oi_4 _11436_ (.A1(_03965_),
    .A2(_03939_),
    .B1(_04017_),
    .C1(_04018_),
    .Y(_04019_));
 sky130_fd_sc_hd__o211a_1 _11437_ (.A1(_04018_),
    .A2(_04017_),
    .B1(_03939_),
    .C1(_03965_),
    .X(_04020_));
 sky130_fd_sc_hd__a31o_1 _11438_ (.A1(_03944_),
    .A2(_03022_),
    .A3(_03955_),
    .B1(_03958_),
    .X(_04021_));
 sky130_fd_sc_hd__o21ba_1 _11439_ (.A1(_03917_),
    .A2(_03935_),
    .B1_N(_03934_),
    .X(_04022_));
 sky130_fd_sc_hd__a31o_1 _11440_ (.A1(_03945_),
    .A2(_03029_),
    .A3(_03929_),
    .B1(_03928_),
    .X(_04023_));
 sky130_fd_sc_hd__nand2_1 _11441_ (.A(_03942_),
    .B(_02953_),
    .Y(_04024_));
 sky130_fd_sc_hd__xnor2_1 _11442_ (.A(_04023_),
    .B(_04024_),
    .Y(_04025_));
 sky130_fd_sc_hd__and3_1 _11443_ (.A(_03954_),
    .B(_03040_),
    .C(_04025_),
    .X(_04026_));
 sky130_fd_sc_hd__a21oi_1 _11444_ (.A1(_03959_),
    .A2(_03040_),
    .B1(_04025_),
    .Y(_04027_));
 sky130_fd_sc_hd__nor2_1 _11445_ (.A(_04026_),
    .B(_04027_),
    .Y(_04028_));
 sky130_fd_sc_hd__xnor2_1 _11446_ (.A(_04022_),
    .B(_04028_),
    .Y(_04029_));
 sky130_fd_sc_hd__xnor2_1 _11447_ (.A(_04021_),
    .B(_04029_),
    .Y(_04030_));
 sky130_fd_sc_hd__o21ai_1 _11448_ (.A1(_04019_),
    .A2(_04020_),
    .B1(_04030_),
    .Y(_04031_));
 sky130_fd_sc_hd__or3_1 _11449_ (.A(_04019_),
    .B(_04020_),
    .C(_04030_),
    .X(_04032_));
 sky130_fd_sc_hd__o211a_1 _11450_ (.A1(_03940_),
    .A2(_03964_),
    .B1(_04031_),
    .C1(_04032_),
    .X(_04033_));
 sky130_fd_sc_hd__inv_2 _11451_ (.A(_04033_),
    .Y(_04034_));
 sky130_fd_sc_hd__or3_1 _11452_ (.A(_03958_),
    .B(_03953_),
    .C(_03960_),
    .X(_04035_));
 sky130_fd_sc_hd__nand2_1 _11453_ (.A(_03952_),
    .B(_03962_),
    .Y(_04036_));
 sky130_fd_sc_hd__a211oi_2 _11454_ (.A1(_04032_),
    .A2(_04031_),
    .B1(_03964_),
    .C1(_03940_),
    .Y(_04037_));
 sky130_fd_sc_hd__a211o_1 _11455_ (.A1(_04035_),
    .A2(_04036_),
    .B1(_04033_),
    .C1(_04037_),
    .X(_04038_));
 sky130_fd_sc_hd__or3_1 _11456_ (.A(_04026_),
    .B(_04022_),
    .C(_04027_),
    .X(_04039_));
 sky130_fd_sc_hd__nand2_1 _11457_ (.A(_04021_),
    .B(_04029_),
    .Y(_04040_));
 sky130_fd_sc_hd__nor3_1 _11458_ (.A(_04019_),
    .B(_04020_),
    .C(_04030_),
    .Y(_04041_));
 sky130_fd_sc_hd__or3b_1 _11459_ (.A(_03968_),
    .B(_03598_),
    .C_N(_03677_),
    .X(_04042_));
 sky130_fd_sc_hd__nand4_1 _11460_ (.A(_04042_),
    .B(_03682_),
    .C(_03688_),
    .D(_03689_),
    .Y(_04043_));
 sky130_fd_sc_hd__a22o_1 _11461_ (.A1(_04042_),
    .A2(_03682_),
    .B1(_03688_),
    .B2(_03689_),
    .X(_04044_));
 sky130_fd_sc_hd__and3_1 _11462_ (.A(_03888_),
    .B(_03968_),
    .C(_03966_),
    .X(_04045_));
 sky130_fd_sc_hd__a31o_1 _11463_ (.A1(_03969_),
    .A2(_03973_),
    .A3(_03974_),
    .B1(_04045_),
    .X(_04046_));
 sky130_fd_sc_hd__nand3_2 _11464_ (.A(_04043_),
    .B(_04044_),
    .C(_04046_),
    .Y(_04047_));
 sky130_fd_sc_hd__a21o_1 _11465_ (.A1(_04043_),
    .A2(_04044_),
    .B1(_04046_),
    .X(_04048_));
 sky130_fd_sc_hd__nand2_1 _11466_ (.A(_03984_),
    .B(_03986_),
    .Y(_04049_));
 sky130_fd_sc_hd__o21bai_2 _11467_ (.A1(_03970_),
    .A2(_03971_),
    .B1_N(_03972_),
    .Y(_04050_));
 sky130_fd_sc_hd__a22o_1 _11468_ (.A1(_03239_),
    .A2(_03229_),
    .B1(_03694_),
    .B2(_03695_),
    .X(_04051_));
 sky130_fd_sc_hd__nand3_1 _11469_ (.A(_04050_),
    .B(_03696_),
    .C(_04051_),
    .Y(_04052_));
 sky130_fd_sc_hd__a21o_1 _11470_ (.A1(_03696_),
    .A2(_04051_),
    .B1(_04050_),
    .X(_04053_));
 sky130_fd_sc_hd__nand3_1 _11471_ (.A(_04049_),
    .B(_04052_),
    .C(_04053_),
    .Y(_04054_));
 sky130_fd_sc_hd__a21o_1 _11472_ (.A1(_04052_),
    .A2(_04053_),
    .B1(_04049_),
    .X(_04055_));
 sky130_fd_sc_hd__nand4_4 _11473_ (.A(_04047_),
    .B(_04048_),
    .C(_04054_),
    .D(_04055_),
    .Y(_04056_));
 sky130_fd_sc_hd__a22o_1 _11474_ (.A1(_04047_),
    .A2(_04048_),
    .B1(_04054_),
    .B2(_04055_),
    .X(_04057_));
 sky130_fd_sc_hd__o211a_1 _11475_ (.A1(_03979_),
    .A2(_03992_),
    .B1(_04056_),
    .C1(_04057_),
    .X(_04058_));
 sky130_fd_sc_hd__a211oi_1 _11476_ (.A1(_04056_),
    .A2(_04057_),
    .B1(_03979_),
    .C1(_03992_),
    .Y(_04059_));
 sky130_fd_sc_hd__a21bo_1 _11477_ (.A1(_03981_),
    .A2(_03989_),
    .B1_N(_03988_),
    .X(_04060_));
 sky130_fd_sc_hd__nand3_1 _11478_ (.A(_03709_),
    .B(_03711_),
    .C(_03710_),
    .Y(_04061_));
 sky130_fd_sc_hd__a21o_1 _11479_ (.A1(_03711_),
    .A2(_03710_),
    .B1(_03709_),
    .X(_04062_));
 sky130_fd_sc_hd__o21bai_1 _11480_ (.A1(_03997_),
    .A2(_03999_),
    .B1_N(_03998_),
    .Y(_04063_));
 sky130_fd_sc_hd__nand3_2 _11481_ (.A(_04061_),
    .B(_04062_),
    .C(_04063_),
    .Y(_04064_));
 sky130_fd_sc_hd__a21o_1 _11482_ (.A1(_04061_),
    .A2(_04062_),
    .B1(_04063_),
    .X(_04065_));
 sky130_fd_sc_hd__nand2_1 _11483_ (.A(_03490_),
    .B(_02951_),
    .Y(_04066_));
 sky130_fd_sc_hd__a22oi_1 _11484_ (.A1(_03873_),
    .A2(_03038_),
    .B1(_03093_),
    .B2(_03872_),
    .Y(_04067_));
 sky130_fd_sc_hd__and4_1 _11485_ (.A(_03633_),
    .B(_02899_),
    .C(_03038_),
    .D(_03093_),
    .X(_04068_));
 sky130_fd_sc_hd__or2_1 _11486_ (.A(_04067_),
    .B(_04068_),
    .X(_04069_));
 sky130_fd_sc_hd__xor2_2 _11487_ (.A(_04066_),
    .B(_04069_),
    .X(_04070_));
 sky130_fd_sc_hd__nand3_2 _11488_ (.A(_04064_),
    .B(_04065_),
    .C(_04070_),
    .Y(_04071_));
 sky130_fd_sc_hd__a21o_1 _11489_ (.A1(_04064_),
    .A2(_04065_),
    .B1(_04070_),
    .X(_04072_));
 sky130_fd_sc_hd__and3_1 _11490_ (.A(_04060_),
    .B(_04071_),
    .C(_04072_),
    .X(_04073_));
 sky130_fd_sc_hd__a21oi_1 _11491_ (.A1(_04071_),
    .A2(_04072_),
    .B1(_04060_),
    .Y(_04074_));
 sky130_fd_sc_hd__a211oi_2 _11492_ (.A1(_04003_),
    .A2(_04010_),
    .B1(_04073_),
    .C1(_04074_),
    .Y(_04075_));
 sky130_fd_sc_hd__o211a_1 _11493_ (.A1(_04073_),
    .A2(_04074_),
    .B1(_04003_),
    .C1(_04010_),
    .X(_04076_));
 sky130_fd_sc_hd__or4_2 _11494_ (.A(_04058_),
    .B(_04059_),
    .C(_04075_),
    .D(_04076_),
    .X(_04077_));
 sky130_fd_sc_hd__o22ai_2 _11495_ (.A1(_04058_),
    .A2(_04059_),
    .B1(_04075_),
    .B2(_04076_),
    .Y(_04078_));
 sky130_fd_sc_hd__o211a_1 _11496_ (.A1(_03994_),
    .A2(_04018_),
    .B1(_04077_),
    .C1(_04078_),
    .X(_04079_));
 sky130_fd_sc_hd__a211oi_2 _11497_ (.A1(_04077_),
    .A2(_04078_),
    .B1(_03994_),
    .C1(_04018_),
    .Y(_04080_));
 sky130_fd_sc_hd__buf_8 _11498_ (.A(_03943_),
    .X(_04081_));
 sky130_fd_sc_hd__a31o_1 _11499_ (.A1(_04081_),
    .A2(_02953_),
    .A3(_04023_),
    .B1(_04026_),
    .X(_04082_));
 sky130_fd_sc_hd__and3_1 _11500_ (.A(_03996_),
    .B(_04010_),
    .C(_04011_),
    .X(_04083_));
 sky130_fd_sc_hd__a21oi_2 _11501_ (.A1(_04014_),
    .A2(_04013_),
    .B1(_04083_),
    .Y(_04084_));
 sky130_fd_sc_hd__nand2_1 _11502_ (.A(_03959_),
    .B(_03029_),
    .Y(_04085_));
 sky130_fd_sc_hd__nor2_1 _11503_ (.A(_04005_),
    .B(_04008_),
    .Y(_04086_));
 sky130_fd_sc_hd__o21a_1 _11504_ (.A1(_04007_),
    .A2(_04086_),
    .B1(_02890_),
    .X(_04087_));
 sky130_fd_sc_hd__or3_1 _11505_ (.A(_02890_),
    .B(_04007_),
    .C(_04086_),
    .X(_04088_));
 sky130_fd_sc_hd__and2b_1 _11506_ (.A_N(_04087_),
    .B(_04088_),
    .X(_04089_));
 sky130_fd_sc_hd__xnor2_2 _11507_ (.A(_04085_),
    .B(_04089_),
    .Y(_04090_));
 sky130_fd_sc_hd__xnor2_1 _11508_ (.A(_04084_),
    .B(_04090_),
    .Y(_04091_));
 sky130_fd_sc_hd__xnor2_1 _11509_ (.A(_04082_),
    .B(_04091_),
    .Y(_04092_));
 sky130_fd_sc_hd__o21ai_1 _11510_ (.A1(_04079_),
    .A2(_04080_),
    .B1(_04092_),
    .Y(_04093_));
 sky130_fd_sc_hd__or3_1 _11511_ (.A(_04079_),
    .B(_04080_),
    .C(_04092_),
    .X(_04094_));
 sky130_fd_sc_hd__o211a_1 _11512_ (.A1(_04019_),
    .A2(_04041_),
    .B1(_04093_),
    .C1(_04094_),
    .X(_04095_));
 sky130_fd_sc_hd__a211oi_2 _11513_ (.A1(_04094_),
    .A2(_04093_),
    .B1(_04041_),
    .C1(_04019_),
    .Y(_04096_));
 sky130_fd_sc_hd__a211oi_2 _11514_ (.A1(_04039_),
    .A2(_04040_),
    .B1(_04095_),
    .C1(_04096_),
    .Y(_04097_));
 sky130_fd_sc_hd__o211a_1 _11515_ (.A1(_04095_),
    .A2(_04096_),
    .B1(_04039_),
    .C1(_04040_),
    .X(_04098_));
 sky130_fd_sc_hd__a211oi_2 _11516_ (.A1(_04034_),
    .A2(_04038_),
    .B1(_04097_),
    .C1(_04098_),
    .Y(_04099_));
 sky130_fd_sc_hd__o211a_1 _11517_ (.A1(_04097_),
    .A2(_04098_),
    .B1(_04034_),
    .C1(_04038_),
    .X(_04100_));
 sky130_fd_sc_hd__nor2_2 _11518_ (.A(_04099_),
    .B(_04100_),
    .Y(_04101_));
 sky130_fd_sc_hd__clkbuf_4 _11519_ (.A(net2),
    .X(_04102_));
 sky130_fd_sc_hd__nand4_1 _11520_ (.A(_03678_),
    .B(_03018_),
    .C(_03233_),
    .D(_04102_),
    .Y(_04103_));
 sky130_fd_sc_hd__or3b_1 _11521_ (.A(_03766_),
    .B(_04103_),
    .C_N(_03779_),
    .X(_04104_));
 sky130_fd_sc_hd__nand4_1 _11522_ (.A(_04104_),
    .B(_03781_),
    .C(_03785_),
    .D(_03786_),
    .Y(_04105_));
 sky130_fd_sc_hd__a22o_1 _11523_ (.A1(_03757_),
    .A2(net16),
    .B1(net2),
    .B2(_03756_),
    .X(_04106_));
 sky130_fd_sc_hd__and4_1 _11524_ (.A(\wfg_stim_mem_top.cfg_gain_q[23] ),
    .B(\wfg_stim_mem_top.cfg_gain_q[10] ),
    .C(net15),
    .D(net32),
    .X(_04107_));
 sky130_fd_sc_hd__a21o_1 _11525_ (.A1(_04103_),
    .A2(_04106_),
    .B1(_04107_),
    .X(_04108_));
 sky130_fd_sc_hd__and2_1 _11526_ (.A(\wfg_stim_mem_top.cfg_gain_q[20] ),
    .B(_03770_),
    .X(_04109_));
 sky130_fd_sc_hd__nand4_1 _11527_ (.A(_02963_),
    .B(_02965_),
    .C(_03762_),
    .D(_03760_),
    .Y(_04110_));
 sky130_fd_sc_hd__a22o_1 _11528_ (.A1(_03773_),
    .A2(_03762_),
    .B1(_03760_),
    .B2(_03774_),
    .X(_04111_));
 sky130_fd_sc_hd__nand3_1 _11529_ (.A(_04109_),
    .B(_04110_),
    .C(_04111_),
    .Y(_04112_));
 sky130_fd_sc_hd__a21o_1 _11530_ (.A1(_04110_),
    .A2(_04111_),
    .B1(_04109_),
    .X(_04113_));
 sky130_fd_sc_hd__and3_1 _11531_ (.A(_04103_),
    .B(_04107_),
    .C(_04106_),
    .X(_04114_));
 sky130_fd_sc_hd__a31o_1 _11532_ (.A1(_04108_),
    .A2(_04112_),
    .A3(_04113_),
    .B1(_04114_),
    .X(_04115_));
 sky130_fd_sc_hd__a22o_1 _11533_ (.A1(_04104_),
    .A2(_03781_),
    .B1(_03785_),
    .B2(_03786_),
    .X(_04116_));
 sky130_fd_sc_hd__and3_2 _11534_ (.A(_04105_),
    .B(_04115_),
    .C(_04116_),
    .X(_04117_));
 sky130_fd_sc_hd__nand3_1 _11535_ (.A(_04105_),
    .B(_04115_),
    .C(_04116_),
    .Y(_04118_));
 sky130_fd_sc_hd__a21o_1 _11536_ (.A1(_04105_),
    .A2(_04116_),
    .B1(_04115_),
    .X(_04119_));
 sky130_fd_sc_hd__nand4_1 _11537_ (.A(_02943_),
    .B(_02940_),
    .C(_03680_),
    .D(_03769_),
    .Y(_04120_));
 sky130_fd_sc_hd__a22o_1 _11538_ (.A1(_02937_),
    .A2(_03680_),
    .B1(_03769_),
    .B2(_03143_),
    .X(_04121_));
 sky130_fd_sc_hd__nand4_1 _11539_ (.A(_03798_),
    .B(_03675_),
    .C(_04120_),
    .D(_04121_),
    .Y(_04122_));
 sky130_fd_sc_hd__nand2_1 _11540_ (.A(_04120_),
    .B(_04122_),
    .Y(_04123_));
 sky130_fd_sc_hd__a21bo_1 _11541_ (.A1(_04109_),
    .A2(_04111_),
    .B1_N(_04110_),
    .X(_04124_));
 sky130_fd_sc_hd__o21ai_1 _11542_ (.A1(_03792_),
    .A2(_03795_),
    .B1(_03794_),
    .Y(_04125_));
 sky130_fd_sc_hd__nand3_1 _11543_ (.A(_03796_),
    .B(_04124_),
    .C(_04125_),
    .Y(_04126_));
 sky130_fd_sc_hd__a21o_1 _11544_ (.A1(_03796_),
    .A2(_04125_),
    .B1(_04124_),
    .X(_04127_));
 sky130_fd_sc_hd__nand3_1 _11545_ (.A(_04123_),
    .B(_04126_),
    .C(_04127_),
    .Y(_04128_));
 sky130_fd_sc_hd__a21o_1 _11546_ (.A1(_04126_),
    .A2(_04127_),
    .B1(_04123_),
    .X(_04129_));
 sky130_fd_sc_hd__and4_2 _11547_ (.A(_04118_),
    .B(_04119_),
    .C(_04128_),
    .D(_04129_),
    .X(_04130_));
 sky130_fd_sc_hd__a22o_1 _11548_ (.A1(_03790_),
    .A2(_03791_),
    .B1(_03807_),
    .B2(_03808_),
    .X(_04131_));
 sky130_fd_sc_hd__o211ai_4 _11549_ (.A1(_04117_),
    .A2(_04130_),
    .B1(_04131_),
    .C1(_03809_),
    .Y(_04132_));
 sky130_fd_sc_hd__o211a_1 _11550_ (.A1(_04117_),
    .A2(_04130_),
    .B1(_04131_),
    .C1(_03809_),
    .X(_04133_));
 sky130_fd_sc_hd__a211oi_2 _11551_ (.A1(_03809_),
    .A2(_04131_),
    .B1(_04130_),
    .C1(_04117_),
    .Y(_04134_));
 sky130_fd_sc_hd__or3_1 _11552_ (.A(_03849_),
    .B(_03847_),
    .C(_03848_),
    .X(_04135_));
 sky130_fd_sc_hd__and2_1 _11553_ (.A(\wfg_stim_mem_top.cfg_gain_q[14] ),
    .B(_03286_),
    .X(_04136_));
 sky130_fd_sc_hd__a22o_1 _11554_ (.A1(_03209_),
    .A2(_03436_),
    .B1(_03793_),
    .B2(_02919_),
    .X(_04137_));
 sky130_fd_sc_hd__nand4_1 _11555_ (.A(_03217_),
    .B(_03212_),
    .C(_03436_),
    .D(_03793_),
    .Y(_04138_));
 sky130_fd_sc_hd__a21bo_1 _11556_ (.A1(_04136_),
    .A2(_04137_),
    .B1_N(_04138_),
    .X(_04139_));
 sky130_fd_sc_hd__o21ai_1 _11557_ (.A1(_03849_),
    .A2(_03848_),
    .B1(_03847_),
    .Y(_04140_));
 sky130_fd_sc_hd__nand3_1 _11558_ (.A(_04135_),
    .B(_04139_),
    .C(_04140_),
    .Y(_04141_));
 sky130_fd_sc_hd__a21o_1 _11559_ (.A1(_04135_),
    .A2(_04140_),
    .B1(_04139_),
    .X(_04142_));
 sky130_fd_sc_hd__nand2_1 _11560_ (.A(_02892_),
    .B(_03128_),
    .Y(_04143_));
 sky130_fd_sc_hd__a22oi_1 _11561_ (.A1(_02896_),
    .A2(_03228_),
    .B1(_03236_),
    .B2(_02894_),
    .Y(_04144_));
 sky130_fd_sc_hd__and4_1 _11562_ (.A(_03633_),
    .B(_02899_),
    .C(_03228_),
    .D(_03230_),
    .X(_04145_));
 sky130_fd_sc_hd__nor2_1 _11563_ (.A(_04144_),
    .B(_04145_),
    .Y(_04146_));
 sky130_fd_sc_hd__xnor2_2 _11564_ (.A(_04143_),
    .B(_04146_),
    .Y(_04147_));
 sky130_fd_sc_hd__nand3_1 _11565_ (.A(_04141_),
    .B(_04142_),
    .C(_04147_),
    .Y(_04148_));
 sky130_fd_sc_hd__and2_1 _11566_ (.A(_04141_),
    .B(_04148_),
    .X(_04149_));
 sky130_fd_sc_hd__a21bo_1 _11567_ (.A1(_04123_),
    .A2(_04127_),
    .B1_N(_04126_),
    .X(_04150_));
 sky130_fd_sc_hd__a21o_1 _11568_ (.A1(_03852_),
    .A2(_03853_),
    .B1(_03858_),
    .X(_04151_));
 sky130_fd_sc_hd__and3_1 _11569_ (.A(_03859_),
    .B(_04150_),
    .C(_04151_),
    .X(_04152_));
 sky130_fd_sc_hd__a21oi_1 _11570_ (.A1(_03859_),
    .A2(_04151_),
    .B1(_04150_),
    .Y(_04153_));
 sky130_fd_sc_hd__nor3_1 _11571_ (.A(_04149_),
    .B(_04152_),
    .C(_04153_),
    .Y(_04154_));
 sky130_fd_sc_hd__o21a_1 _11572_ (.A1(_04152_),
    .A2(_04153_),
    .B1(_04149_),
    .X(_04155_));
 sky130_fd_sc_hd__or4_4 _11573_ (.A(_04133_),
    .B(_04134_),
    .C(_04154_),
    .D(_04155_),
    .X(_04156_));
 sky130_fd_sc_hd__o22a_1 _11574_ (.A1(_03841_),
    .A2(_03842_),
    .B1(_03882_),
    .B2(_03883_),
    .X(_04157_));
 sky130_fd_sc_hd__a211oi_4 _11575_ (.A1(_04132_),
    .A2(_04156_),
    .B1(_04157_),
    .C1(_03884_),
    .Y(_04158_));
 sky130_fd_sc_hd__o211a_1 _11576_ (.A1(_03884_),
    .A2(_04157_),
    .B1(_04156_),
    .C1(_04132_),
    .X(_04159_));
 sky130_fd_sc_hd__a31o_1 _11577_ (.A1(_03869_),
    .A2(_03129_),
    .A3(_04146_),
    .B1(_04145_),
    .X(_04160_));
 sky130_fd_sc_hd__nand2_1 _11578_ (.A(_02887_),
    .B(_03040_),
    .Y(_04161_));
 sky130_fd_sc_hd__xnor2_1 _11579_ (.A(_04160_),
    .B(_04161_),
    .Y(_04162_));
 sky130_fd_sc_hd__and3_1 _11580_ (.A(_02907_),
    .B(_03274_),
    .C(_04162_),
    .X(_04163_));
 sky130_fd_sc_hd__a31o_1 _11581_ (.A1(_03944_),
    .A2(_03040_),
    .A3(_04160_),
    .B1(_04163_),
    .X(_04164_));
 sky130_fd_sc_hd__o21ba_1 _11582_ (.A1(_04149_),
    .A2(_04153_),
    .B1_N(_04152_),
    .X(_04165_));
 sky130_fd_sc_hd__a21oi_1 _11583_ (.A1(_02908_),
    .A2(_03129_),
    .B1(_03950_),
    .Y(_04166_));
 sky130_fd_sc_hd__nor2_1 _11584_ (.A(_03951_),
    .B(_04166_),
    .Y(_04167_));
 sky130_fd_sc_hd__xnor2_1 _11585_ (.A(_04165_),
    .B(_04167_),
    .Y(_04168_));
 sky130_fd_sc_hd__xnor2_1 _11586_ (.A(_04164_),
    .B(_04168_),
    .Y(_04169_));
 sky130_fd_sc_hd__nor3_2 _11587_ (.A(_04158_),
    .B(_04159_),
    .C(_04169_),
    .Y(_04170_));
 sky130_fd_sc_hd__o21ai_2 _11588_ (.A1(_03940_),
    .A2(_03941_),
    .B1(_03963_),
    .Y(_04171_));
 sky130_fd_sc_hd__or3_1 _11589_ (.A(_03940_),
    .B(_03941_),
    .C(_03963_),
    .X(_04172_));
 sky130_fd_sc_hd__o211ai_4 _11590_ (.A1(_04158_),
    .A2(_04170_),
    .B1(_04171_),
    .C1(_04172_),
    .Y(_04173_));
 sky130_fd_sc_hd__and2b_1 _11591_ (.A_N(_04165_),
    .B(_04167_),
    .X(_04174_));
 sky130_fd_sc_hd__and2_1 _11592_ (.A(_04164_),
    .B(_04168_),
    .X(_04175_));
 sky130_fd_sc_hd__a211o_1 _11593_ (.A1(_04172_),
    .A2(_04171_),
    .B1(_04170_),
    .C1(_04158_),
    .X(_04176_));
 sky130_fd_sc_hd__o211ai_4 _11594_ (.A1(_04174_),
    .A2(_04175_),
    .B1(_04173_),
    .C1(_04176_),
    .Y(_04177_));
 sky130_fd_sc_hd__a211oi_1 _11595_ (.A1(_04035_),
    .A2(_04036_),
    .B1(_04033_),
    .C1(_04037_),
    .Y(_04178_));
 sky130_fd_sc_hd__o211a_1 _11596_ (.A1(_04033_),
    .A2(_04037_),
    .B1(_04035_),
    .C1(_04036_),
    .X(_04179_));
 sky130_fd_sc_hd__a211oi_2 _11597_ (.A1(_04173_),
    .A2(_04177_),
    .B1(_04178_),
    .C1(_04179_),
    .Y(_04180_));
 sky130_fd_sc_hd__o211a_1 _11598_ (.A1(_04178_),
    .A2(_04179_),
    .B1(_04173_),
    .C1(_04177_),
    .X(_04181_));
 sky130_fd_sc_hd__nor2_2 _11599_ (.A(_04180_),
    .B(_04181_),
    .Y(_04182_));
 sky130_fd_sc_hd__nand2_1 _11600_ (.A(_04101_),
    .B(_04182_),
    .Y(_04183_));
 sky130_fd_sc_hd__a211o_1 _11601_ (.A1(_04173_),
    .A2(_04176_),
    .B1(_04174_),
    .C1(_04175_),
    .X(_04184_));
 sky130_fd_sc_hd__clkbuf_4 _11602_ (.A(net32),
    .X(_04185_));
 sky130_fd_sc_hd__nand4_1 _11603_ (.A(_03678_),
    .B(_03679_),
    .C(net15),
    .D(_04185_),
    .Y(_04186_));
 sky130_fd_sc_hd__or3b_1 _11604_ (.A(_03780_),
    .B(_04186_),
    .C_N(_04106_),
    .X(_04187_));
 sky130_fd_sc_hd__nand4_2 _11605_ (.A(_04187_),
    .B(_04108_),
    .C(_04112_),
    .D(_04113_),
    .Y(_04188_));
 sky130_fd_sc_hd__a22o_1 _11606_ (.A1(_03757_),
    .A2(net15),
    .B1(_04185_),
    .B2(_03756_),
    .X(_04189_));
 sky130_fd_sc_hd__and4_1 _11607_ (.A(_03013_),
    .B(_03757_),
    .C(net14),
    .D(net31),
    .X(_04190_));
 sky130_fd_sc_hd__a21o_1 _11608_ (.A1(_04186_),
    .A2(_04189_),
    .B1(_04190_),
    .X(_04191_));
 sky130_fd_sc_hd__nand2_1 _11609_ (.A(\wfg_stim_mem_top.cfg_gain_q[20] ),
    .B(_03762_),
    .Y(_04192_));
 sky130_fd_sc_hd__and4_1 _11610_ (.A(_02959_),
    .B(\wfg_stim_mem_top.cfg_gain_q[21] ),
    .C(net3),
    .D(net2),
    .X(_04193_));
 sky130_fd_sc_hd__a22oi_2 _11611_ (.A1(_02954_),
    .A2(net3),
    .B1(_04102_),
    .B2(_02959_),
    .Y(_04194_));
 sky130_fd_sc_hd__or3_1 _11612_ (.A(_04192_),
    .B(_04193_),
    .C(_04194_),
    .X(_04195_));
 sky130_fd_sc_hd__o21ai_1 _11613_ (.A1(_04193_),
    .A2(_04194_),
    .B1(_04192_),
    .Y(_04196_));
 sky130_fd_sc_hd__and3_1 _11614_ (.A(_04186_),
    .B(_04190_),
    .C(_04189_),
    .X(_04197_));
 sky130_fd_sc_hd__a31o_1 _11615_ (.A1(_04191_),
    .A2(_04195_),
    .A3(_04196_),
    .B1(_04197_),
    .X(_04198_));
 sky130_fd_sc_hd__a22o_1 _11616_ (.A1(_04187_),
    .A2(_04108_),
    .B1(_04112_),
    .B2(_04113_),
    .X(_04199_));
 sky130_fd_sc_hd__nand3_4 _11617_ (.A(_04188_),
    .B(_04198_),
    .C(_04199_),
    .Y(_04200_));
 sky130_fd_sc_hd__a21o_1 _11618_ (.A1(_04188_),
    .A2(_04199_),
    .B1(_04198_),
    .X(_04201_));
 sky130_fd_sc_hd__and4_1 _11619_ (.A(\wfg_stim_mem_top.cfg_gain_q[19] ),
    .B(\wfg_stim_mem_top.cfg_gain_q[18] ),
    .C(net6),
    .D(net5),
    .X(_04202_));
 sky130_fd_sc_hd__nand2_1 _11620_ (.A(\wfg_stim_mem_top.cfg_gain_q[17] ),
    .B(_03680_),
    .Y(_04203_));
 sky130_fd_sc_hd__a22oi_1 _11621_ (.A1(_02937_),
    .A2(_03769_),
    .B1(_03770_),
    .B2(_03143_),
    .Y(_04204_));
 sky130_fd_sc_hd__or3_1 _11622_ (.A(_04202_),
    .B(_04203_),
    .C(_04204_),
    .X(_04205_));
 sky130_fd_sc_hd__or2b_1 _11623_ (.A(_04202_),
    .B_N(_04205_),
    .X(_04206_));
 sky130_fd_sc_hd__o21bai_1 _11624_ (.A1(_04192_),
    .A2(_04194_),
    .B1_N(_04193_),
    .Y(_04207_));
 sky130_fd_sc_hd__a22o_1 _11625_ (.A1(_02934_),
    .A2(_03597_),
    .B1(_04120_),
    .B2(_04121_),
    .X(_04208_));
 sky130_fd_sc_hd__nand3_1 _11626_ (.A(_04122_),
    .B(_04207_),
    .C(_04208_),
    .Y(_04209_));
 sky130_fd_sc_hd__a21o_1 _11627_ (.A1(_04122_),
    .A2(_04208_),
    .B1(_04207_),
    .X(_04210_));
 sky130_fd_sc_hd__nand3_1 _11628_ (.A(_04206_),
    .B(_04209_),
    .C(_04210_),
    .Y(_04211_));
 sky130_fd_sc_hd__a21o_1 _11629_ (.A1(_04209_),
    .A2(_04210_),
    .B1(_04206_),
    .X(_04212_));
 sky130_fd_sc_hd__nand4_4 _11630_ (.A(_04200_),
    .B(_04201_),
    .C(_04211_),
    .D(_04212_),
    .Y(_04213_));
 sky130_fd_sc_hd__a22oi_4 _11631_ (.A1(_04118_),
    .A2(_04119_),
    .B1(_04128_),
    .B2(_04129_),
    .Y(_04214_));
 sky130_fd_sc_hd__a211oi_4 _11632_ (.A1(_04200_),
    .A2(_04213_),
    .B1(_04214_),
    .C1(_04130_),
    .Y(_04215_));
 sky130_fd_sc_hd__o211a_1 _11633_ (.A1(_04130_),
    .A2(_04214_),
    .B1(_04213_),
    .C1(_04200_),
    .X(_04216_));
 sky130_fd_sc_hd__nand3_1 _11634_ (.A(_04138_),
    .B(_04136_),
    .C(_04137_),
    .Y(_04217_));
 sky130_fd_sc_hd__nand2_1 _11635_ (.A(\wfg_stim_mem_top.cfg_gain_q[14] ),
    .B(_03436_),
    .Y(_04218_));
 sky130_fd_sc_hd__a22oi_2 _11636_ (.A1(_03209_),
    .A2(_03793_),
    .B1(_03674_),
    .B2(_03217_),
    .Y(_04219_));
 sky130_fd_sc_hd__and4_1 _11637_ (.A(_02919_),
    .B(\wfg_stim_mem_top.cfg_gain_q[15] ),
    .C(net9),
    .D(_03674_),
    .X(_04220_));
 sky130_fd_sc_hd__o21bai_1 _11638_ (.A1(_04218_),
    .A2(_04219_),
    .B1_N(_04220_),
    .Y(_04221_));
 sky130_fd_sc_hd__a22o_1 _11639_ (.A1(_03529_),
    .A2(_03287_),
    .B1(_04138_),
    .B2(_04137_),
    .X(_04222_));
 sky130_fd_sc_hd__nand3_1 _11640_ (.A(_04217_),
    .B(_04221_),
    .C(_04222_),
    .Y(_04223_));
 sky130_fd_sc_hd__a21o_1 _11641_ (.A1(_04217_),
    .A2(_04222_),
    .B1(_04221_),
    .X(_04224_));
 sky130_fd_sc_hd__nand2_1 _11642_ (.A(\wfg_stim_mem_top.cfg_gain_q[9] ),
    .B(_03248_),
    .Y(_04225_));
 sky130_fd_sc_hd__a22oi_1 _11643_ (.A1(_02899_),
    .A2(_03230_),
    .B1(_03279_),
    .B2(_03633_),
    .Y(_04226_));
 sky130_fd_sc_hd__and4_1 _11644_ (.A(\wfg_stim_mem_top.cfg_gain_q[13] ),
    .B(\wfg_stim_mem_top.cfg_gain_q[12] ),
    .C(_03230_),
    .D(_03279_),
    .X(_04227_));
 sky130_fd_sc_hd__nor2_1 _11645_ (.A(_04226_),
    .B(_04227_),
    .Y(_04228_));
 sky130_fd_sc_hd__xnor2_2 _11646_ (.A(_04225_),
    .B(_04228_),
    .Y(_04229_));
 sky130_fd_sc_hd__nand3_1 _11647_ (.A(_04223_),
    .B(_04224_),
    .C(_04229_),
    .Y(_04230_));
 sky130_fd_sc_hd__nand2_1 _11648_ (.A(_04223_),
    .B(_04230_),
    .Y(_04231_));
 sky130_fd_sc_hd__a21bo_1 _11649_ (.A1(_04206_),
    .A2(_04210_),
    .B1_N(_04209_),
    .X(_04232_));
 sky130_fd_sc_hd__a21o_1 _11650_ (.A1(_04141_),
    .A2(_04142_),
    .B1(_04147_),
    .X(_04233_));
 sky130_fd_sc_hd__nand3_1 _11651_ (.A(_04148_),
    .B(_04232_),
    .C(_04233_),
    .Y(_04234_));
 sky130_fd_sc_hd__a21o_1 _11652_ (.A1(_04148_),
    .A2(_04233_),
    .B1(_04232_),
    .X(_04235_));
 sky130_fd_sc_hd__and3_1 _11653_ (.A(_04231_),
    .B(_04234_),
    .C(_04235_),
    .X(_04236_));
 sky130_fd_sc_hd__a21oi_2 _11654_ (.A1(_04234_),
    .A2(_04235_),
    .B1(_04231_),
    .Y(_04237_));
 sky130_fd_sc_hd__nor4_4 _11655_ (.A(_04215_),
    .B(_04216_),
    .C(_04236_),
    .D(_04237_),
    .Y(_04238_));
 sky130_fd_sc_hd__o22ai_2 _11656_ (.A1(_04133_),
    .A2(_04134_),
    .B1(_04154_),
    .B2(_04155_),
    .Y(_04239_));
 sky130_fd_sc_hd__o211a_2 _11657_ (.A1(_04215_),
    .A2(_04238_),
    .B1(_04239_),
    .C1(_04156_),
    .X(_04240_));
 sky130_fd_sc_hd__a211oi_2 _11658_ (.A1(_04156_),
    .A2(_04239_),
    .B1(_04238_),
    .C1(_04215_),
    .Y(_04241_));
 sky130_fd_sc_hd__a31o_1 _11659_ (.A1(_03869_),
    .A2(_03274_),
    .A3(_04228_),
    .B1(_04227_),
    .X(_04242_));
 sky130_fd_sc_hd__nand2_1 _11660_ (.A(_02887_),
    .B(_03095_),
    .Y(_04243_));
 sky130_fd_sc_hd__xnor2_1 _11661_ (.A(_04242_),
    .B(_04243_),
    .Y(_04244_));
 sky130_fd_sc_hd__and3_1 _11662_ (.A(_02907_),
    .B(_03234_),
    .C(_04244_),
    .X(_04245_));
 sky130_fd_sc_hd__a31o_1 _11663_ (.A1(_03943_),
    .A2(_03095_),
    .A3(_04242_),
    .B1(_04245_),
    .X(_04246_));
 sky130_fd_sc_hd__a21boi_2 _11664_ (.A1(_04231_),
    .A2(_04235_),
    .B1_N(_04234_),
    .Y(_04247_));
 sky130_fd_sc_hd__a21oi_1 _11665_ (.A1(_03947_),
    .A2(_03274_),
    .B1(_04162_),
    .Y(_04248_));
 sky130_fd_sc_hd__nor2_1 _11666_ (.A(_04163_),
    .B(_04248_),
    .Y(_04249_));
 sky130_fd_sc_hd__xnor2_1 _11667_ (.A(_04247_),
    .B(_04249_),
    .Y(_04250_));
 sky130_fd_sc_hd__xnor2_1 _11668_ (.A(_04246_),
    .B(_04250_),
    .Y(_04251_));
 sky130_fd_sc_hd__nor3_1 _11669_ (.A(_04240_),
    .B(_04241_),
    .C(_04251_),
    .Y(_04252_));
 sky130_fd_sc_hd__o21ai_1 _11670_ (.A1(_04158_),
    .A2(_04159_),
    .B1(_04169_),
    .Y(_04253_));
 sky130_fd_sc_hd__or3_1 _11671_ (.A(_04158_),
    .B(_04159_),
    .C(_04169_),
    .X(_04254_));
 sky130_fd_sc_hd__o211ai_2 _11672_ (.A1(_04240_),
    .A2(_04252_),
    .B1(_04253_),
    .C1(_04254_),
    .Y(_04255_));
 sky130_fd_sc_hd__inv_2 _11673_ (.A(_04255_),
    .Y(_04256_));
 sky130_fd_sc_hd__and2b_1 _11674_ (.A_N(_04247_),
    .B(_04249_),
    .X(_04257_));
 sky130_fd_sc_hd__and2_1 _11675_ (.A(_04246_),
    .B(_04250_),
    .X(_04258_));
 sky130_fd_sc_hd__a211o_1 _11676_ (.A1(_04254_),
    .A2(_04253_),
    .B1(_04252_),
    .C1(_04240_),
    .X(_04259_));
 sky130_fd_sc_hd__o211a_1 _11677_ (.A1(_04257_),
    .A2(_04258_),
    .B1(_04255_),
    .C1(_04259_),
    .X(_04260_));
 sky130_fd_sc_hd__a211o_1 _11678_ (.A1(_04177_),
    .A2(_04184_),
    .B1(_04256_),
    .C1(_04260_),
    .X(_04261_));
 sky130_fd_sc_hd__o211a_1 _11679_ (.A1(_04256_),
    .A2(_04260_),
    .B1(_04177_),
    .C1(_04184_),
    .X(_04262_));
 sky130_fd_sc_hd__inv_2 _11680_ (.A(_04262_),
    .Y(_04263_));
 sky130_fd_sc_hd__nand2_2 _11681_ (.A(_04261_),
    .B(_04263_),
    .Y(_04264_));
 sky130_fd_sc_hd__a211oi_1 _11682_ (.A1(_04255_),
    .A2(_04259_),
    .B1(_04257_),
    .C1(_04258_),
    .Y(_04265_));
 sky130_fd_sc_hd__nor2_1 _11683_ (.A(_04260_),
    .B(_04265_),
    .Y(_04266_));
 sky130_fd_sc_hd__nand4_1 _11684_ (.A(_03013_),
    .B(_03018_),
    .C(net14),
    .D(net31),
    .Y(_04267_));
 sky130_fd_sc_hd__or3b_1 _11685_ (.A(_04107_),
    .B(_04267_),
    .C_N(_04189_),
    .X(_04268_));
 sky130_fd_sc_hd__nand4_1 _11686_ (.A(_04268_),
    .B(_04191_),
    .C(_04195_),
    .D(_04196_),
    .Y(_04269_));
 sky130_fd_sc_hd__clkbuf_4 _11687_ (.A(net31),
    .X(_04270_));
 sky130_fd_sc_hd__a22o_1 _11688_ (.A1(_03018_),
    .A2(_03230_),
    .B1(_04270_),
    .B2(_03013_),
    .X(_04271_));
 sky130_fd_sc_hd__and4_1 _11689_ (.A(_03756_),
    .B(_03757_),
    .C(net13),
    .D(net30),
    .X(_04272_));
 sky130_fd_sc_hd__a21o_1 _11690_ (.A1(_04267_),
    .A2(_04271_),
    .B1(_04272_),
    .X(_04273_));
 sky130_fd_sc_hd__and2_1 _11691_ (.A(\wfg_stim_mem_top.cfg_gain_q[20] ),
    .B(_03760_),
    .X(_04274_));
 sky130_fd_sc_hd__nand4_1 _11692_ (.A(_02963_),
    .B(_03773_),
    .C(_04102_),
    .D(_04185_),
    .Y(_04275_));
 sky130_fd_sc_hd__a22o_1 _11693_ (.A1(_02954_),
    .A2(_04102_),
    .B1(_04185_),
    .B2(_03774_),
    .X(_04276_));
 sky130_fd_sc_hd__nand3_1 _11694_ (.A(_04274_),
    .B(_04275_),
    .C(_04276_),
    .Y(_04277_));
 sky130_fd_sc_hd__a21o_1 _11695_ (.A1(_04275_),
    .A2(_04276_),
    .B1(_04274_),
    .X(_04278_));
 sky130_fd_sc_hd__and3_1 _11696_ (.A(_04267_),
    .B(_04272_),
    .C(_04271_),
    .X(_04279_));
 sky130_fd_sc_hd__a31o_1 _11697_ (.A1(_04273_),
    .A2(_04277_),
    .A3(_04278_),
    .B1(_04279_),
    .X(_04280_));
 sky130_fd_sc_hd__a22o_1 _11698_ (.A1(_04268_),
    .A2(_04191_),
    .B1(_04195_),
    .B2(_04196_),
    .X(_04281_));
 sky130_fd_sc_hd__and3_2 _11699_ (.A(_04269_),
    .B(_04280_),
    .C(_04281_),
    .X(_04282_));
 sky130_fd_sc_hd__nand3_1 _11700_ (.A(_04269_),
    .B(_04280_),
    .C(_04281_),
    .Y(_04283_));
 sky130_fd_sc_hd__a21o_1 _11701_ (.A1(_04269_),
    .A2(_04281_),
    .B1(_04280_),
    .X(_04284_));
 sky130_fd_sc_hd__nand4_1 _11702_ (.A(_03799_),
    .B(_03830_),
    .C(_03771_),
    .D(_03762_),
    .Y(_04285_));
 sky130_fd_sc_hd__clkbuf_4 _11703_ (.A(_03812_),
    .X(_04286_));
 sky130_fd_sc_hd__a22o_1 _11704_ (.A1(_02940_),
    .A2(_03770_),
    .B1(_03762_),
    .B2(_02943_),
    .X(_04287_));
 sky130_fd_sc_hd__nand4_1 _11705_ (.A(_03798_),
    .B(_04286_),
    .C(_04285_),
    .D(_04287_),
    .Y(_04288_));
 sky130_fd_sc_hd__nand2_1 _11706_ (.A(_04285_),
    .B(_04288_),
    .Y(_04289_));
 sky130_fd_sc_hd__a21bo_1 _11707_ (.A1(_04274_),
    .A2(_04276_),
    .B1_N(_04275_),
    .X(_04290_));
 sky130_fd_sc_hd__o21ai_1 _11708_ (.A1(_04202_),
    .A2(_04204_),
    .B1(_04203_),
    .Y(_04291_));
 sky130_fd_sc_hd__nand3_1 _11709_ (.A(_04205_),
    .B(_04290_),
    .C(_04291_),
    .Y(_04292_));
 sky130_fd_sc_hd__a21o_1 _11710_ (.A1(_04205_),
    .A2(_04291_),
    .B1(_04290_),
    .X(_04293_));
 sky130_fd_sc_hd__nand3_1 _11711_ (.A(_04289_),
    .B(_04292_),
    .C(_04293_),
    .Y(_04294_));
 sky130_fd_sc_hd__a21o_1 _11712_ (.A1(_04292_),
    .A2(_04293_),
    .B1(_04289_),
    .X(_04295_));
 sky130_fd_sc_hd__and4_2 _11713_ (.A(_04283_),
    .B(_04284_),
    .C(_04294_),
    .D(_04295_),
    .X(_04296_));
 sky130_fd_sc_hd__a22o_1 _11714_ (.A1(_04200_),
    .A2(_04201_),
    .B1(_04211_),
    .B2(_04212_),
    .X(_04297_));
 sky130_fd_sc_hd__o211ai_4 _11715_ (.A1(_04282_),
    .A2(_04296_),
    .B1(_04297_),
    .C1(_04213_),
    .Y(_04298_));
 sky130_fd_sc_hd__o211a_1 _11716_ (.A1(_04282_),
    .A2(_04296_),
    .B1(_04297_),
    .C1(_04213_),
    .X(_04299_));
 sky130_fd_sc_hd__a211oi_2 _11717_ (.A1(_04213_),
    .A2(_04297_),
    .B1(_04296_),
    .C1(_04282_),
    .Y(_04300_));
 sky130_fd_sc_hd__or3_1 _11718_ (.A(_04220_),
    .B(_04218_),
    .C(_04219_),
    .X(_04301_));
 sky130_fd_sc_hd__and2_1 _11719_ (.A(\wfg_stim_mem_top.cfg_gain_q[14] ),
    .B(_03793_),
    .X(_04302_));
 sky130_fd_sc_hd__a22o_1 _11720_ (.A1(_03209_),
    .A2(_03674_),
    .B1(_03680_),
    .B2(_02919_),
    .X(_04303_));
 sky130_fd_sc_hd__nand4_1 _11721_ (.A(_02920_),
    .B(_02922_),
    .C(_03597_),
    .D(_03894_),
    .Y(_04304_));
 sky130_fd_sc_hd__a21bo_1 _11722_ (.A1(_04302_),
    .A2(_04303_),
    .B1_N(_04304_),
    .X(_04305_));
 sky130_fd_sc_hd__o21ai_1 _11723_ (.A1(_04220_),
    .A2(_04219_),
    .B1(_04218_),
    .Y(_04306_));
 sky130_fd_sc_hd__nand3_1 _11724_ (.A(_04301_),
    .B(_04305_),
    .C(_04306_),
    .Y(_04307_));
 sky130_fd_sc_hd__a21o_1 _11725_ (.A1(_04301_),
    .A2(_04306_),
    .B1(_04305_),
    .X(_04308_));
 sky130_fd_sc_hd__nand2_1 _11726_ (.A(_02892_),
    .B(_03271_),
    .Y(_04309_));
 sky130_fd_sc_hd__a22oi_1 _11727_ (.A1(_02896_),
    .A2(_03280_),
    .B1(_03287_),
    .B2(_03636_),
    .Y(_04310_));
 sky130_fd_sc_hd__and4_1 _11728_ (.A(_03633_),
    .B(_02899_),
    .C(_03279_),
    .D(_03286_),
    .X(_04311_));
 sky130_fd_sc_hd__nor2_1 _11729_ (.A(_04310_),
    .B(_04311_),
    .Y(_04312_));
 sky130_fd_sc_hd__xnor2_1 _11730_ (.A(_04309_),
    .B(_04312_),
    .Y(_04313_));
 sky130_fd_sc_hd__nand3_1 _11731_ (.A(_04307_),
    .B(_04308_),
    .C(_04313_),
    .Y(_04314_));
 sky130_fd_sc_hd__and2_1 _11732_ (.A(_04307_),
    .B(_04314_),
    .X(_04315_));
 sky130_fd_sc_hd__a21bo_1 _11733_ (.A1(_04289_),
    .A2(_04293_),
    .B1_N(_04292_),
    .X(_04316_));
 sky130_fd_sc_hd__a21o_1 _11734_ (.A1(_04223_),
    .A2(_04224_),
    .B1(_04229_),
    .X(_04317_));
 sky130_fd_sc_hd__and3_1 _11735_ (.A(_04230_),
    .B(_04316_),
    .C(_04317_),
    .X(_04318_));
 sky130_fd_sc_hd__a21oi_1 _11736_ (.A1(_04230_),
    .A2(_04317_),
    .B1(_04316_),
    .Y(_04319_));
 sky130_fd_sc_hd__nor3_1 _11737_ (.A(_04315_),
    .B(_04318_),
    .C(_04319_),
    .Y(_04320_));
 sky130_fd_sc_hd__o21a_1 _11738_ (.A1(_04318_),
    .A2(_04319_),
    .B1(_04315_),
    .X(_04321_));
 sky130_fd_sc_hd__or4_4 _11739_ (.A(_04299_),
    .B(_04300_),
    .C(_04320_),
    .D(_04321_),
    .X(_04322_));
 sky130_fd_sc_hd__o22a_1 _11740_ (.A1(_04215_),
    .A2(_04216_),
    .B1(_04236_),
    .B2(_04237_),
    .X(_04323_));
 sky130_fd_sc_hd__a211oi_4 _11741_ (.A1(_04298_),
    .A2(_04322_),
    .B1(_04323_),
    .C1(_04238_),
    .Y(_04324_));
 sky130_fd_sc_hd__o211a_1 _11742_ (.A1(_04238_),
    .A2(_04323_),
    .B1(_04322_),
    .C1(_04298_),
    .X(_04325_));
 sky130_fd_sc_hd__a31o_1 _11743_ (.A1(_03869_),
    .A2(_03234_),
    .A3(_04312_),
    .B1(_04311_),
    .X(_04326_));
 sky130_fd_sc_hd__nand2_1 _11744_ (.A(_02886_),
    .B(_03129_),
    .Y(_04327_));
 sky130_fd_sc_hd__xnor2_1 _11745_ (.A(_04326_),
    .B(_04327_),
    .Y(_04328_));
 sky130_fd_sc_hd__and3_1 _11746_ (.A(_02907_),
    .B(_03314_),
    .C(_04328_),
    .X(_04329_));
 sky130_fd_sc_hd__a31o_1 _11747_ (.A1(_03943_),
    .A2(_03129_),
    .A3(_04326_),
    .B1(_04329_),
    .X(_04330_));
 sky130_fd_sc_hd__o21ba_1 _11748_ (.A1(_04315_),
    .A2(_04319_),
    .B1_N(_04318_),
    .X(_04331_));
 sky130_fd_sc_hd__a21oi_1 _11749_ (.A1(_02907_),
    .A2(_03234_),
    .B1(_04244_),
    .Y(_04332_));
 sky130_fd_sc_hd__nor2_1 _11750_ (.A(_04245_),
    .B(_04332_),
    .Y(_04333_));
 sky130_fd_sc_hd__xnor2_1 _11751_ (.A(_04331_),
    .B(_04333_),
    .Y(_04334_));
 sky130_fd_sc_hd__xnor2_1 _11752_ (.A(_04330_),
    .B(_04334_),
    .Y(_04335_));
 sky130_fd_sc_hd__nor3_1 _11753_ (.A(_04324_),
    .B(_04325_),
    .C(_04335_),
    .Y(_04336_));
 sky130_fd_sc_hd__o21ai_1 _11754_ (.A1(_04240_),
    .A2(_04241_),
    .B1(_04251_),
    .Y(_04337_));
 sky130_fd_sc_hd__or3_1 _11755_ (.A(_04240_),
    .B(_04241_),
    .C(_04251_),
    .X(_04338_));
 sky130_fd_sc_hd__o211a_1 _11756_ (.A1(_04324_),
    .A2(_04336_),
    .B1(_04337_),
    .C1(_04338_),
    .X(_04339_));
 sky130_fd_sc_hd__or3_1 _11757_ (.A(_04245_),
    .B(_04331_),
    .C(_04332_),
    .X(_04340_));
 sky130_fd_sc_hd__nand2_1 _11758_ (.A(_04330_),
    .B(_04334_),
    .Y(_04341_));
 sky130_fd_sc_hd__a211oi_1 _11759_ (.A1(_04338_),
    .A2(_04337_),
    .B1(_04336_),
    .C1(_04324_),
    .Y(_04342_));
 sky130_fd_sc_hd__a211oi_2 _11760_ (.A1(_04340_),
    .A2(_04341_),
    .B1(_04339_),
    .C1(_04342_),
    .Y(_04343_));
 sky130_fd_sc_hd__nor2_1 _11761_ (.A(_04339_),
    .B(_04343_),
    .Y(_04344_));
 sky130_fd_sc_hd__xor2_2 _11762_ (.A(_04266_),
    .B(_04344_),
    .X(_04345_));
 sky130_fd_sc_hd__clkbuf_4 _11763_ (.A(net30),
    .X(_04346_));
 sky130_fd_sc_hd__nand4_1 _11764_ (.A(_03759_),
    .B(_03679_),
    .C(_03279_),
    .D(_04346_),
    .Y(_04347_));
 sky130_fd_sc_hd__or3b_1 _11765_ (.A(_04190_),
    .B(_04347_),
    .C_N(_04271_),
    .X(_04348_));
 sky130_fd_sc_hd__nand4_2 _11766_ (.A(_04348_),
    .B(_04273_),
    .C(_04277_),
    .D(_04278_),
    .Y(_04349_));
 sky130_fd_sc_hd__a22o_1 _11767_ (.A1(_03757_),
    .A2(net13),
    .B1(net30),
    .B2(_03756_),
    .X(_04350_));
 sky130_fd_sc_hd__and4_1 _11768_ (.A(_03013_),
    .B(_03018_),
    .C(net11),
    .D(net29),
    .X(_04351_));
 sky130_fd_sc_hd__a21o_1 _11769_ (.A1(_04347_),
    .A2(_04350_),
    .B1(_04351_),
    .X(_04352_));
 sky130_fd_sc_hd__nand2_1 _11770_ (.A(\wfg_stim_mem_top.cfg_gain_q[20] ),
    .B(_04102_),
    .Y(_04353_));
 sky130_fd_sc_hd__a22oi_2 _11771_ (.A1(_02954_),
    .A2(_04185_),
    .B1(_04270_),
    .B2(_02959_),
    .Y(_04354_));
 sky130_fd_sc_hd__and4_1 _11772_ (.A(_02959_),
    .B(_02954_),
    .C(net32),
    .D(net31),
    .X(_04355_));
 sky130_fd_sc_hd__or3_1 _11773_ (.A(_04353_),
    .B(_04354_),
    .C(_04355_),
    .X(_04356_));
 sky130_fd_sc_hd__o21ai_1 _11774_ (.A1(_04354_),
    .A2(_04355_),
    .B1(_04353_),
    .Y(_04357_));
 sky130_fd_sc_hd__and3_1 _11775_ (.A(_04347_),
    .B(_04351_),
    .C(_04350_),
    .X(_04358_));
 sky130_fd_sc_hd__a31o_1 _11776_ (.A1(_04352_),
    .A2(_04356_),
    .A3(_04357_),
    .B1(_04358_),
    .X(_04359_));
 sky130_fd_sc_hd__a22o_1 _11777_ (.A1(_04348_),
    .A2(_04273_),
    .B1(_04277_),
    .B2(_04278_),
    .X(_04360_));
 sky130_fd_sc_hd__nand3_4 _11778_ (.A(_04349_),
    .B(_04359_),
    .C(_04360_),
    .Y(_04361_));
 sky130_fd_sc_hd__a21o_1 _11779_ (.A1(_04349_),
    .A2(_04360_),
    .B1(_04359_),
    .X(_04362_));
 sky130_fd_sc_hd__and4_1 _11780_ (.A(_03143_),
    .B(_02937_),
    .C(net4),
    .D(net3),
    .X(_04363_));
 sky130_fd_sc_hd__nand2_1 _11781_ (.A(_02934_),
    .B(_03770_),
    .Y(_04364_));
 sky130_fd_sc_hd__a22oi_1 _11782_ (.A1(_02940_),
    .A2(_03762_),
    .B1(_03760_),
    .B2(_02943_),
    .Y(_04365_));
 sky130_fd_sc_hd__or3_1 _11783_ (.A(_04363_),
    .B(_04364_),
    .C(_04365_),
    .X(_04366_));
 sky130_fd_sc_hd__or2b_1 _11784_ (.A(_04363_),
    .B_N(_04366_),
    .X(_04367_));
 sky130_fd_sc_hd__o21bai_2 _11785_ (.A1(_04353_),
    .A2(_04354_),
    .B1_N(_04355_),
    .Y(_04368_));
 sky130_fd_sc_hd__a22o_1 _11786_ (.A1(_02934_),
    .A2(_03812_),
    .B1(_04285_),
    .B2(_04287_),
    .X(_04369_));
 sky130_fd_sc_hd__nand3_1 _11787_ (.A(_04288_),
    .B(_04368_),
    .C(_04369_),
    .Y(_04370_));
 sky130_fd_sc_hd__a21o_1 _11788_ (.A1(_04288_),
    .A2(_04369_),
    .B1(_04368_),
    .X(_04371_));
 sky130_fd_sc_hd__nand3_1 _11789_ (.A(_04367_),
    .B(_04370_),
    .C(_04371_),
    .Y(_04372_));
 sky130_fd_sc_hd__a21o_1 _11790_ (.A1(_04370_),
    .A2(_04371_),
    .B1(_04367_),
    .X(_04373_));
 sky130_fd_sc_hd__nand4_4 _11791_ (.A(_04361_),
    .B(_04362_),
    .C(_04372_),
    .D(_04373_),
    .Y(_04374_));
 sky130_fd_sc_hd__a22oi_4 _11792_ (.A1(_04283_),
    .A2(_04284_),
    .B1(_04294_),
    .B2(_04295_),
    .Y(_04375_));
 sky130_fd_sc_hd__a211oi_4 _11793_ (.A1(_04361_),
    .A2(_04374_),
    .B1(_04375_),
    .C1(_04296_),
    .Y(_04376_));
 sky130_fd_sc_hd__o211a_1 _11794_ (.A1(_04296_),
    .A2(_04375_),
    .B1(_04374_),
    .C1(_04361_),
    .X(_04377_));
 sky130_fd_sc_hd__nand3_1 _11795_ (.A(_04304_),
    .B(_04302_),
    .C(_04303_),
    .Y(_04378_));
 sky130_fd_sc_hd__nand2_1 _11796_ (.A(_03529_),
    .B(_03597_),
    .Y(_04379_));
 sky130_fd_sc_hd__a22oi_2 _11797_ (.A1(_02922_),
    .A2(_03894_),
    .B1(_03812_),
    .B2(_02920_),
    .Y(_04380_));
 sky130_fd_sc_hd__and4_1 _11798_ (.A(_03217_),
    .B(_03209_),
    .C(_03680_),
    .D(_03769_),
    .X(_04381_));
 sky130_fd_sc_hd__o21bai_1 _11799_ (.A1(_04379_),
    .A2(_04380_),
    .B1_N(_04381_),
    .Y(_04382_));
 sky130_fd_sc_hd__a22o_1 _11800_ (.A1(_02926_),
    .A2(_03551_),
    .B1(_04304_),
    .B2(_04303_),
    .X(_04383_));
 sky130_fd_sc_hd__nand3_1 _11801_ (.A(_04378_),
    .B(_04382_),
    .C(_04383_),
    .Y(_04384_));
 sky130_fd_sc_hd__a21o_1 _11802_ (.A1(_04378_),
    .A2(_04383_),
    .B1(_04382_),
    .X(_04385_));
 sky130_fd_sc_hd__nand2_1 _11803_ (.A(_02892_),
    .B(_03229_),
    .Y(_04386_));
 sky130_fd_sc_hd__a22oi_1 _11804_ (.A1(_03637_),
    .A2(_03287_),
    .B1(_03684_),
    .B2(_03636_),
    .Y(_04387_));
 sky130_fd_sc_hd__and4_1 _11805_ (.A(\wfg_stim_mem_top.cfg_gain_q[13] ),
    .B(\wfg_stim_mem_top.cfg_gain_q[12] ),
    .C(_03286_),
    .D(_03436_),
    .X(_04388_));
 sky130_fd_sc_hd__nor2_1 _11806_ (.A(_04387_),
    .B(_04388_),
    .Y(_04389_));
 sky130_fd_sc_hd__xnor2_1 _11807_ (.A(_04386_),
    .B(_04389_),
    .Y(_04390_));
 sky130_fd_sc_hd__nand3_1 _11808_ (.A(_04384_),
    .B(_04385_),
    .C(_04390_),
    .Y(_04391_));
 sky130_fd_sc_hd__nand2_1 _11809_ (.A(_04384_),
    .B(_04391_),
    .Y(_04392_));
 sky130_fd_sc_hd__a21bo_1 _11810_ (.A1(_04367_),
    .A2(_04371_),
    .B1_N(_04370_),
    .X(_04393_));
 sky130_fd_sc_hd__a21o_1 _11811_ (.A1(_04307_),
    .A2(_04308_),
    .B1(_04313_),
    .X(_04394_));
 sky130_fd_sc_hd__nand3_1 _11812_ (.A(_04314_),
    .B(_04393_),
    .C(_04394_),
    .Y(_04395_));
 sky130_fd_sc_hd__a21o_1 _11813_ (.A1(_04314_),
    .A2(_04394_),
    .B1(_04393_),
    .X(_04396_));
 sky130_fd_sc_hd__and3_1 _11814_ (.A(_04392_),
    .B(_04395_),
    .C(_04396_),
    .X(_04397_));
 sky130_fd_sc_hd__a21oi_2 _11815_ (.A1(_04395_),
    .A2(_04396_),
    .B1(_04392_),
    .Y(_04398_));
 sky130_fd_sc_hd__nor4_4 _11816_ (.A(_04376_),
    .B(_04377_),
    .C(_04397_),
    .D(_04398_),
    .Y(_04399_));
 sky130_fd_sc_hd__o22ai_2 _11817_ (.A1(_04299_),
    .A2(_04300_),
    .B1(_04320_),
    .B2(_04321_),
    .Y(_04400_));
 sky130_fd_sc_hd__o211a_1 _11818_ (.A1(_04376_),
    .A2(_04399_),
    .B1(_04400_),
    .C1(_04322_),
    .X(_04401_));
 sky130_fd_sc_hd__a211oi_2 _11819_ (.A1(_04322_),
    .A2(_04400_),
    .B1(_04399_),
    .C1(_04376_),
    .Y(_04402_));
 sky130_fd_sc_hd__a31o_1 _11820_ (.A1(_03491_),
    .A2(_03314_),
    .A3(_04389_),
    .B1(_04388_),
    .X(_04403_));
 sky130_fd_sc_hd__nand2_1 _11821_ (.A(_02887_),
    .B(_03274_),
    .Y(_04404_));
 sky130_fd_sc_hd__xnor2_1 _11822_ (.A(_04403_),
    .B(_04404_),
    .Y(_04405_));
 sky130_fd_sc_hd__and3_1 _11823_ (.A(_02907_),
    .B(_03231_),
    .C(_04405_),
    .X(_04406_));
 sky130_fd_sc_hd__a31o_1 _11824_ (.A1(_03943_),
    .A2(_03274_),
    .A3(_04403_),
    .B1(_04406_),
    .X(_04407_));
 sky130_fd_sc_hd__a21boi_2 _11825_ (.A1(_04392_),
    .A2(_04396_),
    .B1_N(_04395_),
    .Y(_04408_));
 sky130_fd_sc_hd__a21oi_1 _11826_ (.A1(_02907_),
    .A2(_03314_),
    .B1(_04328_),
    .Y(_04409_));
 sky130_fd_sc_hd__nor2_1 _11827_ (.A(_04329_),
    .B(_04409_),
    .Y(_04410_));
 sky130_fd_sc_hd__xnor2_1 _11828_ (.A(_04408_),
    .B(_04410_),
    .Y(_04411_));
 sky130_fd_sc_hd__xnor2_1 _11829_ (.A(_04407_),
    .B(_04411_),
    .Y(_04412_));
 sky130_fd_sc_hd__nor3_1 _11830_ (.A(_04401_),
    .B(_04402_),
    .C(_04412_),
    .Y(_04413_));
 sky130_fd_sc_hd__o21ai_1 _11831_ (.A1(_04324_),
    .A2(_04325_),
    .B1(_04335_),
    .Y(_04414_));
 sky130_fd_sc_hd__or3_1 _11832_ (.A(_04324_),
    .B(_04325_),
    .C(_04335_),
    .X(_04415_));
 sky130_fd_sc_hd__o211ai_1 _11833_ (.A1(_04401_),
    .A2(_04413_),
    .B1(_04414_),
    .C1(_04415_),
    .Y(_04416_));
 sky130_fd_sc_hd__or3_1 _11834_ (.A(_04329_),
    .B(_04408_),
    .C(_04409_),
    .X(_04417_));
 sky130_fd_sc_hd__nand2_1 _11835_ (.A(_04407_),
    .B(_04411_),
    .Y(_04418_));
 sky130_fd_sc_hd__o211a_1 _11836_ (.A1(_04401_),
    .A2(_04413_),
    .B1(_04414_),
    .C1(_04415_),
    .X(_04419_));
 sky130_fd_sc_hd__a211oi_1 _11837_ (.A1(_04415_),
    .A2(_04414_),
    .B1(_04413_),
    .C1(_04401_),
    .Y(_04420_));
 sky130_fd_sc_hd__a211o_1 _11838_ (.A1(_04417_),
    .A2(_04418_),
    .B1(_04419_),
    .C1(_04420_),
    .X(_04421_));
 sky130_fd_sc_hd__o211a_1 _11839_ (.A1(_04339_),
    .A2(_04342_),
    .B1(_04340_),
    .C1(_04341_),
    .X(_04422_));
 sky130_fd_sc_hd__a211oi_1 _11840_ (.A1(_04416_),
    .A2(_04421_),
    .B1(_04343_),
    .C1(_04422_),
    .Y(_04423_));
 sky130_fd_sc_hd__o211ai_1 _11841_ (.A1(_04343_),
    .A2(_04422_),
    .B1(_04416_),
    .C1(_04421_),
    .Y(_04424_));
 sky130_fd_sc_hd__or2b_2 _11842_ (.A(_04423_),
    .B_N(_04424_),
    .X(_04425_));
 sky130_fd_sc_hd__clkbuf_4 _11843_ (.A(net29),
    .X(_04426_));
 sky130_fd_sc_hd__nand4_1 _11844_ (.A(_03678_),
    .B(_03679_),
    .C(net11),
    .D(_04426_),
    .Y(_04427_));
 sky130_fd_sc_hd__or3b_1 _11845_ (.A(_04272_),
    .B(_04427_),
    .C_N(_04350_),
    .X(_04428_));
 sky130_fd_sc_hd__nand4_2 _11846_ (.A(_04428_),
    .B(_04352_),
    .C(_04356_),
    .D(_04357_),
    .Y(_04429_));
 sky130_fd_sc_hd__a22o_1 _11847_ (.A1(_03679_),
    .A2(_03286_),
    .B1(_04426_),
    .B2(_03678_),
    .X(_04430_));
 sky130_fd_sc_hd__and4_1 _11848_ (.A(_03013_),
    .B(_03018_),
    .C(net10),
    .D(net28),
    .X(_04431_));
 sky130_fd_sc_hd__a21o_1 _11849_ (.A1(_04427_),
    .A2(_04430_),
    .B1(_04431_),
    .X(_04432_));
 sky130_fd_sc_hd__and2_1 _11850_ (.A(_02948_),
    .B(_04185_),
    .X(_04433_));
 sky130_fd_sc_hd__a22o_1 _11851_ (.A1(_03773_),
    .A2(_04270_),
    .B1(_04346_),
    .B2(_03774_),
    .X(_04434_));
 sky130_fd_sc_hd__nand4_1 _11852_ (.A(_02963_),
    .B(_02965_),
    .C(_04270_),
    .D(_04346_),
    .Y(_04435_));
 sky130_fd_sc_hd__nand3_1 _11853_ (.A(_04433_),
    .B(_04434_),
    .C(_04435_),
    .Y(_04436_));
 sky130_fd_sc_hd__a21o_1 _11854_ (.A1(_04434_),
    .A2(_04435_),
    .B1(_04433_),
    .X(_04437_));
 sky130_fd_sc_hd__and3_1 _11855_ (.A(_04427_),
    .B(_04431_),
    .C(_04430_),
    .X(_04438_));
 sky130_fd_sc_hd__a31o_1 _11856_ (.A1(_04432_),
    .A2(_04436_),
    .A3(_04437_),
    .B1(_04438_),
    .X(_04439_));
 sky130_fd_sc_hd__a22o_1 _11857_ (.A1(_04428_),
    .A2(_04352_),
    .B1(_04356_),
    .B2(_04357_),
    .X(_04440_));
 sky130_fd_sc_hd__and3_2 _11858_ (.A(_04429_),
    .B(_04439_),
    .C(_04440_),
    .X(_04441_));
 sky130_fd_sc_hd__nand3_1 _11859_ (.A(_04429_),
    .B(_04439_),
    .C(_04440_),
    .Y(_04442_));
 sky130_fd_sc_hd__a21o_1 _11860_ (.A1(_04429_),
    .A2(_04440_),
    .B1(_04439_),
    .X(_04443_));
 sky130_fd_sc_hd__buf_2 _11861_ (.A(_03760_),
    .X(_04444_));
 sky130_fd_sc_hd__clkbuf_4 _11862_ (.A(_04102_),
    .X(_04445_));
 sky130_fd_sc_hd__nand4_1 _11863_ (.A(_03144_),
    .B(_02938_),
    .C(_04444_),
    .D(_04445_),
    .Y(_04446_));
 sky130_fd_sc_hd__clkbuf_4 _11864_ (.A(_03762_),
    .X(_04447_));
 sky130_fd_sc_hd__buf_4 _11865_ (.A(_04447_),
    .X(_04448_));
 sky130_fd_sc_hd__a22o_1 _11866_ (.A1(_03830_),
    .A2(_03760_),
    .B1(_04102_),
    .B2(_03799_),
    .X(_04449_));
 sky130_fd_sc_hd__nand4_1 _11867_ (.A(_03798_),
    .B(_04448_),
    .C(_04446_),
    .D(_04449_),
    .Y(_04450_));
 sky130_fd_sc_hd__nand2_1 _11868_ (.A(_04446_),
    .B(_04450_),
    .Y(_04451_));
 sky130_fd_sc_hd__a21bo_1 _11869_ (.A1(_04433_),
    .A2(_04434_),
    .B1_N(_04435_),
    .X(_04452_));
 sky130_fd_sc_hd__o21ai_1 _11870_ (.A1(_04363_),
    .A2(_04365_),
    .B1(_04364_),
    .Y(_04453_));
 sky130_fd_sc_hd__nand3_1 _11871_ (.A(_04366_),
    .B(_04452_),
    .C(_04453_),
    .Y(_04454_));
 sky130_fd_sc_hd__a21o_1 _11872_ (.A1(_04366_),
    .A2(_04453_),
    .B1(_04452_),
    .X(_04455_));
 sky130_fd_sc_hd__nand3_1 _11873_ (.A(_04451_),
    .B(_04454_),
    .C(_04455_),
    .Y(_04456_));
 sky130_fd_sc_hd__a21o_1 _11874_ (.A1(_04454_),
    .A2(_04455_),
    .B1(_04451_),
    .X(_04457_));
 sky130_fd_sc_hd__and4_2 _11875_ (.A(_04442_),
    .B(_04443_),
    .C(_04456_),
    .D(_04457_),
    .X(_04458_));
 sky130_fd_sc_hd__a22o_1 _11876_ (.A1(_04361_),
    .A2(_04362_),
    .B1(_04372_),
    .B2(_04373_),
    .X(_04459_));
 sky130_fd_sc_hd__o211ai_4 _11877_ (.A1(_04441_),
    .A2(_04458_),
    .B1(_04459_),
    .C1(_04374_),
    .Y(_04460_));
 sky130_fd_sc_hd__o211a_1 _11878_ (.A1(_04441_),
    .A2(_04458_),
    .B1(_04459_),
    .C1(_04374_),
    .X(_04461_));
 sky130_fd_sc_hd__a211oi_2 _11879_ (.A1(_04374_),
    .A2(_04459_),
    .B1(_04458_),
    .C1(_04441_),
    .Y(_04462_));
 sky130_fd_sc_hd__or3_1 _11880_ (.A(_04381_),
    .B(_04379_),
    .C(_04380_),
    .X(_04463_));
 sky130_fd_sc_hd__and2_1 _11881_ (.A(_03529_),
    .B(_03894_),
    .X(_04464_));
 sky130_fd_sc_hd__a22o_1 _11882_ (.A1(_03531_),
    .A2(_03812_),
    .B1(_03771_),
    .B2(_03532_),
    .X(_04465_));
 sky130_fd_sc_hd__nand4_1 _11883_ (.A(_03218_),
    .B(_03210_),
    .C(_03812_),
    .D(_03771_),
    .Y(_04466_));
 sky130_fd_sc_hd__a21bo_1 _11884_ (.A1(_04464_),
    .A2(_04465_),
    .B1_N(_04466_),
    .X(_04467_));
 sky130_fd_sc_hd__o21ai_1 _11885_ (.A1(_04381_),
    .A2(_04380_),
    .B1(_04379_),
    .Y(_04468_));
 sky130_fd_sc_hd__nand3_1 _11886_ (.A(_04463_),
    .B(_04467_),
    .C(_04468_),
    .Y(_04469_));
 sky130_fd_sc_hd__a21o_1 _11887_ (.A1(_04463_),
    .A2(_04468_),
    .B1(_04467_),
    .X(_04470_));
 sky130_fd_sc_hd__nand2_1 _11888_ (.A(_03490_),
    .B(_03231_),
    .Y(_04471_));
 sky130_fd_sc_hd__a22oi_1 _11889_ (.A1(_03873_),
    .A2(_03684_),
    .B1(_03685_),
    .B2(_03872_),
    .Y(_04472_));
 sky130_fd_sc_hd__and4_1 _11890_ (.A(_03636_),
    .B(_03637_),
    .C(_03684_),
    .D(_03551_),
    .X(_04473_));
 sky130_fd_sc_hd__nor2_1 _11891_ (.A(_04472_),
    .B(_04473_),
    .Y(_04474_));
 sky130_fd_sc_hd__xnor2_1 _11892_ (.A(_04471_),
    .B(_04474_),
    .Y(_04475_));
 sky130_fd_sc_hd__nand3_1 _11893_ (.A(_04469_),
    .B(_04470_),
    .C(_04475_),
    .Y(_04476_));
 sky130_fd_sc_hd__and2_1 _11894_ (.A(_04469_),
    .B(_04476_),
    .X(_04477_));
 sky130_fd_sc_hd__a21bo_1 _11895_ (.A1(_04451_),
    .A2(_04455_),
    .B1_N(_04454_),
    .X(_04478_));
 sky130_fd_sc_hd__a21o_1 _11896_ (.A1(_04384_),
    .A2(_04385_),
    .B1(_04390_),
    .X(_04479_));
 sky130_fd_sc_hd__and3_1 _11897_ (.A(_04391_),
    .B(_04478_),
    .C(_04479_),
    .X(_04480_));
 sky130_fd_sc_hd__a21oi_1 _11898_ (.A1(_04391_),
    .A2(_04479_),
    .B1(_04478_),
    .Y(_04481_));
 sky130_fd_sc_hd__nor3_1 _11899_ (.A(_04477_),
    .B(_04480_),
    .C(_04481_),
    .Y(_04482_));
 sky130_fd_sc_hd__o21a_1 _11900_ (.A1(_04480_),
    .A2(_04481_),
    .B1(_04477_),
    .X(_04483_));
 sky130_fd_sc_hd__or4_4 _11901_ (.A(_04461_),
    .B(_04462_),
    .C(_04482_),
    .D(_04483_),
    .X(_04484_));
 sky130_fd_sc_hd__o22a_1 _11902_ (.A1(_04376_),
    .A2(_04377_),
    .B1(_04397_),
    .B2(_04398_),
    .X(_04485_));
 sky130_fd_sc_hd__a211oi_4 _11903_ (.A1(_04460_),
    .A2(_04484_),
    .B1(_04485_),
    .C1(_04399_),
    .Y(_04486_));
 sky130_fd_sc_hd__o211a_1 _11904_ (.A1(_04399_),
    .A2(_04485_),
    .B1(_04484_),
    .C1(_04460_),
    .X(_04487_));
 sky130_fd_sc_hd__a31o_1 _11905_ (.A1(_03491_),
    .A2(_03231_),
    .A3(_04474_),
    .B1(_04473_),
    .X(_04488_));
 sky130_fd_sc_hd__nand2_1 _11906_ (.A(_03948_),
    .B(_03234_),
    .Y(_04489_));
 sky130_fd_sc_hd__xnor2_1 _11907_ (.A(_04488_),
    .B(_04489_),
    .Y(_04490_));
 sky130_fd_sc_hd__and3_1 _11908_ (.A(_03947_),
    .B(_03281_),
    .C(_04490_),
    .X(_04491_));
 sky130_fd_sc_hd__a31o_1 _11909_ (.A1(_03943_),
    .A2(_03234_),
    .A3(_04488_),
    .B1(_04491_),
    .X(_04492_));
 sky130_fd_sc_hd__o21ba_1 _11910_ (.A1(_04477_),
    .A2(_04481_),
    .B1_N(_04480_),
    .X(_04493_));
 sky130_fd_sc_hd__a21oi_1 _11911_ (.A1(_03954_),
    .A2(_03231_),
    .B1(_04405_),
    .Y(_04494_));
 sky130_fd_sc_hd__nor2_1 _11912_ (.A(_04406_),
    .B(_04494_),
    .Y(_04495_));
 sky130_fd_sc_hd__xnor2_1 _11913_ (.A(_04493_),
    .B(_04495_),
    .Y(_04496_));
 sky130_fd_sc_hd__xnor2_1 _11914_ (.A(_04492_),
    .B(_04496_),
    .Y(_04497_));
 sky130_fd_sc_hd__nor3_1 _11915_ (.A(_04486_),
    .B(_04487_),
    .C(_04497_),
    .Y(_04498_));
 sky130_fd_sc_hd__o21ai_1 _11916_ (.A1(_04401_),
    .A2(_04402_),
    .B1(_04412_),
    .Y(_04499_));
 sky130_fd_sc_hd__or3_1 _11917_ (.A(_04401_),
    .B(_04402_),
    .C(_04412_),
    .X(_04500_));
 sky130_fd_sc_hd__o211a_1 _11918_ (.A1(_04486_),
    .A2(_04498_),
    .B1(_04499_),
    .C1(_04500_),
    .X(_04501_));
 sky130_fd_sc_hd__or3_1 _11919_ (.A(_04406_),
    .B(_04493_),
    .C(_04494_),
    .X(_04502_));
 sky130_fd_sc_hd__nand2_1 _11920_ (.A(_04492_),
    .B(_04496_),
    .Y(_04503_));
 sky130_fd_sc_hd__a211oi_1 _11921_ (.A1(_04500_),
    .A2(_04499_),
    .B1(_04498_),
    .C1(_04486_),
    .Y(_04504_));
 sky130_fd_sc_hd__a211oi_1 _11922_ (.A1(_04502_),
    .A2(_04503_),
    .B1(_04501_),
    .C1(_04504_),
    .Y(_04505_));
 sky130_fd_sc_hd__o211ai_1 _11923_ (.A1(_04419_),
    .A2(_04420_),
    .B1(_04417_),
    .C1(_04418_),
    .Y(_04506_));
 sky130_fd_sc_hd__o211a_1 _11924_ (.A1(_04501_),
    .A2(_04505_),
    .B1(_04421_),
    .C1(_04506_),
    .X(_04507_));
 sky130_fd_sc_hd__a211oi_1 _11925_ (.A1(_04421_),
    .A2(_04506_),
    .B1(_04501_),
    .C1(_04505_),
    .Y(_04508_));
 sky130_fd_sc_hd__or2_2 _11926_ (.A(_04507_),
    .B(_04508_),
    .X(_04509_));
 sky130_fd_sc_hd__o211a_1 _11927_ (.A1(_04501_),
    .A2(_04504_),
    .B1(_04502_),
    .C1(_04503_),
    .X(_04510_));
 sky130_fd_sc_hd__or2_2 _11928_ (.A(_04505_),
    .B(_04510_),
    .X(_04511_));
 sky130_fd_sc_hd__buf_4 _11929_ (.A(net28),
    .X(_04512_));
 sky130_fd_sc_hd__nand4_1 _11930_ (.A(_03014_),
    .B(_03019_),
    .C(_03684_),
    .D(_04512_),
    .Y(_04513_));
 sky130_fd_sc_hd__or3b_1 _11931_ (.A(_04351_),
    .B(_04513_),
    .C_N(_04430_),
    .X(_04514_));
 sky130_fd_sc_hd__nand4_2 _11932_ (.A(_04514_),
    .B(_04432_),
    .C(_04436_),
    .D(_04437_),
    .Y(_04515_));
 sky130_fd_sc_hd__a22o_1 _11933_ (.A1(_03596_),
    .A2(_03436_),
    .B1(_04512_),
    .B2(_03759_),
    .X(_04516_));
 sky130_fd_sc_hd__clkbuf_4 _11934_ (.A(net27),
    .X(_04517_));
 sky130_fd_sc_hd__and4_1 _11935_ (.A(_03678_),
    .B(_03679_),
    .C(net9),
    .D(_04517_),
    .X(_04518_));
 sky130_fd_sc_hd__a21o_1 _11936_ (.A1(_04513_),
    .A2(_04516_),
    .B1(_04518_),
    .X(_04519_));
 sky130_fd_sc_hd__buf_4 _11937_ (.A(_04270_),
    .X(_04520_));
 sky130_fd_sc_hd__and2_1 _11938_ (.A(_02948_),
    .B(_04520_),
    .X(_04521_));
 sky130_fd_sc_hd__buf_4 _11939_ (.A(net30),
    .X(_04522_));
 sky130_fd_sc_hd__a22o_1 _11940_ (.A1(_02955_),
    .A2(_04522_),
    .B1(_04426_),
    .B2(_02960_),
    .X(_04523_));
 sky130_fd_sc_hd__buf_4 _11941_ (.A(_04426_),
    .X(_04524_));
 sky130_fd_sc_hd__nand4_1 _11942_ (.A(_02960_),
    .B(_02955_),
    .C(_04522_),
    .D(_04524_),
    .Y(_04525_));
 sky130_fd_sc_hd__nand3_1 _11943_ (.A(_04521_),
    .B(_04523_),
    .C(_04525_),
    .Y(_04526_));
 sky130_fd_sc_hd__a21o_1 _11944_ (.A1(_04523_),
    .A2(_04525_),
    .B1(_04521_),
    .X(_04527_));
 sky130_fd_sc_hd__and3_1 _11945_ (.A(_04513_),
    .B(_04518_),
    .C(_04516_),
    .X(_04528_));
 sky130_fd_sc_hd__a31o_1 _11946_ (.A1(_04519_),
    .A2(_04526_),
    .A3(_04527_),
    .B1(_04528_),
    .X(_04529_));
 sky130_fd_sc_hd__a22o_1 _11947_ (.A1(_04514_),
    .A2(_04432_),
    .B1(_04436_),
    .B2(_04437_),
    .X(_04530_));
 sky130_fd_sc_hd__nand3_4 _11948_ (.A(_04515_),
    .B(_04529_),
    .C(_04530_),
    .Y(_04531_));
 sky130_fd_sc_hd__a21o_1 _11949_ (.A1(_04515_),
    .A2(_04530_),
    .B1(_04529_),
    .X(_04532_));
 sky130_fd_sc_hd__clkbuf_4 _11950_ (.A(_04185_),
    .X(_04533_));
 sky130_fd_sc_hd__nand4_1 _11951_ (.A(_02944_),
    .B(_02938_),
    .C(_04445_),
    .D(_04533_),
    .Y(_04534_));
 sky130_fd_sc_hd__buf_4 _11952_ (.A(_04444_),
    .X(_04535_));
 sky130_fd_sc_hd__a22o_1 _11953_ (.A1(_02938_),
    .A2(_04445_),
    .B1(_04533_),
    .B2(_03144_),
    .X(_04536_));
 sky130_fd_sc_hd__nand4_1 _11954_ (.A(_02935_),
    .B(_04535_),
    .C(_04534_),
    .D(_04536_),
    .Y(_04537_));
 sky130_fd_sc_hd__nand2_1 _11955_ (.A(_04534_),
    .B(_04537_),
    .Y(_04538_));
 sky130_fd_sc_hd__a21bo_1 _11956_ (.A1(_04521_),
    .A2(_04523_),
    .B1_N(_04525_),
    .X(_04539_));
 sky130_fd_sc_hd__a22o_1 _11957_ (.A1(_02935_),
    .A2(_04448_),
    .B1(_04446_),
    .B2(_04449_),
    .X(_04540_));
 sky130_fd_sc_hd__nand3_1 _11958_ (.A(_04450_),
    .B(_04539_),
    .C(_04540_),
    .Y(_04541_));
 sky130_fd_sc_hd__a21o_1 _11959_ (.A1(_04450_),
    .A2(_04540_),
    .B1(_04539_),
    .X(_04542_));
 sky130_fd_sc_hd__nand3_1 _11960_ (.A(_04538_),
    .B(_04541_),
    .C(_04542_),
    .Y(_04543_));
 sky130_fd_sc_hd__a21o_1 _11961_ (.A1(_04541_),
    .A2(_04542_),
    .B1(_04538_),
    .X(_04544_));
 sky130_fd_sc_hd__nand4_4 _11962_ (.A(_04531_),
    .B(_04532_),
    .C(_04543_),
    .D(_04544_),
    .Y(_04545_));
 sky130_fd_sc_hd__a22oi_4 _11963_ (.A1(_04442_),
    .A2(_04443_),
    .B1(_04456_),
    .B2(_04457_),
    .Y(_04546_));
 sky130_fd_sc_hd__a211oi_4 _11964_ (.A1(_04531_),
    .A2(_04545_),
    .B1(_04546_),
    .C1(_04458_),
    .Y(_04547_));
 sky130_fd_sc_hd__o211a_1 _11965_ (.A1(_04458_),
    .A2(_04546_),
    .B1(_04545_),
    .C1(_04531_),
    .X(_04548_));
 sky130_fd_sc_hd__nand3_1 _11966_ (.A(_04466_),
    .B(_04464_),
    .C(_04465_),
    .Y(_04549_));
 sky130_fd_sc_hd__and2_1 _11967_ (.A(_02926_),
    .B(_04286_),
    .X(_04550_));
 sky130_fd_sc_hd__buf_4 _11968_ (.A(_03770_),
    .X(_04551_));
 sky130_fd_sc_hd__a22o_1 _11969_ (.A1(_03213_),
    .A2(_04551_),
    .B1(_04447_),
    .B2(_03218_),
    .X(_04552_));
 sky130_fd_sc_hd__nand4_1 _11970_ (.A(_02921_),
    .B(_03213_),
    .C(_04551_),
    .D(_04447_),
    .Y(_04553_));
 sky130_fd_sc_hd__a21bo_1 _11971_ (.A1(_04550_),
    .A2(_04552_),
    .B1_N(_04553_),
    .X(_04554_));
 sky130_fd_sc_hd__clkbuf_4 _11972_ (.A(_03894_),
    .X(_04555_));
 sky130_fd_sc_hd__a22o_1 _11973_ (.A1(_02927_),
    .A2(_04555_),
    .B1(_04466_),
    .B2(_04465_),
    .X(_04556_));
 sky130_fd_sc_hd__nand3_1 _11974_ (.A(_04549_),
    .B(_04554_),
    .C(_04556_),
    .Y(_04557_));
 sky130_fd_sc_hd__a21o_1 _11975_ (.A1(_04549_),
    .A2(_04556_),
    .B1(_04554_),
    .X(_04558_));
 sky130_fd_sc_hd__nand2_1 _11976_ (.A(_03490_),
    .B(_03281_),
    .Y(_04559_));
 sky130_fd_sc_hd__and3_1 _11977_ (.A(_02894_),
    .B(_02896_),
    .C(_03597_),
    .X(_04560_));
 sky130_fd_sc_hd__a22o_1 _11978_ (.A1(_02896_),
    .A2(_03551_),
    .B1(_03675_),
    .B2(_02894_),
    .X(_04561_));
 sky130_fd_sc_hd__a21bo_1 _11979_ (.A1(_03685_),
    .A2(_04560_),
    .B1_N(_04561_),
    .X(_04562_));
 sky130_fd_sc_hd__xor2_1 _11980_ (.A(_04559_),
    .B(_04562_),
    .X(_04563_));
 sky130_fd_sc_hd__nand3_1 _11981_ (.A(_04557_),
    .B(_04558_),
    .C(_04563_),
    .Y(_04564_));
 sky130_fd_sc_hd__nand2_1 _11982_ (.A(_04557_),
    .B(_04564_),
    .Y(_04565_));
 sky130_fd_sc_hd__a21bo_1 _11983_ (.A1(_04538_),
    .A2(_04542_),
    .B1_N(_04541_),
    .X(_04566_));
 sky130_fd_sc_hd__a21o_1 _11984_ (.A1(_04469_),
    .A2(_04470_),
    .B1(_04475_),
    .X(_04567_));
 sky130_fd_sc_hd__nand3_1 _11985_ (.A(_04476_),
    .B(_04566_),
    .C(_04567_),
    .Y(_04568_));
 sky130_fd_sc_hd__a21o_1 _11986_ (.A1(_04476_),
    .A2(_04567_),
    .B1(_04566_),
    .X(_04569_));
 sky130_fd_sc_hd__and3_1 _11987_ (.A(_04565_),
    .B(_04568_),
    .C(_04569_),
    .X(_04570_));
 sky130_fd_sc_hd__a21oi_2 _11988_ (.A1(_04568_),
    .A2(_04569_),
    .B1(_04565_),
    .Y(_04571_));
 sky130_fd_sc_hd__nor4_4 _11989_ (.A(_04547_),
    .B(_04548_),
    .C(_04570_),
    .D(_04571_),
    .Y(_04572_));
 sky130_fd_sc_hd__o22ai_2 _11990_ (.A1(_04461_),
    .A2(_04462_),
    .B1(_04482_),
    .B2(_04483_),
    .Y(_04573_));
 sky130_fd_sc_hd__o211a_2 _11991_ (.A1(_04547_),
    .A2(_04572_),
    .B1(_04573_),
    .C1(_04484_),
    .X(_04574_));
 sky130_fd_sc_hd__a211oi_2 _11992_ (.A1(_04484_),
    .A2(_04573_),
    .B1(_04572_),
    .C1(_04547_),
    .Y(_04575_));
 sky130_fd_sc_hd__a32o_1 _11993_ (.A1(_03869_),
    .A2(_03281_),
    .A3(_04561_),
    .B1(_04560_),
    .B2(_03685_),
    .X(_04576_));
 sky130_fd_sc_hd__and3_1 _11994_ (.A(_03948_),
    .B(_03314_),
    .C(_04576_),
    .X(_04577_));
 sky130_fd_sc_hd__a21oi_1 _11995_ (.A1(_03942_),
    .A2(_03314_),
    .B1(_04576_),
    .Y(_04578_));
 sky130_fd_sc_hd__nor2_1 _11996_ (.A(_04577_),
    .B(_04578_),
    .Y(_04579_));
 sky130_fd_sc_hd__and3_1 _11997_ (.A(_03954_),
    .B(_03288_),
    .C(_04579_),
    .X(_04580_));
 sky130_fd_sc_hd__or2_1 _11998_ (.A(_04577_),
    .B(_04580_),
    .X(_04581_));
 sky130_fd_sc_hd__a21boi_2 _11999_ (.A1(_04565_),
    .A2(_04569_),
    .B1_N(_04568_),
    .Y(_04582_));
 sky130_fd_sc_hd__a21oi_1 _12000_ (.A1(_02908_),
    .A2(_03281_),
    .B1(_04490_),
    .Y(_04583_));
 sky130_fd_sc_hd__nor2_1 _12001_ (.A(_04491_),
    .B(_04583_),
    .Y(_04584_));
 sky130_fd_sc_hd__xnor2_1 _12002_ (.A(_04582_),
    .B(_04584_),
    .Y(_04585_));
 sky130_fd_sc_hd__xnor2_2 _12003_ (.A(_04581_),
    .B(_04585_),
    .Y(_04586_));
 sky130_fd_sc_hd__nor3_2 _12004_ (.A(_04574_),
    .B(_04575_),
    .C(_04586_),
    .Y(_04587_));
 sky130_fd_sc_hd__o21ai_2 _12005_ (.A1(_04486_),
    .A2(_04487_),
    .B1(_04497_),
    .Y(_04588_));
 sky130_fd_sc_hd__or3_1 _12006_ (.A(_04486_),
    .B(_04487_),
    .C(_04497_),
    .X(_04589_));
 sky130_fd_sc_hd__o211ai_4 _12007_ (.A1(_04574_),
    .A2(_04587_),
    .B1(_04588_),
    .C1(_04589_),
    .Y(_04590_));
 sky130_fd_sc_hd__inv_2 _12008_ (.A(_04590_),
    .Y(_04591_));
 sky130_fd_sc_hd__and2b_1 _12009_ (.A_N(_04582_),
    .B(_04584_),
    .X(_04592_));
 sky130_fd_sc_hd__and2_1 _12010_ (.A(_04581_),
    .B(_04585_),
    .X(_04593_));
 sky130_fd_sc_hd__a211o_1 _12011_ (.A1(_04589_),
    .A2(_04588_),
    .B1(_04587_),
    .C1(_04574_),
    .X(_04594_));
 sky130_fd_sc_hd__o211a_1 _12012_ (.A1(_04592_),
    .A2(_04593_),
    .B1(_04590_),
    .C1(_04594_),
    .X(_04595_));
 sky130_fd_sc_hd__nor2_1 _12013_ (.A(_04591_),
    .B(_04595_),
    .Y(_04596_));
 sky130_fd_sc_hd__xor2_2 _12014_ (.A(_04511_),
    .B(_04596_),
    .X(_04597_));
 sky130_fd_sc_hd__a211oi_1 _12015_ (.A1(_04590_),
    .A2(_04594_),
    .B1(_04592_),
    .C1(_04593_),
    .Y(_04598_));
 sky130_fd_sc_hd__nor2_1 _12016_ (.A(_04595_),
    .B(_04598_),
    .Y(_04599_));
 sky130_fd_sc_hd__nand3_1 _12017_ (.A(_04553_),
    .B(_04550_),
    .C(_04552_),
    .Y(_04600_));
 sky130_fd_sc_hd__and2_1 _12018_ (.A(_03529_),
    .B(_03771_),
    .X(_04601_));
 sky130_fd_sc_hd__a22o_1 _12019_ (.A1(_02922_),
    .A2(_04447_),
    .B1(_04444_),
    .B2(_02920_),
    .X(_04602_));
 sky130_fd_sc_hd__nand4_1 _12020_ (.A(_03208_),
    .B(_03210_),
    .C(_04447_),
    .D(_04444_),
    .Y(_04603_));
 sky130_fd_sc_hd__a21bo_1 _12021_ (.A1(_04601_),
    .A2(_04602_),
    .B1_N(_04603_),
    .X(_04604_));
 sky130_fd_sc_hd__a21o_1 _12022_ (.A1(_04553_),
    .A2(_04552_),
    .B1(_04550_),
    .X(_04605_));
 sky130_fd_sc_hd__nand3_1 _12023_ (.A(_04600_),
    .B(_04604_),
    .C(_04605_),
    .Y(_04606_));
 sky130_fd_sc_hd__a21o_1 _12024_ (.A1(_04600_),
    .A2(_04605_),
    .B1(_04604_),
    .X(_04607_));
 sky130_fd_sc_hd__nand2_1 _12025_ (.A(_03869_),
    .B(_03288_),
    .Y(_04608_));
 sky130_fd_sc_hd__a22o_1 _12026_ (.A1(_03873_),
    .A2(_03675_),
    .B1(_04555_),
    .B2(_03872_),
    .X(_04609_));
 sky130_fd_sc_hd__a21bo_1 _12027_ (.A1(_04555_),
    .A2(_04560_),
    .B1_N(_04609_),
    .X(_04610_));
 sky130_fd_sc_hd__xor2_1 _12028_ (.A(_04608_),
    .B(_04610_),
    .X(_04611_));
 sky130_fd_sc_hd__nand3_1 _12029_ (.A(_04606_),
    .B(_04607_),
    .C(_04611_),
    .Y(_04612_));
 sky130_fd_sc_hd__and2_1 _12030_ (.A(_04606_),
    .B(_04612_),
    .X(_04613_));
 sky130_fd_sc_hd__a21o_1 _12031_ (.A1(_04557_),
    .A2(_04558_),
    .B1(_04563_),
    .X(_04614_));
 sky130_fd_sc_hd__nand4_1 _12032_ (.A(_03144_),
    .B(_02938_),
    .C(_04533_),
    .D(_04520_),
    .Y(_04615_));
 sky130_fd_sc_hd__buf_4 _12033_ (.A(_04445_),
    .X(_04616_));
 sky130_fd_sc_hd__a22o_1 _12034_ (.A1(_03830_),
    .A2(_04185_),
    .B1(_04270_),
    .B2(_03799_),
    .X(_04617_));
 sky130_fd_sc_hd__nand4_1 _12035_ (.A(_02935_),
    .B(_04616_),
    .C(_04615_),
    .D(_04617_),
    .Y(_04618_));
 sky130_fd_sc_hd__nand2_1 _12036_ (.A(_04615_),
    .B(_04618_),
    .Y(_04619_));
 sky130_fd_sc_hd__a22o_1 _12037_ (.A1(_03798_),
    .A2(_04535_),
    .B1(_04534_),
    .B2(_04536_),
    .X(_04620_));
 sky130_fd_sc_hd__and2_1 _12038_ (.A(_02948_),
    .B(_04522_),
    .X(_04621_));
 sky130_fd_sc_hd__a22o_1 _12039_ (.A1(_02965_),
    .A2(_04426_),
    .B1(_04512_),
    .B2(_02963_),
    .X(_04622_));
 sky130_fd_sc_hd__nand4_1 _12040_ (.A(_02960_),
    .B(_02955_),
    .C(_04426_),
    .D(_04512_),
    .Y(_04623_));
 sky130_fd_sc_hd__a21bo_1 _12041_ (.A1(_04621_),
    .A2(_04622_),
    .B1_N(_04623_),
    .X(_04624_));
 sky130_fd_sc_hd__a21o_1 _12042_ (.A1(_04537_),
    .A2(_04620_),
    .B1(_04624_),
    .X(_04625_));
 sky130_fd_sc_hd__nand3_1 _12043_ (.A(_04537_),
    .B(_04624_),
    .C(_04620_),
    .Y(_04626_));
 sky130_fd_sc_hd__a21bo_1 _12044_ (.A1(_04619_),
    .A2(_04625_),
    .B1_N(_04626_),
    .X(_04627_));
 sky130_fd_sc_hd__a21oi_1 _12045_ (.A1(_04564_),
    .A2(_04614_),
    .B1(_04627_),
    .Y(_04628_));
 sky130_fd_sc_hd__and3_1 _12046_ (.A(_04564_),
    .B(_04627_),
    .C(_04614_),
    .X(_04629_));
 sky130_fd_sc_hd__o21ba_1 _12047_ (.A1(_04613_),
    .A2(_04628_),
    .B1_N(_04629_),
    .X(_04630_));
 sky130_fd_sc_hd__a21oi_1 _12048_ (.A1(_03959_),
    .A2(_03288_),
    .B1(_04579_),
    .Y(_04631_));
 sky130_fd_sc_hd__a32o_1 _12049_ (.A1(_03492_),
    .A2(_03288_),
    .A3(_04609_),
    .B1(_04560_),
    .B2(_04555_),
    .X(_04632_));
 sky130_fd_sc_hd__nand2_1 _12050_ (.A(_03942_),
    .B(_03231_),
    .Y(_04633_));
 sky130_fd_sc_hd__xnor2_1 _12051_ (.A(_04632_),
    .B(_04633_),
    .Y(_04634_));
 sky130_fd_sc_hd__and3_1 _12052_ (.A(_02908_),
    .B(_03437_),
    .C(_04634_),
    .X(_04635_));
 sky130_fd_sc_hd__a31o_1 _12053_ (.A1(_03944_),
    .A2(_03231_),
    .A3(_04632_),
    .B1(_04635_),
    .X(_04636_));
 sky130_fd_sc_hd__nor2_1 _12054_ (.A(_04580_),
    .B(_04631_),
    .Y(_04637_));
 sky130_fd_sc_hd__xnor2_1 _12055_ (.A(_04630_),
    .B(_04637_),
    .Y(_04638_));
 sky130_fd_sc_hd__nand2_1 _12056_ (.A(_04636_),
    .B(_04638_),
    .Y(_04639_));
 sky130_fd_sc_hd__o31a_1 _12057_ (.A1(_04580_),
    .A2(_04630_),
    .A3(_04631_),
    .B1(_04639_),
    .X(_04640_));
 sky130_fd_sc_hd__or3_1 _12058_ (.A(_04574_),
    .B(_04575_),
    .C(_04586_),
    .X(_04641_));
 sky130_fd_sc_hd__o21ai_1 _12059_ (.A1(_04574_),
    .A2(_04575_),
    .B1(_04586_),
    .Y(_04642_));
 sky130_fd_sc_hd__buf_4 _12060_ (.A(_04517_),
    .X(_04643_));
 sky130_fd_sc_hd__nand4_2 _12061_ (.A(_03014_),
    .B(_03019_),
    .C(_03551_),
    .D(_04643_),
    .Y(_04644_));
 sky130_fd_sc_hd__or3b_1 _12062_ (.A(_04431_),
    .B(_04644_),
    .C_N(_04516_),
    .X(_04645_));
 sky130_fd_sc_hd__nand4_1 _12063_ (.A(_04645_),
    .B(_04519_),
    .C(_04526_),
    .D(_04527_),
    .Y(_04646_));
 sky130_fd_sc_hd__a22o_1 _12064_ (.A1(_03679_),
    .A2(_03793_),
    .B1(_04517_),
    .B2(_03678_),
    .X(_04647_));
 sky130_fd_sc_hd__and4_1 _12065_ (.A(_03013_),
    .B(_03018_),
    .C(net8),
    .D(net26),
    .X(_04648_));
 sky130_fd_sc_hd__a21o_1 _12066_ (.A1(_04644_),
    .A2(_04647_),
    .B1(_04648_),
    .X(_04649_));
 sky130_fd_sc_hd__nand3_1 _12067_ (.A(_04621_),
    .B(_04623_),
    .C(_04622_),
    .Y(_04650_));
 sky130_fd_sc_hd__a21o_1 _12068_ (.A1(_04623_),
    .A2(_04622_),
    .B1(_04621_),
    .X(_04651_));
 sky130_fd_sc_hd__and3_1 _12069_ (.A(_04644_),
    .B(_04647_),
    .C(_04648_),
    .X(_04652_));
 sky130_fd_sc_hd__a31o_1 _12070_ (.A1(_04649_),
    .A2(_04650_),
    .A3(_04651_),
    .B1(_04652_),
    .X(_04653_));
 sky130_fd_sc_hd__a22o_1 _12071_ (.A1(_04645_),
    .A2(_04519_),
    .B1(_04526_),
    .B2(_04527_),
    .X(_04654_));
 sky130_fd_sc_hd__and3_2 _12072_ (.A(_04646_),
    .B(_04653_),
    .C(_04654_),
    .X(_04655_));
 sky130_fd_sc_hd__nand3_1 _12073_ (.A(_04646_),
    .B(_04653_),
    .C(_04654_),
    .Y(_04656_));
 sky130_fd_sc_hd__a21o_1 _12074_ (.A1(_04646_),
    .A2(_04654_),
    .B1(_04653_),
    .X(_04657_));
 sky130_fd_sc_hd__nand3_1 _12075_ (.A(_04619_),
    .B(_04626_),
    .C(_04625_),
    .Y(_04658_));
 sky130_fd_sc_hd__a21o_1 _12076_ (.A1(_04626_),
    .A2(_04625_),
    .B1(_04619_),
    .X(_04659_));
 sky130_fd_sc_hd__and4_2 _12077_ (.A(_04656_),
    .B(_04657_),
    .C(_04658_),
    .D(_04659_),
    .X(_04660_));
 sky130_fd_sc_hd__a22o_1 _12078_ (.A1(_04531_),
    .A2(_04532_),
    .B1(_04543_),
    .B2(_04544_),
    .X(_04661_));
 sky130_fd_sc_hd__o211ai_4 _12079_ (.A1(_04655_),
    .A2(_04660_),
    .B1(_04661_),
    .C1(_04545_),
    .Y(_04662_));
 sky130_fd_sc_hd__o211a_1 _12080_ (.A1(_04655_),
    .A2(_04660_),
    .B1(_04661_),
    .C1(_04545_),
    .X(_04663_));
 sky130_fd_sc_hd__a211oi_2 _12081_ (.A1(_04545_),
    .A2(_04661_),
    .B1(_04660_),
    .C1(_04655_),
    .Y(_04664_));
 sky130_fd_sc_hd__nor3_1 _12082_ (.A(_04613_),
    .B(_04629_),
    .C(_04628_),
    .Y(_04665_));
 sky130_fd_sc_hd__o21a_1 _12083_ (.A1(_04629_),
    .A2(_04628_),
    .B1(_04613_),
    .X(_04666_));
 sky130_fd_sc_hd__or4_4 _12084_ (.A(_04663_),
    .B(_04664_),
    .C(_04665_),
    .D(_04666_),
    .X(_04667_));
 sky130_fd_sc_hd__o22a_1 _12085_ (.A1(_04547_),
    .A2(_04548_),
    .B1(_04570_),
    .B2(_04571_),
    .X(_04668_));
 sky130_fd_sc_hd__a211oi_4 _12086_ (.A1(_04662_),
    .A2(_04667_),
    .B1(_04668_),
    .C1(_04572_),
    .Y(_04669_));
 sky130_fd_sc_hd__o211a_1 _12087_ (.A1(_04572_),
    .A2(_04668_),
    .B1(_04667_),
    .C1(_04662_),
    .X(_04670_));
 sky130_fd_sc_hd__xnor2_1 _12088_ (.A(_04636_),
    .B(_04638_),
    .Y(_04671_));
 sky130_fd_sc_hd__nor3_1 _12089_ (.A(_04669_),
    .B(_04670_),
    .C(_04671_),
    .Y(_04672_));
 sky130_fd_sc_hd__a211oi_2 _12090_ (.A1(_04641_),
    .A2(_04642_),
    .B1(_04672_),
    .C1(_04669_),
    .Y(_04673_));
 sky130_fd_sc_hd__o211a_1 _12091_ (.A1(_04669_),
    .A2(_04672_),
    .B1(_04642_),
    .C1(_04641_),
    .X(_04674_));
 sky130_fd_sc_hd__o21bai_2 _12092_ (.A1(_04640_),
    .A2(_04673_),
    .B1_N(_04674_),
    .Y(_04675_));
 sky130_fd_sc_hd__xor2_2 _12093_ (.A(_04599_),
    .B(_04675_),
    .X(_04676_));
 sky130_fd_sc_hd__or4bb_1 _12094_ (.A(_04425_),
    .B(_04509_),
    .C_N(_04597_),
    .D_N(_04676_),
    .X(_04677_));
 sky130_fd_sc_hd__or4_2 _12095_ (.A(_04183_),
    .B(_04264_),
    .C(_04345_),
    .D(_04677_),
    .X(_04678_));
 sky130_fd_sc_hd__nor3_1 _12096_ (.A(_04674_),
    .B(_04640_),
    .C(_04673_),
    .Y(_04679_));
 sky130_fd_sc_hd__o21a_1 _12097_ (.A1(_04674_),
    .A2(_04673_),
    .B1(_04640_),
    .X(_04680_));
 sky130_fd_sc_hd__buf_4 _12098_ (.A(net26),
    .X(_04681_));
 sky130_fd_sc_hd__nand4_1 _12099_ (.A(_03759_),
    .B(_03596_),
    .C(_03674_),
    .D(_04681_),
    .Y(_04682_));
 sky130_fd_sc_hd__or3b_1 _12100_ (.A(_04518_),
    .B(_04682_),
    .C_N(_04647_),
    .X(_04683_));
 sky130_fd_sc_hd__nand4_2 _12101_ (.A(_04683_),
    .B(_04649_),
    .C(_04650_),
    .D(_04651_),
    .Y(_04684_));
 sky130_fd_sc_hd__a22o_1 _12102_ (.A1(_03679_),
    .A2(_03674_),
    .B1(_04681_),
    .B2(_03678_),
    .X(_04685_));
 sky130_fd_sc_hd__clkbuf_4 _12103_ (.A(net23),
    .X(_04686_));
 sky130_fd_sc_hd__and4_1 _12104_ (.A(_03759_),
    .B(_03596_),
    .C(_03680_),
    .D(_04686_),
    .X(_04687_));
 sky130_fd_sc_hd__a21o_1 _12105_ (.A1(_04682_),
    .A2(_04685_),
    .B1(_04687_),
    .X(_04688_));
 sky130_fd_sc_hd__nand2_1 _12106_ (.A(_02948_),
    .B(_04426_),
    .Y(_04689_));
 sky130_fd_sc_hd__a22oi_2 _12107_ (.A1(_03773_),
    .A2(net28),
    .B1(_04517_),
    .B2(_02963_),
    .Y(_04690_));
 sky130_fd_sc_hd__and4_1 _12108_ (.A(_03774_),
    .B(_03773_),
    .C(net28),
    .D(_04517_),
    .X(_04691_));
 sky130_fd_sc_hd__or3_1 _12109_ (.A(_04689_),
    .B(_04690_),
    .C(_04691_),
    .X(_04692_));
 sky130_fd_sc_hd__o21ai_1 _12110_ (.A1(_04690_),
    .A2(_04691_),
    .B1(_04689_),
    .Y(_04693_));
 sky130_fd_sc_hd__and3_1 _12111_ (.A(_04682_),
    .B(_04687_),
    .C(_04685_),
    .X(_04694_));
 sky130_fd_sc_hd__a31o_1 _12112_ (.A1(_04688_),
    .A2(_04692_),
    .A3(_04693_),
    .B1(_04694_),
    .X(_04695_));
 sky130_fd_sc_hd__a22o_1 _12113_ (.A1(_04683_),
    .A2(_04649_),
    .B1(_04650_),
    .B2(_04651_),
    .X(_04696_));
 sky130_fd_sc_hd__nand3_4 _12114_ (.A(_04684_),
    .B(_04695_),
    .C(_04696_),
    .Y(_04697_));
 sky130_fd_sc_hd__a21o_1 _12115_ (.A1(_04684_),
    .A2(_04696_),
    .B1(_04695_),
    .X(_04698_));
 sky130_fd_sc_hd__and4_1 _12116_ (.A(_03143_),
    .B(_02937_),
    .C(_04270_),
    .D(_04346_),
    .X(_04699_));
 sky130_fd_sc_hd__nand2_1 _12117_ (.A(_02934_),
    .B(_04533_),
    .Y(_04700_));
 sky130_fd_sc_hd__a22oi_1 _12118_ (.A1(_02940_),
    .A2(_04270_),
    .B1(_04346_),
    .B2(_03799_),
    .Y(_04701_));
 sky130_fd_sc_hd__or3_1 _12119_ (.A(_04699_),
    .B(_04700_),
    .C(_04701_),
    .X(_04702_));
 sky130_fd_sc_hd__or2b_1 _12120_ (.A(_04699_),
    .B_N(_04702_),
    .X(_04703_));
 sky130_fd_sc_hd__o21bai_1 _12121_ (.A1(_04689_),
    .A2(_04690_),
    .B1_N(_04691_),
    .Y(_04704_));
 sky130_fd_sc_hd__a22o_1 _12122_ (.A1(_03798_),
    .A2(_04616_),
    .B1(_04615_),
    .B2(_04617_),
    .X(_04705_));
 sky130_fd_sc_hd__nand3_1 _12123_ (.A(_04618_),
    .B(_04704_),
    .C(_04705_),
    .Y(_04706_));
 sky130_fd_sc_hd__a21o_1 _12124_ (.A1(_04618_),
    .A2(_04705_),
    .B1(_04704_),
    .X(_04707_));
 sky130_fd_sc_hd__nand3_1 _12125_ (.A(_04703_),
    .B(_04706_),
    .C(_04707_),
    .Y(_04708_));
 sky130_fd_sc_hd__a21o_1 _12126_ (.A1(_04706_),
    .A2(_04707_),
    .B1(_04703_),
    .X(_04709_));
 sky130_fd_sc_hd__nand4_4 _12127_ (.A(_04697_),
    .B(_04698_),
    .C(_04708_),
    .D(_04709_),
    .Y(_04710_));
 sky130_fd_sc_hd__a22oi_4 _12128_ (.A1(_04656_),
    .A2(_04657_),
    .B1(_04658_),
    .B2(_04659_),
    .Y(_04711_));
 sky130_fd_sc_hd__a211oi_4 _12129_ (.A1(_04697_),
    .A2(_04710_),
    .B1(_04711_),
    .C1(_04660_),
    .Y(_04712_));
 sky130_fd_sc_hd__o211a_1 _12130_ (.A1(_04660_),
    .A2(_04711_),
    .B1(_04710_),
    .C1(_04697_),
    .X(_04713_));
 sky130_fd_sc_hd__nand3_1 _12131_ (.A(_04603_),
    .B(_04601_),
    .C(_04602_),
    .Y(_04714_));
 sky130_fd_sc_hd__nand2_1 _12132_ (.A(_03529_),
    .B(_04447_),
    .Y(_04715_));
 sky130_fd_sc_hd__a22oi_2 _12133_ (.A1(_02922_),
    .A2(_03760_),
    .B1(_04445_),
    .B2(_02920_),
    .Y(_04716_));
 sky130_fd_sc_hd__and4_1 _12134_ (.A(_03217_),
    .B(_03212_),
    .C(_03760_),
    .D(_04102_),
    .X(_04717_));
 sky130_fd_sc_hd__o21bai_1 _12135_ (.A1(_04715_),
    .A2(_04716_),
    .B1_N(_04717_),
    .Y(_04718_));
 sky130_fd_sc_hd__a22o_1 _12136_ (.A1(_02917_),
    .A2(_04551_),
    .B1(_04603_),
    .B2(_04602_),
    .X(_04719_));
 sky130_fd_sc_hd__nand3_1 _12137_ (.A(_04714_),
    .B(_04718_),
    .C(_04719_),
    .Y(_04720_));
 sky130_fd_sc_hd__a21o_1 _12138_ (.A1(_04714_),
    .A2(_04719_),
    .B1(_04718_),
    .X(_04721_));
 sky130_fd_sc_hd__nand2_1 _12139_ (.A(_03490_),
    .B(_03437_),
    .Y(_04722_));
 sky130_fd_sc_hd__a22oi_1 _12140_ (.A1(_03873_),
    .A2(_03894_),
    .B1(_04286_),
    .B2(_03872_),
    .Y(_04723_));
 sky130_fd_sc_hd__and4_1 _12141_ (.A(_03636_),
    .B(_03637_),
    .C(_03894_),
    .D(_03812_),
    .X(_04724_));
 sky130_fd_sc_hd__nor2_1 _12142_ (.A(_04723_),
    .B(_04724_),
    .Y(_04725_));
 sky130_fd_sc_hd__xnor2_1 _12143_ (.A(_04722_),
    .B(_04725_),
    .Y(_04726_));
 sky130_fd_sc_hd__nand3_1 _12144_ (.A(_04720_),
    .B(_04721_),
    .C(_04726_),
    .Y(_04727_));
 sky130_fd_sc_hd__nand2_1 _12145_ (.A(_04720_),
    .B(_04727_),
    .Y(_04728_));
 sky130_fd_sc_hd__a21bo_1 _12146_ (.A1(_04703_),
    .A2(_04707_),
    .B1_N(_04706_),
    .X(_04729_));
 sky130_fd_sc_hd__a21o_1 _12147_ (.A1(_04606_),
    .A2(_04607_),
    .B1(_04611_),
    .X(_04730_));
 sky130_fd_sc_hd__nand3_1 _12148_ (.A(_04612_),
    .B(_04729_),
    .C(_04730_),
    .Y(_04731_));
 sky130_fd_sc_hd__a21o_1 _12149_ (.A1(_04612_),
    .A2(_04730_),
    .B1(_04729_),
    .X(_04732_));
 sky130_fd_sc_hd__and3_1 _12150_ (.A(_04728_),
    .B(_04731_),
    .C(_04732_),
    .X(_04733_));
 sky130_fd_sc_hd__a21oi_2 _12151_ (.A1(_04731_),
    .A2(_04732_),
    .B1(_04728_),
    .Y(_04734_));
 sky130_fd_sc_hd__nor4_4 _12152_ (.A(_04712_),
    .B(_04713_),
    .C(_04733_),
    .D(_04734_),
    .Y(_04735_));
 sky130_fd_sc_hd__o22ai_2 _12153_ (.A1(_04663_),
    .A2(_04664_),
    .B1(_04665_),
    .B2(_04666_),
    .Y(_04736_));
 sky130_fd_sc_hd__o211a_1 _12154_ (.A1(_04712_),
    .A2(_04735_),
    .B1(_04736_),
    .C1(_04667_),
    .X(_04737_));
 sky130_fd_sc_hd__a211oi_2 _12155_ (.A1(_04667_),
    .A2(_04736_),
    .B1(_04735_),
    .C1(_04712_),
    .Y(_04738_));
 sky130_fd_sc_hd__a31o_1 _12156_ (.A1(_03492_),
    .A2(_03437_),
    .A3(_04725_),
    .B1(_04724_),
    .X(_04739_));
 sky130_fd_sc_hd__nand2_1 _12157_ (.A(_03942_),
    .B(_03281_),
    .Y(_04740_));
 sky130_fd_sc_hd__xnor2_1 _12158_ (.A(_04739_),
    .B(_04740_),
    .Y(_04741_));
 sky130_fd_sc_hd__and3_1 _12159_ (.A(_02908_),
    .B(_03685_),
    .C(_04741_),
    .X(_04742_));
 sky130_fd_sc_hd__a31o_1 _12160_ (.A1(_04081_),
    .A2(_03281_),
    .A3(_04739_),
    .B1(_04742_),
    .X(_04743_));
 sky130_fd_sc_hd__a21boi_1 _12161_ (.A1(_04728_),
    .A2(_04732_),
    .B1_N(_04731_),
    .Y(_04744_));
 sky130_fd_sc_hd__a21oi_1 _12162_ (.A1(_03959_),
    .A2(_03437_),
    .B1(_04634_),
    .Y(_04745_));
 sky130_fd_sc_hd__nor2_1 _12163_ (.A(_04635_),
    .B(_04745_),
    .Y(_04746_));
 sky130_fd_sc_hd__xnor2_1 _12164_ (.A(_04744_),
    .B(_04746_),
    .Y(_04747_));
 sky130_fd_sc_hd__xnor2_1 _12165_ (.A(_04743_),
    .B(_04747_),
    .Y(_04748_));
 sky130_fd_sc_hd__nor3_1 _12166_ (.A(_04737_),
    .B(_04738_),
    .C(_04748_),
    .Y(_04749_));
 sky130_fd_sc_hd__o21ai_1 _12167_ (.A1(_04669_),
    .A2(_04670_),
    .B1(_04671_),
    .Y(_04750_));
 sky130_fd_sc_hd__or3_1 _12168_ (.A(_04669_),
    .B(_04670_),
    .C(_04671_),
    .X(_04751_));
 sky130_fd_sc_hd__o211ai_1 _12169_ (.A1(_04737_),
    .A2(_04749_),
    .B1(_04750_),
    .C1(_04751_),
    .Y(_04752_));
 sky130_fd_sc_hd__or3_1 _12170_ (.A(_04635_),
    .B(_04744_),
    .C(_04745_),
    .X(_04753_));
 sky130_fd_sc_hd__nand2_1 _12171_ (.A(_04743_),
    .B(_04747_),
    .Y(_04754_));
 sky130_fd_sc_hd__o211a_1 _12172_ (.A1(_04737_),
    .A2(_04749_),
    .B1(_04750_),
    .C1(_04751_),
    .X(_04755_));
 sky130_fd_sc_hd__a211oi_1 _12173_ (.A1(_04751_),
    .A2(_04750_),
    .B1(_04749_),
    .C1(_04737_),
    .Y(_04756_));
 sky130_fd_sc_hd__a211o_1 _12174_ (.A1(_04753_),
    .A2(_04754_),
    .B1(_04755_),
    .C1(_04756_),
    .X(_04757_));
 sky130_fd_sc_hd__o211a_1 _12175_ (.A1(_04679_),
    .A2(_04680_),
    .B1(_04752_),
    .C1(_04757_),
    .X(_04758_));
 sky130_fd_sc_hd__a211oi_1 _12176_ (.A1(_04752_),
    .A2(_04757_),
    .B1(_04679_),
    .C1(_04680_),
    .Y(_04759_));
 sky130_fd_sc_hd__nor2_2 _12177_ (.A(_04758_),
    .B(_04759_),
    .Y(_04760_));
 sky130_fd_sc_hd__nand4_2 _12178_ (.A(_03013_),
    .B(_03018_),
    .C(net7),
    .D(net23),
    .Y(_04761_));
 sky130_fd_sc_hd__or3b_1 _12179_ (.A(_04648_),
    .B(_04761_),
    .C_N(_04685_),
    .X(_04762_));
 sky130_fd_sc_hd__nand4_1 _12180_ (.A(_04762_),
    .B(_04688_),
    .C(_04692_),
    .D(_04693_),
    .Y(_04763_));
 sky130_fd_sc_hd__a22o_1 _12181_ (.A1(_03757_),
    .A2(net7),
    .B1(net23),
    .B2(_03756_),
    .X(_04764_));
 sky130_fd_sc_hd__and4_1 _12182_ (.A(\wfg_stim_mem_top.cfg_gain_q[23] ),
    .B(\wfg_stim_mem_top.cfg_gain_q[10] ),
    .C(net6),
    .D(net12),
    .X(_04765_));
 sky130_fd_sc_hd__a21o_1 _12183_ (.A1(_04761_),
    .A2(_04764_),
    .B1(_04765_),
    .X(_04766_));
 sky130_fd_sc_hd__and2_1 _12184_ (.A(\wfg_stim_mem_top.cfg_gain_q[20] ),
    .B(net28),
    .X(_04767_));
 sky130_fd_sc_hd__nand4_1 _12185_ (.A(_02963_),
    .B(_02965_),
    .C(_04517_),
    .D(_04681_),
    .Y(_04768_));
 sky130_fd_sc_hd__a22o_1 _12186_ (.A1(_03773_),
    .A2(net27),
    .B1(_04681_),
    .B2(_03774_),
    .X(_04769_));
 sky130_fd_sc_hd__nand3_1 _12187_ (.A(_04767_),
    .B(_04768_),
    .C(_04769_),
    .Y(_04770_));
 sky130_fd_sc_hd__a21o_1 _12188_ (.A1(_04768_),
    .A2(_04769_),
    .B1(_04767_),
    .X(_04771_));
 sky130_fd_sc_hd__and3_1 _12189_ (.A(_04761_),
    .B(_04765_),
    .C(_04764_),
    .X(_04772_));
 sky130_fd_sc_hd__a31o_1 _12190_ (.A1(_04766_),
    .A2(_04770_),
    .A3(_04771_),
    .B1(_04772_),
    .X(_04773_));
 sky130_fd_sc_hd__a22o_1 _12191_ (.A1(_04762_),
    .A2(_04688_),
    .B1(_04692_),
    .B2(_04693_),
    .X(_04774_));
 sky130_fd_sc_hd__and3_2 _12192_ (.A(_04763_),
    .B(_04773_),
    .C(_04774_),
    .X(_04775_));
 sky130_fd_sc_hd__nand3_2 _12193_ (.A(_04763_),
    .B(_04773_),
    .C(_04774_),
    .Y(_04776_));
 sky130_fd_sc_hd__a21o_1 _12194_ (.A1(_04763_),
    .A2(_04774_),
    .B1(_04773_),
    .X(_04777_));
 sky130_fd_sc_hd__nand4_2 _12195_ (.A(_03799_),
    .B(_03830_),
    .C(_04346_),
    .D(_04426_),
    .Y(_04778_));
 sky130_fd_sc_hd__a22o_1 _12196_ (.A1(_02940_),
    .A2(_04346_),
    .B1(_04426_),
    .B2(_02943_),
    .X(_04779_));
 sky130_fd_sc_hd__nand4_2 _12197_ (.A(_03798_),
    .B(_04520_),
    .C(_04778_),
    .D(_04779_),
    .Y(_04780_));
 sky130_fd_sc_hd__nand2_1 _12198_ (.A(_04778_),
    .B(_04780_),
    .Y(_04781_));
 sky130_fd_sc_hd__a21bo_1 _12199_ (.A1(_04767_),
    .A2(_04769_),
    .B1_N(_04768_),
    .X(_04782_));
 sky130_fd_sc_hd__o21ai_1 _12200_ (.A1(_04699_),
    .A2(_04701_),
    .B1(_04700_),
    .Y(_04783_));
 sky130_fd_sc_hd__nand3_1 _12201_ (.A(_04702_),
    .B(_04782_),
    .C(_04783_),
    .Y(_04784_));
 sky130_fd_sc_hd__a21o_1 _12202_ (.A1(_04702_),
    .A2(_04783_),
    .B1(_04782_),
    .X(_04785_));
 sky130_fd_sc_hd__nand3_1 _12203_ (.A(_04781_),
    .B(_04784_),
    .C(_04785_),
    .Y(_04786_));
 sky130_fd_sc_hd__a21o_1 _12204_ (.A1(_04784_),
    .A2(_04785_),
    .B1(_04781_),
    .X(_04787_));
 sky130_fd_sc_hd__and4_4 _12205_ (.A(_04776_),
    .B(_04777_),
    .C(_04786_),
    .D(_04787_),
    .X(_04788_));
 sky130_fd_sc_hd__a22o_2 _12206_ (.A1(_04697_),
    .A2(_04698_),
    .B1(_04708_),
    .B2(_04709_),
    .X(_04789_));
 sky130_fd_sc_hd__o211ai_4 _12207_ (.A1(_04775_),
    .A2(_04788_),
    .B1(_04789_),
    .C1(_04710_),
    .Y(_04790_));
 sky130_fd_sc_hd__o211a_1 _12208_ (.A1(_04775_),
    .A2(_04788_),
    .B1(_04789_),
    .C1(_04710_),
    .X(_04791_));
 sky130_fd_sc_hd__a211oi_2 _12209_ (.A1(_04710_),
    .A2(_04789_),
    .B1(_04788_),
    .C1(_04775_),
    .Y(_04792_));
 sky130_fd_sc_hd__or3_1 _12210_ (.A(_04717_),
    .B(_04715_),
    .C(_04716_),
    .X(_04793_));
 sky130_fd_sc_hd__and2_1 _12211_ (.A(\wfg_stim_mem_top.cfg_gain_q[14] ),
    .B(_04444_),
    .X(_04794_));
 sky130_fd_sc_hd__a22o_1 _12212_ (.A1(_03209_),
    .A2(_04102_),
    .B1(_04185_),
    .B2(_02919_),
    .X(_04795_));
 sky130_fd_sc_hd__nand4_1 _12213_ (.A(_02920_),
    .B(_02922_),
    .C(_04102_),
    .D(_04533_),
    .Y(_04796_));
 sky130_fd_sc_hd__a21bo_1 _12214_ (.A1(_04794_),
    .A2(_04795_),
    .B1_N(_04796_),
    .X(_04797_));
 sky130_fd_sc_hd__o21ai_1 _12215_ (.A1(_04717_),
    .A2(_04716_),
    .B1(_04715_),
    .Y(_04798_));
 sky130_fd_sc_hd__nand3_1 _12216_ (.A(_04793_),
    .B(_04797_),
    .C(_04798_),
    .Y(_04799_));
 sky130_fd_sc_hd__a21o_1 _12217_ (.A1(_04793_),
    .A2(_04798_),
    .B1(_04797_),
    .X(_04800_));
 sky130_fd_sc_hd__nand2_1 _12218_ (.A(_03490_),
    .B(_03685_),
    .Y(_04801_));
 sky130_fd_sc_hd__a22oi_1 _12219_ (.A1(_03873_),
    .A2(_04286_),
    .B1(_04551_),
    .B2(_03872_),
    .Y(_04802_));
 sky130_fd_sc_hd__and4_1 _12220_ (.A(_03636_),
    .B(_03637_),
    .C(_03812_),
    .D(_03771_),
    .X(_04803_));
 sky130_fd_sc_hd__nor2_1 _12221_ (.A(_04802_),
    .B(_04803_),
    .Y(_04804_));
 sky130_fd_sc_hd__xnor2_2 _12222_ (.A(_04801_),
    .B(_04804_),
    .Y(_04805_));
 sky130_fd_sc_hd__nand3_1 _12223_ (.A(_04799_),
    .B(_04800_),
    .C(_04805_),
    .Y(_04806_));
 sky130_fd_sc_hd__and2_1 _12224_ (.A(_04799_),
    .B(_04806_),
    .X(_04807_));
 sky130_fd_sc_hd__a21bo_1 _12225_ (.A1(_04781_),
    .A2(_04785_),
    .B1_N(_04784_),
    .X(_04808_));
 sky130_fd_sc_hd__a21o_1 _12226_ (.A1(_04720_),
    .A2(_04721_),
    .B1(_04726_),
    .X(_04809_));
 sky130_fd_sc_hd__and3_1 _12227_ (.A(_04727_),
    .B(_04808_),
    .C(_04809_),
    .X(_04810_));
 sky130_fd_sc_hd__a21oi_1 _12228_ (.A1(_04727_),
    .A2(_04809_),
    .B1(_04808_),
    .Y(_04811_));
 sky130_fd_sc_hd__nor3_1 _12229_ (.A(_04807_),
    .B(_04810_),
    .C(_04811_),
    .Y(_04812_));
 sky130_fd_sc_hd__o21a_1 _12230_ (.A1(_04810_),
    .A2(_04811_),
    .B1(_04807_),
    .X(_04813_));
 sky130_fd_sc_hd__or4_4 _12231_ (.A(_04791_),
    .B(_04792_),
    .C(_04812_),
    .D(_04813_),
    .X(_04814_));
 sky130_fd_sc_hd__o22a_1 _12232_ (.A1(_04712_),
    .A2(_04713_),
    .B1(_04733_),
    .B2(_04734_),
    .X(_04815_));
 sky130_fd_sc_hd__a211oi_4 _12233_ (.A1(_04790_),
    .A2(_04814_),
    .B1(_04815_),
    .C1(_04735_),
    .Y(_04816_));
 sky130_fd_sc_hd__o211a_1 _12234_ (.A1(_04735_),
    .A2(_04815_),
    .B1(_04814_),
    .C1(_04790_),
    .X(_04817_));
 sky130_fd_sc_hd__a31o_1 _12235_ (.A1(_03945_),
    .A2(_03685_),
    .A3(_04804_),
    .B1(_04803_),
    .X(_04818_));
 sky130_fd_sc_hd__nand2_1 _12236_ (.A(_03948_),
    .B(_03288_),
    .Y(_04819_));
 sky130_fd_sc_hd__xnor2_1 _12237_ (.A(_04818_),
    .B(_04819_),
    .Y(_04820_));
 sky130_fd_sc_hd__and3_1 _12238_ (.A(_03947_),
    .B(_03675_),
    .C(_04820_),
    .X(_04821_));
 sky130_fd_sc_hd__a31o_1 _12239_ (.A1(_04081_),
    .A2(_03288_),
    .A3(_04818_),
    .B1(_04821_),
    .X(_04822_));
 sky130_fd_sc_hd__o21ba_1 _12240_ (.A1(_04807_),
    .A2(_04811_),
    .B1_N(_04810_),
    .X(_04823_));
 sky130_fd_sc_hd__a21oi_1 _12241_ (.A1(_03959_),
    .A2(_03685_),
    .B1(_04741_),
    .Y(_04824_));
 sky130_fd_sc_hd__nor2_1 _12242_ (.A(_04742_),
    .B(_04824_),
    .Y(_04825_));
 sky130_fd_sc_hd__xnor2_1 _12243_ (.A(_04823_),
    .B(_04825_),
    .Y(_04826_));
 sky130_fd_sc_hd__xnor2_1 _12244_ (.A(_04822_),
    .B(_04826_),
    .Y(_04827_));
 sky130_fd_sc_hd__nor3_1 _12245_ (.A(_04816_),
    .B(_04817_),
    .C(_04827_),
    .Y(_04828_));
 sky130_fd_sc_hd__o21ai_1 _12246_ (.A1(_04737_),
    .A2(_04738_),
    .B1(_04748_),
    .Y(_04829_));
 sky130_fd_sc_hd__or3_1 _12247_ (.A(_04737_),
    .B(_04738_),
    .C(_04748_),
    .X(_04830_));
 sky130_fd_sc_hd__o211a_1 _12248_ (.A1(_04816_),
    .A2(_04828_),
    .B1(_04829_),
    .C1(_04830_),
    .X(_04831_));
 sky130_fd_sc_hd__or3_1 _12249_ (.A(_04742_),
    .B(_04823_),
    .C(_04824_),
    .X(_04832_));
 sky130_fd_sc_hd__nand2_1 _12250_ (.A(_04822_),
    .B(_04826_),
    .Y(_04833_));
 sky130_fd_sc_hd__a211oi_2 _12251_ (.A1(_04830_),
    .A2(_04829_),
    .B1(_04828_),
    .C1(_04816_),
    .Y(_04834_));
 sky130_fd_sc_hd__a211oi_1 _12252_ (.A1(_04832_),
    .A2(_04833_),
    .B1(_04831_),
    .C1(_04834_),
    .Y(_04835_));
 sky130_fd_sc_hd__o211ai_1 _12253_ (.A1(_04755_),
    .A2(_04756_),
    .B1(_04753_),
    .C1(_04754_),
    .Y(_04836_));
 sky130_fd_sc_hd__o211a_1 _12254_ (.A1(_04831_),
    .A2(_04835_),
    .B1(_04757_),
    .C1(_04836_),
    .X(_04837_));
 sky130_fd_sc_hd__a211o_1 _12255_ (.A1(_04757_),
    .A2(_04836_),
    .B1(_04831_),
    .C1(_04835_),
    .X(_04838_));
 sky130_fd_sc_hd__nor2b_4 _12256_ (.A(_04837_),
    .B_N(_04838_),
    .Y(_04839_));
 sky130_fd_sc_hd__a211o_1 _12257_ (.A1(_04832_),
    .A2(_04833_),
    .B1(_04831_),
    .C1(_04834_),
    .X(_04840_));
 sky130_fd_sc_hd__o211ai_2 _12258_ (.A1(_04831_),
    .A2(_04834_),
    .B1(_04832_),
    .C1(_04833_),
    .Y(_04841_));
 sky130_fd_sc_hd__a21oi_1 _12259_ (.A1(_04761_),
    .A2(_04764_),
    .B1(_04765_),
    .Y(_04842_));
 sky130_fd_sc_hd__or4bb_2 _12260_ (.A(_04772_),
    .B(_04842_),
    .C_N(_04770_),
    .D_N(_04771_),
    .X(_04843_));
 sky130_fd_sc_hd__nand4_1 _12261_ (.A(_03013_),
    .B(_03018_),
    .C(_03769_),
    .D(net12),
    .Y(_04844_));
 sky130_fd_sc_hd__a22o_1 _12262_ (.A1(\wfg_stim_mem_top.cfg_gain_q[10] ),
    .A2(net6),
    .B1(net12),
    .B2(\wfg_stim_mem_top.cfg_gain_q[23] ),
    .X(_04845_));
 sky130_fd_sc_hd__and4_1 _12263_ (.A(\wfg_stim_mem_top.cfg_gain_q[23] ),
    .B(\wfg_stim_mem_top.cfg_gain_q[10] ),
    .C(net5),
    .D(net1),
    .X(_04846_));
 sky130_fd_sc_hd__a21o_1 _12264_ (.A1(_04844_),
    .A2(_04845_),
    .B1(_04846_),
    .X(_04847_));
 sky130_fd_sc_hd__nand2_1 _12265_ (.A(\wfg_stim_mem_top.cfg_gain_q[20] ),
    .B(net27),
    .Y(_04848_));
 sky130_fd_sc_hd__and4_1 _12266_ (.A(_02959_),
    .B(\wfg_stim_mem_top.cfg_gain_q[21] ),
    .C(net26),
    .D(net23),
    .X(_04849_));
 sky130_fd_sc_hd__a22oi_2 _12267_ (.A1(_02954_),
    .A2(net26),
    .B1(net23),
    .B2(_02959_),
    .Y(_04850_));
 sky130_fd_sc_hd__or3_1 _12268_ (.A(_04848_),
    .B(_04849_),
    .C(_04850_),
    .X(_04851_));
 sky130_fd_sc_hd__o21ai_1 _12269_ (.A1(_04849_),
    .A2(_04850_),
    .B1(_04848_),
    .Y(_04852_));
 sky130_fd_sc_hd__and3_1 _12270_ (.A(_04844_),
    .B(_04846_),
    .C(_04845_),
    .X(_04853_));
 sky130_fd_sc_hd__a31o_1 _12271_ (.A1(_04847_),
    .A2(_04851_),
    .A3(_04852_),
    .B1(_04853_),
    .X(_04854_));
 sky130_fd_sc_hd__a2bb2o_1 _12272_ (.A1_N(_04772_),
    .A2_N(_04842_),
    .B1(_04770_),
    .B2(_04771_),
    .X(_04855_));
 sky130_fd_sc_hd__nand3_4 _12273_ (.A(_04843_),
    .B(_04854_),
    .C(_04855_),
    .Y(_04856_));
 sky130_fd_sc_hd__a21o_1 _12274_ (.A1(_04843_),
    .A2(_04855_),
    .B1(_04854_),
    .X(_04857_));
 sky130_fd_sc_hd__and4_1 _12275_ (.A(_03143_),
    .B(\wfg_stim_mem_top.cfg_gain_q[18] ),
    .C(net29),
    .D(net28),
    .X(_04858_));
 sky130_fd_sc_hd__nand2_1 _12276_ (.A(\wfg_stim_mem_top.cfg_gain_q[17] ),
    .B(_04346_),
    .Y(_04859_));
 sky130_fd_sc_hd__a22oi_1 _12277_ (.A1(_02937_),
    .A2(net29),
    .B1(net28),
    .B2(_02943_),
    .Y(_04860_));
 sky130_fd_sc_hd__or3_1 _12278_ (.A(_04858_),
    .B(_04859_),
    .C(_04860_),
    .X(_04861_));
 sky130_fd_sc_hd__or2b_1 _12279_ (.A(_04858_),
    .B_N(_04861_),
    .X(_04862_));
 sky130_fd_sc_hd__o21bai_1 _12280_ (.A1(_04848_),
    .A2(_04850_),
    .B1_N(_04849_),
    .Y(_04863_));
 sky130_fd_sc_hd__a22o_1 _12281_ (.A1(_02934_),
    .A2(_04520_),
    .B1(_04778_),
    .B2(_04779_),
    .X(_04864_));
 sky130_fd_sc_hd__nand3_1 _12282_ (.A(_04780_),
    .B(_04863_),
    .C(_04864_),
    .Y(_04865_));
 sky130_fd_sc_hd__a21o_1 _12283_ (.A1(_04780_),
    .A2(_04864_),
    .B1(_04863_),
    .X(_04866_));
 sky130_fd_sc_hd__nand3_1 _12284_ (.A(_04862_),
    .B(_04865_),
    .C(_04866_),
    .Y(_04867_));
 sky130_fd_sc_hd__a21o_1 _12285_ (.A1(_04865_),
    .A2(_04866_),
    .B1(_04862_),
    .X(_04868_));
 sky130_fd_sc_hd__nand4_4 _12286_ (.A(_04856_),
    .B(_04857_),
    .C(_04867_),
    .D(_04868_),
    .Y(_04869_));
 sky130_fd_sc_hd__a22oi_4 _12287_ (.A1(_04776_),
    .A2(_04777_),
    .B1(_04786_),
    .B2(_04787_),
    .Y(_04870_));
 sky130_fd_sc_hd__a211oi_4 _12288_ (.A1(_04856_),
    .A2(_04869_),
    .B1(_04870_),
    .C1(_04788_),
    .Y(_04871_));
 sky130_fd_sc_hd__o211a_1 _12289_ (.A1(_04788_),
    .A2(_04870_),
    .B1(_04869_),
    .C1(_04856_),
    .X(_04872_));
 sky130_fd_sc_hd__nand3_1 _12290_ (.A(_04796_),
    .B(_04794_),
    .C(_04795_),
    .Y(_04873_));
 sky130_fd_sc_hd__nand2_1 _12291_ (.A(_03529_),
    .B(_04445_),
    .Y(_04874_));
 sky130_fd_sc_hd__a22oi_2 _12292_ (.A1(_02922_),
    .A2(_04533_),
    .B1(_04520_),
    .B2(_02920_),
    .Y(_04875_));
 sky130_fd_sc_hd__and4_1 _12293_ (.A(_02919_),
    .B(_03209_),
    .C(_04185_),
    .D(_04270_),
    .X(_04876_));
 sky130_fd_sc_hd__o21bai_1 _12294_ (.A1(_04874_),
    .A2(_04875_),
    .B1_N(_04876_),
    .Y(_04877_));
 sky130_fd_sc_hd__a22o_1 _12295_ (.A1(_02926_),
    .A2(_04444_),
    .B1(_04796_),
    .B2(_04795_),
    .X(_04878_));
 sky130_fd_sc_hd__nand3_1 _12296_ (.A(_04873_),
    .B(_04877_),
    .C(_04878_),
    .Y(_04879_));
 sky130_fd_sc_hd__a21o_1 _12297_ (.A1(_04873_),
    .A2(_04878_),
    .B1(_04877_),
    .X(_04880_));
 sky130_fd_sc_hd__nand2_1 _12298_ (.A(_02892_),
    .B(_03675_),
    .Y(_04881_));
 sky130_fd_sc_hd__a22oi_1 _12299_ (.A1(_03637_),
    .A2(_03771_),
    .B1(_04447_),
    .B2(_03636_),
    .Y(_04882_));
 sky130_fd_sc_hd__and4_1 _12300_ (.A(\wfg_stim_mem_top.cfg_gain_q[13] ),
    .B(\wfg_stim_mem_top.cfg_gain_q[12] ),
    .C(_03771_),
    .D(_04447_),
    .X(_04883_));
 sky130_fd_sc_hd__nor2_1 _12301_ (.A(_04882_),
    .B(_04883_),
    .Y(_04884_));
 sky130_fd_sc_hd__xnor2_2 _12302_ (.A(_04881_),
    .B(_04884_),
    .Y(_04885_));
 sky130_fd_sc_hd__nand3_1 _12303_ (.A(_04879_),
    .B(_04880_),
    .C(_04885_),
    .Y(_04886_));
 sky130_fd_sc_hd__nand2_1 _12304_ (.A(_04879_),
    .B(_04886_),
    .Y(_04887_));
 sky130_fd_sc_hd__a21bo_1 _12305_ (.A1(_04862_),
    .A2(_04866_),
    .B1_N(_04865_),
    .X(_04888_));
 sky130_fd_sc_hd__a21o_1 _12306_ (.A1(_04799_),
    .A2(_04800_),
    .B1(_04805_),
    .X(_04889_));
 sky130_fd_sc_hd__nand3_1 _12307_ (.A(_04806_),
    .B(_04888_),
    .C(_04889_),
    .Y(_04890_));
 sky130_fd_sc_hd__a21o_1 _12308_ (.A1(_04806_),
    .A2(_04889_),
    .B1(_04888_),
    .X(_04891_));
 sky130_fd_sc_hd__and3_1 _12309_ (.A(_04887_),
    .B(_04890_),
    .C(_04891_),
    .X(_04892_));
 sky130_fd_sc_hd__a21oi_2 _12310_ (.A1(_04890_),
    .A2(_04891_),
    .B1(_04887_),
    .Y(_04893_));
 sky130_fd_sc_hd__nor4_4 _12311_ (.A(_04871_),
    .B(_04872_),
    .C(_04892_),
    .D(_04893_),
    .Y(_04894_));
 sky130_fd_sc_hd__o22ai_2 _12312_ (.A1(_04791_),
    .A2(_04792_),
    .B1(_04812_),
    .B2(_04813_),
    .Y(_04895_));
 sky130_fd_sc_hd__o211a_1 _12313_ (.A1(_04871_),
    .A2(_04894_),
    .B1(_04895_),
    .C1(_04814_),
    .X(_04896_));
 sky130_fd_sc_hd__a211oi_2 _12314_ (.A1(_04814_),
    .A2(_04895_),
    .B1(_04894_),
    .C1(_04871_),
    .Y(_04897_));
 sky130_fd_sc_hd__a31o_1 _12315_ (.A1(_03491_),
    .A2(_03675_),
    .A3(_04884_),
    .B1(_04883_),
    .X(_04898_));
 sky130_fd_sc_hd__nand2_1 _12316_ (.A(_02887_),
    .B(_03437_),
    .Y(_04899_));
 sky130_fd_sc_hd__xnor2_1 _12317_ (.A(_04898_),
    .B(_04899_),
    .Y(_04900_));
 sky130_fd_sc_hd__and3_1 _12318_ (.A(_02907_),
    .B(_04555_),
    .C(_04900_),
    .X(_04901_));
 sky130_fd_sc_hd__a31o_1 _12319_ (.A1(_03944_),
    .A2(_03437_),
    .A3(_04898_),
    .B1(_04901_),
    .X(_04902_));
 sky130_fd_sc_hd__a21boi_1 _12320_ (.A1(_04887_),
    .A2(_04891_),
    .B1_N(_04890_),
    .Y(_04903_));
 sky130_fd_sc_hd__a21oi_1 _12321_ (.A1(_02908_),
    .A2(_03675_),
    .B1(_04820_),
    .Y(_04904_));
 sky130_fd_sc_hd__nor2_1 _12322_ (.A(_04821_),
    .B(_04904_),
    .Y(_04905_));
 sky130_fd_sc_hd__xnor2_1 _12323_ (.A(_04903_),
    .B(_04905_),
    .Y(_04906_));
 sky130_fd_sc_hd__xnor2_1 _12324_ (.A(_04902_),
    .B(_04906_),
    .Y(_04907_));
 sky130_fd_sc_hd__nor3_1 _12325_ (.A(_04896_),
    .B(_04897_),
    .C(_04907_),
    .Y(_04908_));
 sky130_fd_sc_hd__o21ai_1 _12326_ (.A1(_04816_),
    .A2(_04817_),
    .B1(_04827_),
    .Y(_04909_));
 sky130_fd_sc_hd__or3_1 _12327_ (.A(_04816_),
    .B(_04817_),
    .C(_04827_),
    .X(_04910_));
 sky130_fd_sc_hd__o211a_1 _12328_ (.A1(_04896_),
    .A2(_04908_),
    .B1(_04909_),
    .C1(_04910_),
    .X(_04911_));
 sky130_fd_sc_hd__and2b_1 _12329_ (.A_N(_04903_),
    .B(_04905_),
    .X(_04912_));
 sky130_fd_sc_hd__and2_1 _12330_ (.A(_04902_),
    .B(_04906_),
    .X(_04913_));
 sky130_fd_sc_hd__o211ai_1 _12331_ (.A1(_04896_),
    .A2(_04908_),
    .B1(_04909_),
    .C1(_04910_),
    .Y(_04914_));
 sky130_fd_sc_hd__a211o_1 _12332_ (.A1(_04910_),
    .A2(_04909_),
    .B1(_04908_),
    .C1(_04896_),
    .X(_04915_));
 sky130_fd_sc_hd__o211a_1 _12333_ (.A1(_04912_),
    .A2(_04913_),
    .B1(_04914_),
    .C1(_04915_),
    .X(_04916_));
 sky130_fd_sc_hd__a211oi_2 _12334_ (.A1(_04840_),
    .A2(_04841_),
    .B1(_04911_),
    .C1(_04916_),
    .Y(_04917_));
 sky130_fd_sc_hd__o211a_1 _12335_ (.A1(_04911_),
    .A2(_04916_),
    .B1(_04840_),
    .C1(_04841_),
    .X(_04918_));
 sky130_fd_sc_hd__nor2_4 _12336_ (.A(_04917_),
    .B(_04918_),
    .Y(_04919_));
 sky130_fd_sc_hd__a211oi_2 _12337_ (.A1(_04914_),
    .A2(_04915_),
    .B1(_04912_),
    .C1(_04913_),
    .Y(_04920_));
 sky130_fd_sc_hd__or3_1 _12338_ (.A(_04876_),
    .B(_04874_),
    .C(_04875_),
    .X(_04921_));
 sky130_fd_sc_hd__and2_1 _12339_ (.A(\wfg_stim_mem_top.cfg_gain_q[14] ),
    .B(_04533_),
    .X(_04922_));
 sky130_fd_sc_hd__a22o_1 _12340_ (.A1(_03212_),
    .A2(_04270_),
    .B1(_04346_),
    .B2(_03217_),
    .X(_04923_));
 sky130_fd_sc_hd__nand4_1 _12341_ (.A(_03532_),
    .B(_03531_),
    .C(_04520_),
    .D(_04522_),
    .Y(_04924_));
 sky130_fd_sc_hd__a21bo_1 _12342_ (.A1(_04922_),
    .A2(_04923_),
    .B1_N(_04924_),
    .X(_04925_));
 sky130_fd_sc_hd__o21ai_1 _12343_ (.A1(_04876_),
    .A2(_04875_),
    .B1(_04874_),
    .Y(_04926_));
 sky130_fd_sc_hd__nand3_1 _12344_ (.A(_04921_),
    .B(_04925_),
    .C(_04926_),
    .Y(_04927_));
 sky130_fd_sc_hd__a21o_1 _12345_ (.A1(_04921_),
    .A2(_04926_),
    .B1(_04925_),
    .X(_04928_));
 sky130_fd_sc_hd__nand2_1 _12346_ (.A(_02892_),
    .B(_04555_),
    .Y(_04929_));
 sky130_fd_sc_hd__a22oi_1 _12347_ (.A1(_03873_),
    .A2(_04447_),
    .B1(_04444_),
    .B2(_03872_),
    .Y(_04930_));
 sky130_fd_sc_hd__and4_1 _12348_ (.A(_03636_),
    .B(_03637_),
    .C(_04447_),
    .D(_04444_),
    .X(_04931_));
 sky130_fd_sc_hd__nor2_1 _12349_ (.A(_04930_),
    .B(_04931_),
    .Y(_04932_));
 sky130_fd_sc_hd__xnor2_2 _12350_ (.A(_04929_),
    .B(_04932_),
    .Y(_04933_));
 sky130_fd_sc_hd__nand3_1 _12351_ (.A(_04927_),
    .B(_04928_),
    .C(_04933_),
    .Y(_04934_));
 sky130_fd_sc_hd__and2_1 _12352_ (.A(_04927_),
    .B(_04934_),
    .X(_04935_));
 sky130_fd_sc_hd__a21o_1 _12353_ (.A1(_04879_),
    .A2(_04880_),
    .B1(_04885_),
    .X(_04936_));
 sky130_fd_sc_hd__nand4_1 _12354_ (.A(_03144_),
    .B(_03830_),
    .C(_04512_),
    .D(_04517_),
    .Y(_04937_));
 sky130_fd_sc_hd__a22o_1 _12355_ (.A1(_02940_),
    .A2(net28),
    .B1(_04517_),
    .B2(_02943_),
    .X(_04938_));
 sky130_fd_sc_hd__nand4_1 _12356_ (.A(_03798_),
    .B(_04524_),
    .C(_04937_),
    .D(_04938_),
    .Y(_04939_));
 sky130_fd_sc_hd__nand2_1 _12357_ (.A(_04937_),
    .B(_04939_),
    .Y(_04940_));
 sky130_fd_sc_hd__o21ai_1 _12358_ (.A1(_04858_),
    .A2(_04860_),
    .B1(_04859_),
    .Y(_04941_));
 sky130_fd_sc_hd__and2_1 _12359_ (.A(\wfg_stim_mem_top.cfg_gain_q[20] ),
    .B(net26),
    .X(_04942_));
 sky130_fd_sc_hd__a22o_1 _12360_ (.A1(_02954_),
    .A2(net23),
    .B1(net12),
    .B2(_03774_),
    .X(_04943_));
 sky130_fd_sc_hd__clkbuf_4 _12361_ (.A(net12),
    .X(_04944_));
 sky130_fd_sc_hd__nand4_1 _12362_ (.A(_03774_),
    .B(_03773_),
    .C(_04686_),
    .D(_04944_),
    .Y(_04945_));
 sky130_fd_sc_hd__a21bo_1 _12363_ (.A1(_04942_),
    .A2(_04943_),
    .B1_N(_04945_),
    .X(_04946_));
 sky130_fd_sc_hd__a21o_1 _12364_ (.A1(_04861_),
    .A2(_04941_),
    .B1(_04946_),
    .X(_04947_));
 sky130_fd_sc_hd__nand3_1 _12365_ (.A(_04861_),
    .B(_04946_),
    .C(_04941_),
    .Y(_04948_));
 sky130_fd_sc_hd__a21bo_1 _12366_ (.A1(_04940_),
    .A2(_04947_),
    .B1_N(_04948_),
    .X(_04949_));
 sky130_fd_sc_hd__a21oi_1 _12367_ (.A1(_04886_),
    .A2(_04936_),
    .B1(_04949_),
    .Y(_04950_));
 sky130_fd_sc_hd__and3_1 _12368_ (.A(_04886_),
    .B(_04949_),
    .C(_04936_),
    .X(_04951_));
 sky130_fd_sc_hd__o21ba_1 _12369_ (.A1(_04935_),
    .A2(_04950_),
    .B1_N(_04951_),
    .X(_04952_));
 sky130_fd_sc_hd__a21oi_1 _12370_ (.A1(_03954_),
    .A2(_04555_),
    .B1(_04900_),
    .Y(_04953_));
 sky130_fd_sc_hd__a31o_1 _12371_ (.A1(_03945_),
    .A2(_04555_),
    .A3(_04932_),
    .B1(_04931_),
    .X(_04954_));
 sky130_fd_sc_hd__nand2_1 _12372_ (.A(_03948_),
    .B(_03685_),
    .Y(_04955_));
 sky130_fd_sc_hd__xnor2_1 _12373_ (.A(_04954_),
    .B(_04955_),
    .Y(_04956_));
 sky130_fd_sc_hd__and3_1 _12374_ (.A(_03947_),
    .B(_04286_),
    .C(_04956_),
    .X(_04957_));
 sky130_fd_sc_hd__a31o_1 _12375_ (.A1(_03943_),
    .A2(_03685_),
    .A3(_04954_),
    .B1(_04957_),
    .X(_04958_));
 sky130_fd_sc_hd__nor2_1 _12376_ (.A(_04901_),
    .B(_04953_),
    .Y(_04959_));
 sky130_fd_sc_hd__xnor2_1 _12377_ (.A(_04952_),
    .B(_04959_),
    .Y(_04960_));
 sky130_fd_sc_hd__nand2_1 _12378_ (.A(_04958_),
    .B(_04960_),
    .Y(_04961_));
 sky130_fd_sc_hd__o31a_1 _12379_ (.A1(_04901_),
    .A2(_04952_),
    .A3(_04953_),
    .B1(_04961_),
    .X(_04962_));
 sky130_fd_sc_hd__or3_1 _12380_ (.A(_04896_),
    .B(_04897_),
    .C(_04907_),
    .X(_04963_));
 sky130_fd_sc_hd__o21ai_1 _12381_ (.A1(_04896_),
    .A2(_04897_),
    .B1(_04907_),
    .Y(_04964_));
 sky130_fd_sc_hd__a21oi_1 _12382_ (.A1(_04844_),
    .A2(_04845_),
    .B1(_04846_),
    .Y(_04965_));
 sky130_fd_sc_hd__or4bb_1 _12383_ (.A(_04853_),
    .B(_04965_),
    .C_N(_04851_),
    .D_N(_04852_),
    .X(_04966_));
 sky130_fd_sc_hd__buf_4 _12384_ (.A(net1),
    .X(_04967_));
 sky130_fd_sc_hd__a22oi_2 _12385_ (.A1(_03596_),
    .A2(_03771_),
    .B1(_04967_),
    .B2(_03759_),
    .Y(_04968_));
 sky130_fd_sc_hd__nor2_1 _12386_ (.A(_04846_),
    .B(_04968_),
    .Y(_04969_));
 sky130_fd_sc_hd__nand3_1 _12387_ (.A(_04942_),
    .B(_04943_),
    .C(_04945_),
    .Y(_04970_));
 sky130_fd_sc_hd__a21o_1 _12388_ (.A1(_04943_),
    .A2(_04945_),
    .B1(_04942_),
    .X(_04971_));
 sky130_fd_sc_hd__and3_2 _12389_ (.A(_04969_),
    .B(_04970_),
    .C(_04971_),
    .X(_04972_));
 sky130_fd_sc_hd__a2bb2o_1 _12390_ (.A1_N(_04853_),
    .A2_N(_04965_),
    .B1(_04851_),
    .B2(_04852_),
    .X(_04973_));
 sky130_fd_sc_hd__and3_2 _12391_ (.A(_04966_),
    .B(_04972_),
    .C(_04973_),
    .X(_04974_));
 sky130_fd_sc_hd__nand3_1 _12392_ (.A(_04966_),
    .B(_04972_),
    .C(_04973_),
    .Y(_04975_));
 sky130_fd_sc_hd__a21o_1 _12393_ (.A1(_04966_),
    .A2(_04973_),
    .B1(_04972_),
    .X(_04976_));
 sky130_fd_sc_hd__nand3_1 _12394_ (.A(_04940_),
    .B(_04948_),
    .C(_04947_),
    .Y(_04977_));
 sky130_fd_sc_hd__a21o_1 _12395_ (.A1(_04948_),
    .A2(_04947_),
    .B1(_04940_),
    .X(_04978_));
 sky130_fd_sc_hd__and4_2 _12396_ (.A(_04975_),
    .B(_04976_),
    .C(_04977_),
    .D(_04978_),
    .X(_04979_));
 sky130_fd_sc_hd__a22o_1 _12397_ (.A1(_04856_),
    .A2(_04857_),
    .B1(_04867_),
    .B2(_04868_),
    .X(_04980_));
 sky130_fd_sc_hd__o211ai_4 _12398_ (.A1(_04974_),
    .A2(_04979_),
    .B1(_04980_),
    .C1(_04869_),
    .Y(_04981_));
 sky130_fd_sc_hd__o211a_1 _12399_ (.A1(_04974_),
    .A2(_04979_),
    .B1(_04980_),
    .C1(_04869_),
    .X(_04982_));
 sky130_fd_sc_hd__a211oi_2 _12400_ (.A1(_04869_),
    .A2(_04980_),
    .B1(_04979_),
    .C1(_04974_),
    .Y(_04983_));
 sky130_fd_sc_hd__nor3_1 _12401_ (.A(_04935_),
    .B(_04951_),
    .C(_04950_),
    .Y(_04984_));
 sky130_fd_sc_hd__o21a_1 _12402_ (.A1(_04951_),
    .A2(_04950_),
    .B1(_04935_),
    .X(_04985_));
 sky130_fd_sc_hd__or4_4 _12403_ (.A(_04982_),
    .B(_04983_),
    .C(_04984_),
    .D(_04985_),
    .X(_04986_));
 sky130_fd_sc_hd__o22a_1 _12404_ (.A1(_04871_),
    .A2(_04872_),
    .B1(_04892_),
    .B2(_04893_),
    .X(_04987_));
 sky130_fd_sc_hd__a211oi_4 _12405_ (.A1(_04981_),
    .A2(_04986_),
    .B1(_04987_),
    .C1(_04894_),
    .Y(_04988_));
 sky130_fd_sc_hd__o211a_1 _12406_ (.A1(_04894_),
    .A2(_04987_),
    .B1(_04986_),
    .C1(_04981_),
    .X(_04989_));
 sky130_fd_sc_hd__xnor2_1 _12407_ (.A(_04958_),
    .B(_04960_),
    .Y(_04990_));
 sky130_fd_sc_hd__nor3_1 _12408_ (.A(_04988_),
    .B(_04989_),
    .C(_04990_),
    .Y(_04991_));
 sky130_fd_sc_hd__a211oi_2 _12409_ (.A1(_04963_),
    .A2(_04964_),
    .B1(_04991_),
    .C1(_04988_),
    .Y(_04992_));
 sky130_fd_sc_hd__o211a_1 _12410_ (.A1(_04988_),
    .A2(_04991_),
    .B1(_04964_),
    .C1(_04963_),
    .X(_04993_));
 sky130_fd_sc_hd__o21bai_1 _12411_ (.A1(_04962_),
    .A2(_04992_),
    .B1_N(_04993_),
    .Y(_04994_));
 sky130_fd_sc_hd__nor3b_2 _12412_ (.A(_04916_),
    .B(_04920_),
    .C_N(_04994_),
    .Y(_04995_));
 sky130_fd_sc_hd__o21ba_1 _12413_ (.A1(_04916_),
    .A2(_04920_),
    .B1_N(_04994_),
    .X(_04996_));
 sky130_fd_sc_hd__nor2_4 _12414_ (.A(_04995_),
    .B(_04996_),
    .Y(_04997_));
 sky130_fd_sc_hd__and4_1 _12415_ (.A(_04760_),
    .B(_04839_),
    .C(_04919_),
    .D(_04997_),
    .X(_04998_));
 sky130_fd_sc_hd__and2_1 _12416_ (.A(\wfg_stim_mem_top.cfg_gain_q[20] ),
    .B(net23),
    .X(_04999_));
 sky130_fd_sc_hd__a22o_1 _12417_ (.A1(_03773_),
    .A2(net12),
    .B1(net1),
    .B2(_03774_),
    .X(_05000_));
 sky130_fd_sc_hd__nand4_1 _12418_ (.A(_02963_),
    .B(_02965_),
    .C(_04944_),
    .D(net1),
    .Y(_05001_));
 sky130_fd_sc_hd__nand3_1 _12419_ (.A(_04999_),
    .B(_05000_),
    .C(_05001_),
    .Y(_05002_));
 sky130_fd_sc_hd__a21o_1 _12420_ (.A1(_05000_),
    .A2(_05001_),
    .B1(_04999_),
    .X(_05003_));
 sky130_fd_sc_hd__nand4_2 _12421_ (.A(_03069_),
    .B(_04448_),
    .C(_05002_),
    .D(_05003_),
    .Y(_05004_));
 sky130_fd_sc_hd__a21oi_2 _12422_ (.A1(_04970_),
    .A2(_04971_),
    .B1(_04969_),
    .Y(_05005_));
 sky130_fd_sc_hd__or3_4 _12423_ (.A(_04972_),
    .B(_05004_),
    .C(_05005_),
    .X(_05006_));
 sky130_fd_sc_hd__o21ai_2 _12424_ (.A1(_04972_),
    .A2(_05005_),
    .B1(_05004_),
    .Y(_05007_));
 sky130_fd_sc_hd__and4_1 _12425_ (.A(_03143_),
    .B(_02937_),
    .C(net27),
    .D(net26),
    .X(_05008_));
 sky130_fd_sc_hd__nand2_1 _12426_ (.A(\wfg_stim_mem_top.cfg_gain_q[17] ),
    .B(net28),
    .Y(_05009_));
 sky130_fd_sc_hd__a22oi_1 _12427_ (.A1(_02937_),
    .A2(_04517_),
    .B1(_04681_),
    .B2(_02943_),
    .Y(_05010_));
 sky130_fd_sc_hd__or3_1 _12428_ (.A(_05008_),
    .B(_05009_),
    .C(_05010_),
    .X(_05011_));
 sky130_fd_sc_hd__or2b_1 _12429_ (.A(_05008_),
    .B_N(_05011_),
    .X(_05012_));
 sky130_fd_sc_hd__a21bo_1 _12430_ (.A1(_04999_),
    .A2(_05000_),
    .B1_N(_05001_),
    .X(_05013_));
 sky130_fd_sc_hd__a22o_1 _12431_ (.A1(_03798_),
    .A2(_04524_),
    .B1(_04937_),
    .B2(_04938_),
    .X(_05014_));
 sky130_fd_sc_hd__nand3_1 _12432_ (.A(_04939_),
    .B(_05013_),
    .C(_05014_),
    .Y(_05015_));
 sky130_fd_sc_hd__a21o_1 _12433_ (.A1(_04939_),
    .A2(_05014_),
    .B1(_05013_),
    .X(_05016_));
 sky130_fd_sc_hd__nand3_1 _12434_ (.A(_05012_),
    .B(_05015_),
    .C(_05016_),
    .Y(_05017_));
 sky130_fd_sc_hd__a21o_1 _12435_ (.A1(_05015_),
    .A2(_05016_),
    .B1(_05012_),
    .X(_05018_));
 sky130_fd_sc_hd__nand4_4 _12436_ (.A(_05006_),
    .B(_05007_),
    .C(_05017_),
    .D(_05018_),
    .Y(_05019_));
 sky130_fd_sc_hd__a22oi_4 _12437_ (.A1(_04975_),
    .A2(_04976_),
    .B1(_04977_),
    .B2(_04978_),
    .Y(_05020_));
 sky130_fd_sc_hd__a211oi_4 _12438_ (.A1(_05006_),
    .A2(_05019_),
    .B1(_05020_),
    .C1(_04979_),
    .Y(_05021_));
 sky130_fd_sc_hd__o211a_1 _12439_ (.A1(_04979_),
    .A2(_05020_),
    .B1(_05019_),
    .C1(_05006_),
    .X(_05022_));
 sky130_fd_sc_hd__nand3_1 _12440_ (.A(_04924_),
    .B(_04922_),
    .C(_04923_),
    .Y(_05023_));
 sky130_fd_sc_hd__nand2_1 _12441_ (.A(_03529_),
    .B(_04520_),
    .Y(_05024_));
 sky130_fd_sc_hd__a22oi_2 _12442_ (.A1(_03531_),
    .A2(_04522_),
    .B1(_04524_),
    .B2(_03532_),
    .Y(_05025_));
 sky130_fd_sc_hd__and4_2 _12443_ (.A(_03217_),
    .B(_03212_),
    .C(_04346_),
    .D(_04426_),
    .X(_05026_));
 sky130_fd_sc_hd__o21bai_2 _12444_ (.A1(_05024_),
    .A2(_05025_),
    .B1_N(_05026_),
    .Y(_05027_));
 sky130_fd_sc_hd__a22o_1 _12445_ (.A1(_02926_),
    .A2(_04533_),
    .B1(_04924_),
    .B2(_04923_),
    .X(_05028_));
 sky130_fd_sc_hd__nand3_1 _12446_ (.A(_05023_),
    .B(_05027_),
    .C(_05028_),
    .Y(_05029_));
 sky130_fd_sc_hd__a21o_1 _12447_ (.A1(_05023_),
    .A2(_05028_),
    .B1(_05027_),
    .X(_05030_));
 sky130_fd_sc_hd__nand2_1 _12448_ (.A(_02892_),
    .B(_04286_),
    .Y(_05031_));
 sky130_fd_sc_hd__a22oi_1 _12449_ (.A1(_02896_),
    .A2(_04444_),
    .B1(_04445_),
    .B2(_02894_),
    .Y(_05032_));
 sky130_fd_sc_hd__and4_1 _12450_ (.A(_03633_),
    .B(_02899_),
    .C(_04444_),
    .D(_04445_),
    .X(_05033_));
 sky130_fd_sc_hd__nor2_1 _12451_ (.A(_05032_),
    .B(_05033_),
    .Y(_05034_));
 sky130_fd_sc_hd__xnor2_2 _12452_ (.A(_05031_),
    .B(_05034_),
    .Y(_05035_));
 sky130_fd_sc_hd__nand3_1 _12453_ (.A(_05029_),
    .B(_05030_),
    .C(_05035_),
    .Y(_05036_));
 sky130_fd_sc_hd__nand2_1 _12454_ (.A(_05029_),
    .B(_05036_),
    .Y(_05037_));
 sky130_fd_sc_hd__a21bo_1 _12455_ (.A1(_05012_),
    .A2(_05016_),
    .B1_N(_05015_),
    .X(_05038_));
 sky130_fd_sc_hd__a21o_1 _12456_ (.A1(_04927_),
    .A2(_04928_),
    .B1(_04933_),
    .X(_05039_));
 sky130_fd_sc_hd__nand3_1 _12457_ (.A(_04934_),
    .B(_05038_),
    .C(_05039_),
    .Y(_05040_));
 sky130_fd_sc_hd__a21o_1 _12458_ (.A1(_04934_),
    .A2(_05039_),
    .B1(_05038_),
    .X(_05041_));
 sky130_fd_sc_hd__and3_1 _12459_ (.A(_05037_),
    .B(_05040_),
    .C(_05041_),
    .X(_05042_));
 sky130_fd_sc_hd__a21oi_2 _12460_ (.A1(_05040_),
    .A2(_05041_),
    .B1(_05037_),
    .Y(_05043_));
 sky130_fd_sc_hd__nor4_4 _12461_ (.A(_05021_),
    .B(_05022_),
    .C(_05042_),
    .D(_05043_),
    .Y(_05044_));
 sky130_fd_sc_hd__o22ai_2 _12462_ (.A1(_04982_),
    .A2(_04983_),
    .B1(_04984_),
    .B2(_04985_),
    .Y(_05045_));
 sky130_fd_sc_hd__o211a_2 _12463_ (.A1(_05021_),
    .A2(_05044_),
    .B1(_05045_),
    .C1(_04986_),
    .X(_05046_));
 sky130_fd_sc_hd__a211oi_2 _12464_ (.A1(_04986_),
    .A2(_05045_),
    .B1(_05044_),
    .C1(_05021_),
    .Y(_05047_));
 sky130_fd_sc_hd__a31o_1 _12465_ (.A1(_03491_),
    .A2(_04286_),
    .A3(_05034_),
    .B1(_05033_),
    .X(_05048_));
 sky130_fd_sc_hd__nand2_1 _12466_ (.A(_02887_),
    .B(_03675_),
    .Y(_05049_));
 sky130_fd_sc_hd__xnor2_1 _12467_ (.A(_05048_),
    .B(_05049_),
    .Y(_05050_));
 sky130_fd_sc_hd__and3_1 _12468_ (.A(_03947_),
    .B(_04551_),
    .C(_05050_),
    .X(_05051_));
 sky130_fd_sc_hd__a31o_1 _12469_ (.A1(_03944_),
    .A2(_03675_),
    .A3(_05048_),
    .B1(_05051_),
    .X(_05052_));
 sky130_fd_sc_hd__a21boi_2 _12470_ (.A1(_05037_),
    .A2(_05041_),
    .B1_N(_05040_),
    .Y(_05053_));
 sky130_fd_sc_hd__a21oi_1 _12471_ (.A1(_02908_),
    .A2(_04286_),
    .B1(_04956_),
    .Y(_05054_));
 sky130_fd_sc_hd__nor2_1 _12472_ (.A(_04957_),
    .B(_05054_),
    .Y(_05055_));
 sky130_fd_sc_hd__xnor2_1 _12473_ (.A(_05053_),
    .B(_05055_),
    .Y(_05056_));
 sky130_fd_sc_hd__xnor2_1 _12474_ (.A(_05052_),
    .B(_05056_),
    .Y(_05057_));
 sky130_fd_sc_hd__nor3_1 _12475_ (.A(_05046_),
    .B(_05047_),
    .C(_05057_),
    .Y(_05058_));
 sky130_fd_sc_hd__o21ai_1 _12476_ (.A1(_04988_),
    .A2(_04989_),
    .B1(_04990_),
    .Y(_05059_));
 sky130_fd_sc_hd__or3_1 _12477_ (.A(_04988_),
    .B(_04989_),
    .C(_04990_),
    .X(_05060_));
 sky130_fd_sc_hd__o211a_1 _12478_ (.A1(_05046_),
    .A2(_05058_),
    .B1(_05059_),
    .C1(_05060_),
    .X(_05061_));
 sky130_fd_sc_hd__inv_2 _12479_ (.A(_05061_),
    .Y(_05062_));
 sky130_fd_sc_hd__or3_1 _12480_ (.A(_04957_),
    .B(_05053_),
    .C(_05054_),
    .X(_05063_));
 sky130_fd_sc_hd__nand2_1 _12481_ (.A(_05052_),
    .B(_05056_),
    .Y(_05064_));
 sky130_fd_sc_hd__a211oi_2 _12482_ (.A1(_05060_),
    .A2(_05059_),
    .B1(_05058_),
    .C1(_05046_),
    .Y(_05065_));
 sky130_fd_sc_hd__a211o_1 _12483_ (.A1(_05063_),
    .A2(_05064_),
    .B1(_05061_),
    .C1(_05065_),
    .X(_05066_));
 sky130_fd_sc_hd__nor3_1 _12484_ (.A(_04993_),
    .B(_04962_),
    .C(_04992_),
    .Y(_05067_));
 sky130_fd_sc_hd__o21a_1 _12485_ (.A1(_04993_),
    .A2(_04992_),
    .B1(_04962_),
    .X(_05068_));
 sky130_fd_sc_hd__a211oi_1 _12486_ (.A1(_05062_),
    .A2(_05066_),
    .B1(_05067_),
    .C1(_05068_),
    .Y(_05069_));
 sky130_fd_sc_hd__o211ai_2 _12487_ (.A1(_05067_),
    .A2(_05068_),
    .B1(_05062_),
    .C1(_05066_),
    .Y(_05070_));
 sky130_fd_sc_hd__nand2b_2 _12488_ (.A_N(_05069_),
    .B(_05070_),
    .Y(_05071_));
 sky130_fd_sc_hd__a211oi_2 _12489_ (.A1(_05063_),
    .A2(_05064_),
    .B1(_05061_),
    .C1(_05065_),
    .Y(_05072_));
 sky130_fd_sc_hd__o211a_1 _12490_ (.A1(_05061_),
    .A2(_05065_),
    .B1(_05063_),
    .C1(_05064_),
    .X(_05073_));
 sky130_fd_sc_hd__or3_1 _12491_ (.A(_05026_),
    .B(_05024_),
    .C(_05025_),
    .X(_05074_));
 sky130_fd_sc_hd__and2_1 _12492_ (.A(_03529_),
    .B(_04522_),
    .X(_05075_));
 sky130_fd_sc_hd__a22o_1 _12493_ (.A1(_03210_),
    .A2(_04524_),
    .B1(_04512_),
    .B2(_03208_),
    .X(_05076_));
 sky130_fd_sc_hd__clkbuf_4 _12494_ (.A(_04512_),
    .X(_05077_));
 sky130_fd_sc_hd__nand4_1 _12495_ (.A(_03218_),
    .B(_03213_),
    .C(_04524_),
    .D(_05077_),
    .Y(_05078_));
 sky130_fd_sc_hd__a21bo_1 _12496_ (.A1(_05075_),
    .A2(_05076_),
    .B1_N(_05078_),
    .X(_05079_));
 sky130_fd_sc_hd__o21ai_1 _12497_ (.A1(_05026_),
    .A2(_05025_),
    .B1(_05024_),
    .Y(_05080_));
 sky130_fd_sc_hd__nand3_1 _12498_ (.A(_05074_),
    .B(_05079_),
    .C(_05080_),
    .Y(_05081_));
 sky130_fd_sc_hd__a21o_1 _12499_ (.A1(_05074_),
    .A2(_05080_),
    .B1(_05079_),
    .X(_05082_));
 sky130_fd_sc_hd__nand2_1 _12500_ (.A(_03490_),
    .B(_04551_),
    .Y(_05083_));
 sky130_fd_sc_hd__buf_4 _12501_ (.A(_04533_),
    .X(_05084_));
 sky130_fd_sc_hd__a22oi_1 _12502_ (.A1(_03873_),
    .A2(_04445_),
    .B1(_05084_),
    .B2(_03872_),
    .Y(_05085_));
 sky130_fd_sc_hd__and4_1 _12503_ (.A(_02894_),
    .B(_02896_),
    .C(_04445_),
    .D(_04533_),
    .X(_05086_));
 sky130_fd_sc_hd__nor2_1 _12504_ (.A(_05085_),
    .B(_05086_),
    .Y(_05087_));
 sky130_fd_sc_hd__xnor2_1 _12505_ (.A(_05083_),
    .B(_05087_),
    .Y(_05088_));
 sky130_fd_sc_hd__nand3_1 _12506_ (.A(_05081_),
    .B(_05082_),
    .C(_05088_),
    .Y(_05089_));
 sky130_fd_sc_hd__and2_1 _12507_ (.A(_05081_),
    .B(_05089_),
    .X(_05090_));
 sky130_fd_sc_hd__a21o_1 _12508_ (.A1(_05029_),
    .A2(_05030_),
    .B1(_05035_),
    .X(_05091_));
 sky130_fd_sc_hd__buf_2 _12509_ (.A(_04681_),
    .X(_05092_));
 sky130_fd_sc_hd__clkbuf_4 _12510_ (.A(_04686_),
    .X(_05093_));
 sky130_fd_sc_hd__a22o_1 _12511_ (.A1(_02938_),
    .A2(_05092_),
    .B1(_05093_),
    .B2(_03144_),
    .X(_05094_));
 sky130_fd_sc_hd__and4_1 _12512_ (.A(_03144_),
    .B(_02938_),
    .C(_04681_),
    .D(_04686_),
    .X(_05095_));
 sky130_fd_sc_hd__a31o_2 _12513_ (.A1(_02935_),
    .A2(_04643_),
    .A3(_05094_),
    .B1(_05095_),
    .X(_05096_));
 sky130_fd_sc_hd__o21ai_1 _12514_ (.A1(_05008_),
    .A2(_05010_),
    .B1(_05009_),
    .Y(_05097_));
 sky130_fd_sc_hd__and4_1 _12515_ (.A(_02955_),
    .B(_02948_),
    .C(_04944_),
    .D(net1),
    .X(_05098_));
 sky130_fd_sc_hd__a21o_1 _12516_ (.A1(_05011_),
    .A2(_05097_),
    .B1(_05098_),
    .X(_05099_));
 sky130_fd_sc_hd__nand3_1 _12517_ (.A(_05011_),
    .B(_05098_),
    .C(_05097_),
    .Y(_05100_));
 sky130_fd_sc_hd__a21bo_1 _12518_ (.A1(_05096_),
    .A2(_05099_),
    .B1_N(_05100_),
    .X(_05101_));
 sky130_fd_sc_hd__a21oi_1 _12519_ (.A1(_05036_),
    .A2(_05091_),
    .B1(_05101_),
    .Y(_05102_));
 sky130_fd_sc_hd__and3_1 _12520_ (.A(_05036_),
    .B(_05101_),
    .C(_05091_),
    .X(_05103_));
 sky130_fd_sc_hd__o21ba_1 _12521_ (.A1(_05090_),
    .A2(_05102_),
    .B1_N(_05103_),
    .X(_05104_));
 sky130_fd_sc_hd__a21oi_1 _12522_ (.A1(_03954_),
    .A2(_04551_),
    .B1(_05050_),
    .Y(_05105_));
 sky130_fd_sc_hd__or3_1 _12523_ (.A(_05051_),
    .B(_05104_),
    .C(_05105_),
    .X(_05106_));
 sky130_fd_sc_hd__a31o_1 _12524_ (.A1(_03945_),
    .A2(_04551_),
    .A3(_05087_),
    .B1(_05086_),
    .X(_05107_));
 sky130_fd_sc_hd__nand2_1 _12525_ (.A(_03948_),
    .B(_04555_),
    .Y(_05108_));
 sky130_fd_sc_hd__xnor2_1 _12526_ (.A(_05107_),
    .B(_05108_),
    .Y(_05109_));
 sky130_fd_sc_hd__and3_1 _12527_ (.A(_03947_),
    .B(_04448_),
    .C(_05109_),
    .X(_05110_));
 sky130_fd_sc_hd__a31o_1 _12528_ (.A1(_03943_),
    .A2(_04555_),
    .A3(_05107_),
    .B1(_05110_),
    .X(_05111_));
 sky130_fd_sc_hd__nor2_1 _12529_ (.A(_05051_),
    .B(_05105_),
    .Y(_05112_));
 sky130_fd_sc_hd__xnor2_1 _12530_ (.A(_05104_),
    .B(_05112_),
    .Y(_05113_));
 sky130_fd_sc_hd__nand2_1 _12531_ (.A(_05111_),
    .B(_05113_),
    .Y(_05114_));
 sky130_fd_sc_hd__nand2_1 _12532_ (.A(_05106_),
    .B(_05114_),
    .Y(_05115_));
 sky130_fd_sc_hd__or3_1 _12533_ (.A(_05046_),
    .B(_05047_),
    .C(_05057_),
    .X(_05116_));
 sky130_fd_sc_hd__o21ai_1 _12534_ (.A1(_05046_),
    .A2(_05047_),
    .B1(_05057_),
    .Y(_05117_));
 sky130_fd_sc_hd__clkbuf_4 _12535_ (.A(_04944_),
    .X(_05118_));
 sky130_fd_sc_hd__a22oi_1 _12536_ (.A1(_02949_),
    .A2(_05118_),
    .B1(_04967_),
    .B2(_02955_),
    .Y(_05119_));
 sky130_fd_sc_hd__and4bb_1 _12537_ (.A_N(_05119_),
    .B_N(_05098_),
    .C(_03069_),
    .D(_04535_),
    .X(_05120_));
 sky130_fd_sc_hd__a22o_1 _12538_ (.A1(_03069_),
    .A2(_04448_),
    .B1(_05002_),
    .B2(_05003_),
    .X(_05121_));
 sky130_fd_sc_hd__and3_2 _12539_ (.A(_05004_),
    .B(_05120_),
    .C(_05121_),
    .X(_05122_));
 sky130_fd_sc_hd__a21oi_2 _12540_ (.A1(_05004_),
    .A2(_05121_),
    .B1(_05120_),
    .Y(_05123_));
 sky130_fd_sc_hd__and3_1 _12541_ (.A(_05096_),
    .B(_05100_),
    .C(_05099_),
    .X(_05124_));
 sky130_fd_sc_hd__a21oi_2 _12542_ (.A1(_05100_),
    .A2(_05099_),
    .B1(_05096_),
    .Y(_05125_));
 sky130_fd_sc_hd__nor4_4 _12543_ (.A(_05122_),
    .B(_05123_),
    .C(_05124_),
    .D(_05125_),
    .Y(_05126_));
 sky130_fd_sc_hd__a22o_2 _12544_ (.A1(_05006_),
    .A2(_05007_),
    .B1(_05017_),
    .B2(_05018_),
    .X(_05127_));
 sky130_fd_sc_hd__o211ai_4 _12545_ (.A1(_05122_),
    .A2(_05126_),
    .B1(_05127_),
    .C1(_05019_),
    .Y(_05128_));
 sky130_fd_sc_hd__o211a_1 _12546_ (.A1(_05122_),
    .A2(_05126_),
    .B1(_05127_),
    .C1(_05019_),
    .X(_05129_));
 sky130_fd_sc_hd__a211oi_2 _12547_ (.A1(_05019_),
    .A2(_05127_),
    .B1(_05126_),
    .C1(_05122_),
    .Y(_05130_));
 sky130_fd_sc_hd__nor3_2 _12548_ (.A(_05090_),
    .B(_05103_),
    .C(_05102_),
    .Y(_05131_));
 sky130_fd_sc_hd__o21a_1 _12549_ (.A1(_05103_),
    .A2(_05102_),
    .B1(_05090_),
    .X(_05132_));
 sky130_fd_sc_hd__or4_4 _12550_ (.A(_05129_),
    .B(_05130_),
    .C(_05131_),
    .D(_05132_),
    .X(_05133_));
 sky130_fd_sc_hd__o22a_2 _12551_ (.A1(_05021_),
    .A2(_05022_),
    .B1(_05042_),
    .B2(_05043_),
    .X(_05134_));
 sky130_fd_sc_hd__a211oi_4 _12552_ (.A1(_05128_),
    .A2(_05133_),
    .B1(_05134_),
    .C1(_05044_),
    .Y(_05135_));
 sky130_fd_sc_hd__o211a_1 _12553_ (.A1(_05044_),
    .A2(_05134_),
    .B1(_05133_),
    .C1(_05128_),
    .X(_05136_));
 sky130_fd_sc_hd__xnor2_1 _12554_ (.A(_05111_),
    .B(_05113_),
    .Y(_05137_));
 sky130_fd_sc_hd__nor3_1 _12555_ (.A(_05135_),
    .B(_05136_),
    .C(_05137_),
    .Y(_05138_));
 sky130_fd_sc_hd__a211o_1 _12556_ (.A1(_05116_),
    .A2(_05117_),
    .B1(_05138_),
    .C1(_05135_),
    .X(_05139_));
 sky130_fd_sc_hd__o211a_1 _12557_ (.A1(_05135_),
    .A2(_05138_),
    .B1(_05117_),
    .C1(_05116_),
    .X(_05140_));
 sky130_fd_sc_hd__a21oi_1 _12558_ (.A1(_05115_),
    .A2(_05139_),
    .B1(_05140_),
    .Y(_05141_));
 sky130_fd_sc_hd__nor3_2 _12559_ (.A(_05072_),
    .B(_05073_),
    .C(_05141_),
    .Y(_05142_));
 sky130_fd_sc_hd__o21a_1 _12560_ (.A1(_05072_),
    .A2(_05073_),
    .B1(_05141_),
    .X(_05143_));
 sky130_fd_sc_hd__or2_1 _12561_ (.A(_05142_),
    .B(_05143_),
    .X(_05144_));
 sky130_fd_sc_hd__buf_2 _12562_ (.A(_04967_),
    .X(_05145_));
 sky130_fd_sc_hd__and4_1 _12563_ (.A(_02949_),
    .B(_03069_),
    .C(_04616_),
    .D(_05145_),
    .X(_05146_));
 sky130_fd_sc_hd__clkbuf_4 _12564_ (.A(_05145_),
    .X(_05147_));
 sky130_fd_sc_hd__a22oi_1 _12565_ (.A1(_03434_),
    .A2(_04616_),
    .B1(_05147_),
    .B2(_03100_),
    .Y(_05148_));
 sky130_fd_sc_hd__or2_1 _12566_ (.A(_05146_),
    .B(_05148_),
    .X(_05149_));
 sky130_fd_sc_hd__nand2_1 _12567_ (.A(_03239_),
    .B(_05092_),
    .Y(_05150_));
 sky130_fd_sc_hd__and4_1 _12568_ (.A(_03799_),
    .B(_03830_),
    .C(_04686_),
    .D(_04944_),
    .X(_05151_));
 sky130_fd_sc_hd__a22o_1 _12569_ (.A1(_03830_),
    .A2(_04686_),
    .B1(_04944_),
    .B2(_03144_),
    .X(_05152_));
 sky130_fd_sc_hd__and2b_1 _12570_ (.A_N(_05151_),
    .B(_05152_),
    .X(_05153_));
 sky130_fd_sc_hd__xnor2_1 _12571_ (.A(_05150_),
    .B(_05153_),
    .Y(_05154_));
 sky130_fd_sc_hd__a22o_1 _12572_ (.A1(_03830_),
    .A2(_04944_),
    .B1(_04967_),
    .B2(_03799_),
    .X(_05155_));
 sky130_fd_sc_hd__and4_1 _12573_ (.A(_03799_),
    .B(_03830_),
    .C(_04944_),
    .D(_04967_),
    .X(_05156_));
 sky130_fd_sc_hd__a31o_1 _12574_ (.A1(_03239_),
    .A2(_05093_),
    .A3(_05155_),
    .B1(_05156_),
    .X(_05157_));
 sky130_fd_sc_hd__xor2_1 _12575_ (.A(_05154_),
    .B(_05157_),
    .X(_05158_));
 sky130_fd_sc_hd__or2b_1 _12576_ (.A(_05149_),
    .B_N(_05158_),
    .X(_05159_));
 sky130_fd_sc_hd__o2bb2a_1 _12577_ (.A1_N(_03069_),
    .A2_N(_04535_),
    .B1(_05119_),
    .B2(_05098_),
    .X(_05160_));
 sky130_fd_sc_hd__nor2_2 _12578_ (.A(_05120_),
    .B(_05160_),
    .Y(_05161_));
 sky130_fd_sc_hd__xnor2_1 _12579_ (.A(_05146_),
    .B(_05161_),
    .Y(_05162_));
 sky130_fd_sc_hd__clkbuf_4 _12580_ (.A(_04643_),
    .X(_05163_));
 sky130_fd_sc_hd__nand2_1 _12581_ (.A(_03239_),
    .B(_05163_),
    .Y(_05164_));
 sky130_fd_sc_hd__and2b_1 _12582_ (.A_N(_05095_),
    .B(_05094_),
    .X(_05165_));
 sky130_fd_sc_hd__xnor2_1 _12583_ (.A(_05164_),
    .B(_05165_),
    .Y(_05166_));
 sky130_fd_sc_hd__clkbuf_4 _12584_ (.A(_05092_),
    .X(_05167_));
 sky130_fd_sc_hd__a31o_1 _12585_ (.A1(_03142_),
    .A2(_05167_),
    .A3(_05152_),
    .B1(_05151_),
    .X(_05168_));
 sky130_fd_sc_hd__xor2_1 _12586_ (.A(_05166_),
    .B(_05168_),
    .X(_05169_));
 sky130_fd_sc_hd__xnor2_1 _12587_ (.A(_05162_),
    .B(_05169_),
    .Y(_05170_));
 sky130_fd_sc_hd__and2b_1 _12588_ (.A_N(_05159_),
    .B(_05170_),
    .X(_05171_));
 sky130_fd_sc_hd__xnor2_1 _12589_ (.A(_05159_),
    .B(_05170_),
    .Y(_05172_));
 sky130_fd_sc_hd__and4_2 _12590_ (.A(_02920_),
    .B(_03212_),
    .C(_04512_),
    .D(_04517_),
    .X(_05173_));
 sky130_fd_sc_hd__nand2_1 _12591_ (.A(_03529_),
    .B(_04524_),
    .Y(_05174_));
 sky130_fd_sc_hd__a22oi_2 _12592_ (.A1(_03210_),
    .A2(_04512_),
    .B1(_04643_),
    .B2(_03208_),
    .Y(_05175_));
 sky130_fd_sc_hd__or3_1 _12593_ (.A(_05173_),
    .B(_05174_),
    .C(_05175_),
    .X(_05176_));
 sky130_fd_sc_hd__a22o_1 _12594_ (.A1(_03531_),
    .A2(_04643_),
    .B1(_05092_),
    .B2(_03532_),
    .X(_05177_));
 sky130_fd_sc_hd__and4_1 _12595_ (.A(_03532_),
    .B(_02922_),
    .C(_04643_),
    .D(_04681_),
    .X(_05178_));
 sky130_fd_sc_hd__a31o_1 _12596_ (.A1(_02927_),
    .A2(_05077_),
    .A3(_05177_),
    .B1(_05178_),
    .X(_05179_));
 sky130_fd_sc_hd__o21ai_1 _12597_ (.A1(_05173_),
    .A2(_05175_),
    .B1(_05174_),
    .Y(_05180_));
 sky130_fd_sc_hd__nand3_1 _12598_ (.A(_05176_),
    .B(_05179_),
    .C(_05180_),
    .Y(_05181_));
 sky130_fd_sc_hd__a21o_1 _12599_ (.A1(_05176_),
    .A2(_05180_),
    .B1(_05179_),
    .X(_05182_));
 sky130_fd_sc_hd__nand2_1 _12600_ (.A(_03490_),
    .B(_04535_),
    .Y(_05183_));
 sky130_fd_sc_hd__clkbuf_4 _12601_ (.A(_04522_),
    .X(_05184_));
 sky130_fd_sc_hd__a22oi_1 _12602_ (.A1(_02900_),
    .A2(_04520_),
    .B1(_05184_),
    .B2(_03634_),
    .Y(_05185_));
 sky130_fd_sc_hd__and4_1 _12603_ (.A(_02894_),
    .B(_02896_),
    .C(_04520_),
    .D(_04522_),
    .X(_05186_));
 sky130_fd_sc_hd__nor2_1 _12604_ (.A(_05185_),
    .B(_05186_),
    .Y(_05187_));
 sky130_fd_sc_hd__xnor2_1 _12605_ (.A(_05183_),
    .B(_05187_),
    .Y(_05188_));
 sky130_fd_sc_hd__nand3_1 _12606_ (.A(_05181_),
    .B(_05182_),
    .C(_05188_),
    .Y(_05189_));
 sky130_fd_sc_hd__nand2_1 _12607_ (.A(_05181_),
    .B(_05189_),
    .Y(_05190_));
 sky130_fd_sc_hd__nand3_1 _12608_ (.A(_05078_),
    .B(_05075_),
    .C(_05076_),
    .Y(_05191_));
 sky130_fd_sc_hd__o21bai_1 _12609_ (.A1(_05174_),
    .A2(_05175_),
    .B1_N(_05173_),
    .Y(_05192_));
 sky130_fd_sc_hd__a22o_1 _12610_ (.A1(_02927_),
    .A2(_05184_),
    .B1(_05078_),
    .B2(_05076_),
    .X(_05193_));
 sky130_fd_sc_hd__nand3_1 _12611_ (.A(_05191_),
    .B(_05192_),
    .C(_05193_),
    .Y(_05194_));
 sky130_fd_sc_hd__a21o_1 _12612_ (.A1(_05191_),
    .A2(_05193_),
    .B1(_05192_),
    .X(_05195_));
 sky130_fd_sc_hd__nand2_1 _12613_ (.A(_03491_),
    .B(_04448_),
    .Y(_05196_));
 sky130_fd_sc_hd__buf_2 _12614_ (.A(_04520_),
    .X(_05197_));
 sky130_fd_sc_hd__a22oi_1 _12615_ (.A1(_02897_),
    .A2(_05084_),
    .B1(_05197_),
    .B2(_02895_),
    .Y(_05198_));
 sky130_fd_sc_hd__and4_1 _12616_ (.A(_03634_),
    .B(_02900_),
    .C(_05084_),
    .D(_05197_),
    .X(_05199_));
 sky130_fd_sc_hd__nor2_1 _12617_ (.A(_05198_),
    .B(_05199_),
    .Y(_05200_));
 sky130_fd_sc_hd__xnor2_1 _12618_ (.A(_05196_),
    .B(_05200_),
    .Y(_05201_));
 sky130_fd_sc_hd__nand3_1 _12619_ (.A(_05194_),
    .B(_05195_),
    .C(_05201_),
    .Y(_05202_));
 sky130_fd_sc_hd__and2_1 _12620_ (.A(_05154_),
    .B(_05157_),
    .X(_05203_));
 sky130_fd_sc_hd__a21o_1 _12621_ (.A1(_05194_),
    .A2(_05195_),
    .B1(_05201_),
    .X(_05204_));
 sky130_fd_sc_hd__nand3_1 _12622_ (.A(_05202_),
    .B(_05203_),
    .C(_05204_),
    .Y(_05205_));
 sky130_fd_sc_hd__a21o_1 _12623_ (.A1(_05202_),
    .A2(_05204_),
    .B1(_05203_),
    .X(_05206_));
 sky130_fd_sc_hd__nand3_1 _12624_ (.A(_05190_),
    .B(_05205_),
    .C(_05206_),
    .Y(_05207_));
 sky130_fd_sc_hd__a21o_1 _12625_ (.A1(_05205_),
    .A2(_05206_),
    .B1(_05190_),
    .X(_05208_));
 sky130_fd_sc_hd__and3_1 _12626_ (.A(_05172_),
    .B(_05207_),
    .C(_05208_),
    .X(_05209_));
 sky130_fd_sc_hd__nand2_1 _12627_ (.A(_05146_),
    .B(_05161_),
    .Y(_05210_));
 sky130_fd_sc_hd__or2b_1 _12628_ (.A(_05162_),
    .B_N(_05169_),
    .X(_05211_));
 sky130_fd_sc_hd__o22a_2 _12629_ (.A1(_05122_),
    .A2(_05123_),
    .B1(_05124_),
    .B2(_05125_),
    .X(_05212_));
 sky130_fd_sc_hd__a211oi_4 _12630_ (.A1(_05210_),
    .A2(_05211_),
    .B1(_05212_),
    .C1(_05126_),
    .Y(_05213_));
 sky130_fd_sc_hd__o211a_1 _12631_ (.A1(_05126_),
    .A2(_05212_),
    .B1(_05211_),
    .C1(_05210_),
    .X(_05214_));
 sky130_fd_sc_hd__and2_1 _12632_ (.A(_05166_),
    .B(_05168_),
    .X(_05215_));
 sky130_fd_sc_hd__a21o_1 _12633_ (.A1(_05081_),
    .A2(_05082_),
    .B1(_05088_),
    .X(_05216_));
 sky130_fd_sc_hd__nand3_1 _12634_ (.A(_05089_),
    .B(_05215_),
    .C(_05216_),
    .Y(_05217_));
 sky130_fd_sc_hd__a21o_1 _12635_ (.A1(_05089_),
    .A2(_05216_),
    .B1(_05215_),
    .X(_05218_));
 sky130_fd_sc_hd__nand2_1 _12636_ (.A(_05194_),
    .B(_05202_),
    .Y(_05219_));
 sky130_fd_sc_hd__a21oi_1 _12637_ (.A1(_05217_),
    .A2(_05218_),
    .B1(_05219_),
    .Y(_05220_));
 sky130_fd_sc_hd__and3_1 _12638_ (.A(_05217_),
    .B(_05219_),
    .C(_05218_),
    .X(_05221_));
 sky130_fd_sc_hd__o22ai_2 _12639_ (.A1(_05213_),
    .A2(_05214_),
    .B1(_05220_),
    .B2(_05221_),
    .Y(_05222_));
 sky130_fd_sc_hd__or4_1 _12640_ (.A(_05221_),
    .B(_05213_),
    .C(_05214_),
    .D(_05220_),
    .X(_05223_));
 sky130_fd_sc_hd__o211a_1 _12641_ (.A1(_05171_),
    .A2(_05209_),
    .B1(_05222_),
    .C1(_05223_),
    .X(_05224_));
 sky130_fd_sc_hd__a211oi_1 _12642_ (.A1(_05223_),
    .A2(_05222_),
    .B1(_05209_),
    .C1(_05171_),
    .Y(_05225_));
 sky130_fd_sc_hd__a31o_1 _12643_ (.A1(_03945_),
    .A2(_04535_),
    .A3(_05187_),
    .B1(_05186_),
    .X(_05226_));
 sky130_fd_sc_hd__nand2_1 _12644_ (.A(_03948_),
    .B(_04551_),
    .Y(_05227_));
 sky130_fd_sc_hd__xnor2_1 _12645_ (.A(_05226_),
    .B(_05227_),
    .Y(_05228_));
 sky130_fd_sc_hd__and3_1 _12646_ (.A(_03954_),
    .B(_04616_),
    .C(_05228_),
    .X(_05229_));
 sky130_fd_sc_hd__a31o_1 _12647_ (.A1(_04081_),
    .A2(_04551_),
    .A3(_05226_),
    .B1(_05229_),
    .X(_05230_));
 sky130_fd_sc_hd__a21bo_1 _12648_ (.A1(_05190_),
    .A2(_05206_),
    .B1_N(_05205_),
    .X(_05231_));
 sky130_fd_sc_hd__a31o_1 _12649_ (.A1(_03492_),
    .A2(_04448_),
    .A3(_05200_),
    .B1(_05199_),
    .X(_05232_));
 sky130_fd_sc_hd__nand2_1 _12650_ (.A(_03942_),
    .B(_04286_),
    .Y(_05233_));
 sky130_fd_sc_hd__xnor2_1 _12651_ (.A(_05232_),
    .B(_05233_),
    .Y(_05234_));
 sky130_fd_sc_hd__and3_1 _12652_ (.A(_02908_),
    .B(_04535_),
    .C(_05234_),
    .X(_05235_));
 sky130_fd_sc_hd__a21oi_1 _12653_ (.A1(_03959_),
    .A2(_04535_),
    .B1(_05234_),
    .Y(_05236_));
 sky130_fd_sc_hd__nor2_1 _12654_ (.A(_05235_),
    .B(_05236_),
    .Y(_05237_));
 sky130_fd_sc_hd__xor2_1 _12655_ (.A(_05231_),
    .B(_05237_),
    .X(_05238_));
 sky130_fd_sc_hd__xnor2_1 _12656_ (.A(_05230_),
    .B(_05238_),
    .Y(_05239_));
 sky130_fd_sc_hd__nor3_1 _12657_ (.A(_05224_),
    .B(_05225_),
    .C(_05239_),
    .Y(_05240_));
 sky130_fd_sc_hd__nor4_1 _12658_ (.A(_05221_),
    .B(_05213_),
    .C(_05214_),
    .D(_05220_),
    .Y(_05241_));
 sky130_fd_sc_hd__o22ai_4 _12659_ (.A1(_05129_),
    .A2(_05130_),
    .B1(_05131_),
    .B2(_05132_),
    .Y(_05242_));
 sky130_fd_sc_hd__o211a_1 _12660_ (.A1(_05213_),
    .A2(_05241_),
    .B1(_05242_),
    .C1(_05133_),
    .X(_05243_));
 sky130_fd_sc_hd__a211oi_1 _12661_ (.A1(_05133_),
    .A2(_05242_),
    .B1(_05241_),
    .C1(_05213_),
    .Y(_05244_));
 sky130_fd_sc_hd__a31o_1 _12662_ (.A1(_03944_),
    .A2(_04286_),
    .A3(_05232_),
    .B1(_05235_),
    .X(_05245_));
 sky130_fd_sc_hd__a21boi_1 _12663_ (.A1(_05219_),
    .A2(_05218_),
    .B1_N(_05217_),
    .Y(_05246_));
 sky130_fd_sc_hd__a21oi_1 _12664_ (.A1(_02908_),
    .A2(_04448_),
    .B1(_05109_),
    .Y(_05247_));
 sky130_fd_sc_hd__nor2_1 _12665_ (.A(_05110_),
    .B(_05247_),
    .Y(_05248_));
 sky130_fd_sc_hd__xnor2_1 _12666_ (.A(_05246_),
    .B(_05248_),
    .Y(_05249_));
 sky130_fd_sc_hd__xnor2_1 _12667_ (.A(_05245_),
    .B(_05249_),
    .Y(_05250_));
 sky130_fd_sc_hd__o21ai_1 _12668_ (.A1(_05243_),
    .A2(_05244_),
    .B1(_05250_),
    .Y(_05251_));
 sky130_fd_sc_hd__or3_1 _12669_ (.A(_05243_),
    .B(_05244_),
    .C(_05250_),
    .X(_05252_));
 sky130_fd_sc_hd__o211a_1 _12670_ (.A1(_05224_),
    .A2(_05240_),
    .B1(_05251_),
    .C1(_05252_),
    .X(_05253_));
 sky130_fd_sc_hd__inv_2 _12671_ (.A(_05253_),
    .Y(_05254_));
 sky130_fd_sc_hd__nand2_1 _12672_ (.A(_05231_),
    .B(_05237_),
    .Y(_05255_));
 sky130_fd_sc_hd__nand2_1 _12673_ (.A(_05230_),
    .B(_05238_),
    .Y(_05256_));
 sky130_fd_sc_hd__a211oi_1 _12674_ (.A1(_05252_),
    .A2(_05251_),
    .B1(_05240_),
    .C1(_05224_),
    .Y(_05257_));
 sky130_fd_sc_hd__a211o_1 _12675_ (.A1(_05255_),
    .A2(_05256_),
    .B1(_05253_),
    .C1(_05257_),
    .X(_05258_));
 sky130_fd_sc_hd__or3_2 _12676_ (.A(_05110_),
    .B(_05246_),
    .C(_05247_),
    .X(_05259_));
 sky130_fd_sc_hd__nand2_1 _12677_ (.A(_05245_),
    .B(_05249_),
    .Y(_05260_));
 sky130_fd_sc_hd__nor3_1 _12678_ (.A(_05243_),
    .B(_05244_),
    .C(_05250_),
    .Y(_05261_));
 sky130_fd_sc_hd__o21ai_1 _12679_ (.A1(_05135_),
    .A2(_05136_),
    .B1(_05137_),
    .Y(_05262_));
 sky130_fd_sc_hd__or3_1 _12680_ (.A(_05135_),
    .B(_05136_),
    .C(_05137_),
    .X(_05263_));
 sky130_fd_sc_hd__o211a_2 _12681_ (.A1(_05243_),
    .A2(_05261_),
    .B1(_05262_),
    .C1(_05263_),
    .X(_05264_));
 sky130_fd_sc_hd__a211oi_2 _12682_ (.A1(_05263_),
    .A2(_05262_),
    .B1(_05261_),
    .C1(_05243_),
    .Y(_05265_));
 sky130_fd_sc_hd__a211oi_4 _12683_ (.A1(_05259_),
    .A2(_05260_),
    .B1(_05264_),
    .C1(_05265_),
    .Y(_05266_));
 sky130_fd_sc_hd__o211a_1 _12684_ (.A1(_05264_),
    .A2(_05265_),
    .B1(_05259_),
    .C1(_05260_),
    .X(_05267_));
 sky130_fd_sc_hd__a211oi_1 _12685_ (.A1(_05254_),
    .A2(_05258_),
    .B1(_05266_),
    .C1(_05267_),
    .Y(_05268_));
 sky130_fd_sc_hd__a211oi_1 _12686_ (.A1(_05116_),
    .A2(_05117_),
    .B1(_05138_),
    .C1(_05135_),
    .Y(_05269_));
 sky130_fd_sc_hd__o21bai_1 _12687_ (.A1(_05140_),
    .A2(_05269_),
    .B1_N(_05115_),
    .Y(_05270_));
 sky130_fd_sc_hd__a211o_1 _12688_ (.A1(_05106_),
    .A2(_05114_),
    .B1(_05140_),
    .C1(_05269_),
    .X(_05271_));
 sky130_fd_sc_hd__o211a_1 _12689_ (.A1(_05264_),
    .A2(_05266_),
    .B1(_05270_),
    .C1(_05271_),
    .X(_05272_));
 sky130_fd_sc_hd__a211o_1 _12690_ (.A1(_05271_),
    .A2(_05270_),
    .B1(_05266_),
    .C1(_05264_),
    .X(_05273_));
 sky130_fd_sc_hd__o21ai_1 _12691_ (.A1(_05268_),
    .A2(_05272_),
    .B1(_05273_),
    .Y(_05274_));
 sky130_fd_sc_hd__a21oi_1 _12692_ (.A1(_05070_),
    .A2(_05142_),
    .B1(_05069_),
    .Y(_05275_));
 sky130_fd_sc_hd__o31ai_2 _12693_ (.A1(_05071_),
    .A2(_05144_),
    .A3(_05274_),
    .B1(_05275_),
    .Y(_05276_));
 sky130_fd_sc_hd__o21ba_1 _12694_ (.A1(_04918_),
    .A2(_04995_),
    .B1_N(_04917_),
    .X(_05277_));
 sky130_fd_sc_hd__o21ba_1 _12695_ (.A1(_04759_),
    .A2(_04837_),
    .B1_N(_04758_),
    .X(_05278_));
 sky130_fd_sc_hd__a31o_1 _12696_ (.A1(_04760_),
    .A2(_04839_),
    .A3(_05277_),
    .B1(_05278_),
    .X(_05279_));
 sky130_fd_sc_hd__a21oi_2 _12697_ (.A1(_04998_),
    .A2(_05276_),
    .B1(_05279_),
    .Y(_05280_));
 sky130_fd_sc_hd__and2_1 _12698_ (.A(_04511_),
    .B(_04596_),
    .X(_05281_));
 sky130_fd_sc_hd__nor3b_2 _12699_ (.A(_04595_),
    .B(_04598_),
    .C_N(_04675_),
    .Y(_05282_));
 sky130_fd_sc_hd__o21ba_1 _12700_ (.A1(_04511_),
    .A2(_04596_),
    .B1_N(_05282_),
    .X(_05283_));
 sky130_fd_sc_hd__o21ai_1 _12701_ (.A1(_04423_),
    .A2(_04507_),
    .B1(_04424_),
    .Y(_05284_));
 sky130_fd_sc_hd__o41a_1 _12702_ (.A1(_04425_),
    .A2(_04509_),
    .A3(_05281_),
    .A4(_05283_),
    .B1(_05284_),
    .X(_05285_));
 sky130_fd_sc_hd__or4_1 _12703_ (.A(_04183_),
    .B(_04264_),
    .C(_04345_),
    .D(_05285_),
    .X(_05286_));
 sky130_fd_sc_hd__and2b_1 _12704_ (.A_N(_04344_),
    .B(_04266_),
    .X(_05287_));
 sky130_fd_sc_hd__o21ai_1 _12705_ (.A1(_04262_),
    .A2(_05287_),
    .B1(_04261_),
    .Y(_05288_));
 sky130_fd_sc_hd__nor2_1 _12706_ (.A(_04099_),
    .B(_04180_),
    .Y(_05289_));
 sky130_fd_sc_hd__o22a_1 _12707_ (.A1(_04183_),
    .A2(_05288_),
    .B1(_05289_),
    .B2(_04100_),
    .X(_05290_));
 sky130_fd_sc_hd__o211a_1 _12708_ (.A1(_04678_),
    .A2(_05280_),
    .B1(_05286_),
    .C1(_05290_),
    .X(_05291_));
 sky130_fd_sc_hd__clkbuf_4 _12709_ (.A(_05118_),
    .X(_05292_));
 sky130_fd_sc_hd__and4_1 _12710_ (.A(_03302_),
    .B(_03239_),
    .C(_05292_),
    .D(_05145_),
    .X(_05293_));
 sky130_fd_sc_hd__a22oi_1 _12711_ (.A1(_03239_),
    .A2(_05292_),
    .B1(_05145_),
    .B2(_03302_),
    .Y(_05294_));
 sky130_fd_sc_hd__and4bb_1 _12712_ (.A_N(_05293_),
    .B_N(_05294_),
    .C(_03434_),
    .D(_05197_),
    .X(_05295_));
 sky130_fd_sc_hd__o2bb2a_1 _12713_ (.A1_N(_03434_),
    .A2_N(_05197_),
    .B1(_05293_),
    .B2(_05294_),
    .X(_05296_));
 sky130_fd_sc_hd__nor2_1 _12714_ (.A(_05295_),
    .B(_05296_),
    .Y(_05297_));
 sky130_fd_sc_hd__and4_1 _12715_ (.A(_03142_),
    .B(_03434_),
    .C(_05184_),
    .D(_05147_),
    .X(_05298_));
 sky130_fd_sc_hd__and2_1 _12716_ (.A(_05297_),
    .B(_05298_),
    .X(_05299_));
 sky130_fd_sc_hd__nor2_1 _12717_ (.A(_05297_),
    .B(_05298_),
    .Y(_05300_));
 sky130_fd_sc_hd__or2_1 _12718_ (.A(_05299_),
    .B(_05300_),
    .X(_05301_));
 sky130_fd_sc_hd__nand4_1 _12719_ (.A(_03208_),
    .B(_03531_),
    .C(_05118_),
    .D(_04967_),
    .Y(_05302_));
 sky130_fd_sc_hd__a22o_1 _12720_ (.A1(_03212_),
    .A2(_04944_),
    .B1(_04967_),
    .B2(_03217_),
    .X(_05303_));
 sky130_fd_sc_hd__nand4_1 _12721_ (.A(_02917_),
    .B(_05093_),
    .C(_05302_),
    .D(_05303_),
    .Y(_05304_));
 sky130_fd_sc_hd__and2_1 _12722_ (.A(_05302_),
    .B(_05304_),
    .X(_05305_));
 sky130_fd_sc_hd__and4_1 _12723_ (.A(_03532_),
    .B(_03531_),
    .C(_04686_),
    .D(_05118_),
    .X(_05306_));
 sky130_fd_sc_hd__a22oi_1 _12724_ (.A1(_03213_),
    .A2(_05093_),
    .B1(_05118_),
    .B2(_03218_),
    .Y(_05307_));
 sky130_fd_sc_hd__and4bb_1 _12725_ (.A_N(_05306_),
    .B_N(_05307_),
    .C(_02917_),
    .D(_05092_),
    .X(_05308_));
 sky130_fd_sc_hd__o2bb2a_1 _12726_ (.A1_N(_02917_),
    .A2_N(_05167_),
    .B1(_05306_),
    .B2(_05307_),
    .X(_05309_));
 sky130_fd_sc_hd__nor2_1 _12727_ (.A(_05308_),
    .B(_05309_),
    .Y(_05310_));
 sky130_fd_sc_hd__and2b_1 _12728_ (.A_N(_05305_),
    .B(_05310_),
    .X(_05311_));
 sky130_fd_sc_hd__xnor2_1 _12729_ (.A(_05305_),
    .B(_05310_),
    .Y(_05312_));
 sky130_fd_sc_hd__nand2_1 _12730_ (.A(_03491_),
    .B(_05197_),
    .Y(_05313_));
 sky130_fd_sc_hd__and3_1 _12731_ (.A(_03634_),
    .B(_02900_),
    .C(_05077_),
    .X(_05314_));
 sky130_fd_sc_hd__a22o_1 _12732_ (.A1(_02900_),
    .A2(_05077_),
    .B1(_04643_),
    .B2(_03634_),
    .X(_05315_));
 sky130_fd_sc_hd__a21bo_1 _12733_ (.A1(_05163_),
    .A2(_05314_),
    .B1_N(_05315_),
    .X(_05316_));
 sky130_fd_sc_hd__xor2_1 _12734_ (.A(_05313_),
    .B(_05316_),
    .X(_05317_));
 sky130_fd_sc_hd__and2_1 _12735_ (.A(_05312_),
    .B(_05317_),
    .X(_05318_));
 sky130_fd_sc_hd__nor2_1 _12736_ (.A(_05306_),
    .B(_05308_),
    .Y(_05319_));
 sky130_fd_sc_hd__nand2_1 _12737_ (.A(_02927_),
    .B(_05163_),
    .Y(_05320_));
 sky130_fd_sc_hd__and4_1 _12738_ (.A(_03532_),
    .B(_03531_),
    .C(_04681_),
    .D(_04686_),
    .X(_05321_));
 sky130_fd_sc_hd__a22o_1 _12739_ (.A1(_03531_),
    .A2(_05092_),
    .B1(_05093_),
    .B2(_03208_),
    .X(_05322_));
 sky130_fd_sc_hd__and2b_1 _12740_ (.A_N(_05321_),
    .B(_05322_),
    .X(_05323_));
 sky130_fd_sc_hd__xnor2_1 _12741_ (.A(_05320_),
    .B(_05323_),
    .Y(_05324_));
 sky130_fd_sc_hd__xnor2_1 _12742_ (.A(_05319_),
    .B(_05324_),
    .Y(_05325_));
 sky130_fd_sc_hd__nand2_1 _12743_ (.A(_03491_),
    .B(_05084_),
    .Y(_05326_));
 sky130_fd_sc_hd__clkbuf_4 _12744_ (.A(_04524_),
    .X(_05327_));
 sky130_fd_sc_hd__a22o_1 _12745_ (.A1(_02897_),
    .A2(_05327_),
    .B1(_05077_),
    .B2(_03634_),
    .X(_05328_));
 sky130_fd_sc_hd__a21bo_1 _12746_ (.A1(_05327_),
    .A2(_05314_),
    .B1_N(_05328_),
    .X(_05329_));
 sky130_fd_sc_hd__xor2_1 _12747_ (.A(_05326_),
    .B(_05329_),
    .X(_05330_));
 sky130_fd_sc_hd__xor2_1 _12748_ (.A(_05325_),
    .B(_05330_),
    .X(_05331_));
 sky130_fd_sc_hd__o21a_1 _12749_ (.A1(_05311_),
    .A2(_05318_),
    .B1(_05331_),
    .X(_05332_));
 sky130_fd_sc_hd__nor3_1 _12750_ (.A(_05331_),
    .B(_05311_),
    .C(_05318_),
    .Y(_05333_));
 sky130_fd_sc_hd__nor3_2 _12751_ (.A(_05301_),
    .B(_05332_),
    .C(_05333_),
    .Y(_05334_));
 sky130_fd_sc_hd__and2b_1 _12752_ (.A_N(_05319_),
    .B(_05324_),
    .X(_05335_));
 sky130_fd_sc_hd__and2_1 _12753_ (.A(_05325_),
    .B(_05330_),
    .X(_05336_));
 sky130_fd_sc_hd__a31o_1 _12754_ (.A1(_02918_),
    .A2(_05163_),
    .A3(_05322_),
    .B1(_05321_),
    .X(_05337_));
 sky130_fd_sc_hd__nand2_1 _12755_ (.A(_02927_),
    .B(_05077_),
    .Y(_05338_));
 sky130_fd_sc_hd__and2b_1 _12756_ (.A_N(_05178_),
    .B(_05177_),
    .X(_05339_));
 sky130_fd_sc_hd__xnor2_1 _12757_ (.A(_05338_),
    .B(_05339_),
    .Y(_05340_));
 sky130_fd_sc_hd__xor2_1 _12758_ (.A(_05337_),
    .B(_05340_),
    .X(_05341_));
 sky130_fd_sc_hd__nand2_1 _12759_ (.A(_03945_),
    .B(_04616_),
    .Y(_05342_));
 sky130_fd_sc_hd__a22oi_1 _12760_ (.A1(_02900_),
    .A2(_04522_),
    .B1(_05327_),
    .B2(_03634_),
    .Y(_05343_));
 sky130_fd_sc_hd__and4_1 _12761_ (.A(_03872_),
    .B(_03873_),
    .C(_04522_),
    .D(_04524_),
    .X(_05344_));
 sky130_fd_sc_hd__nor2_1 _12762_ (.A(_05343_),
    .B(_05344_),
    .Y(_05345_));
 sky130_fd_sc_hd__xnor2_1 _12763_ (.A(_05342_),
    .B(_05345_),
    .Y(_05346_));
 sky130_fd_sc_hd__xor2_1 _12764_ (.A(_05341_),
    .B(_05346_),
    .X(_05347_));
 sky130_fd_sc_hd__o21ai_2 _12765_ (.A1(_05335_),
    .A2(_05336_),
    .B1(_05347_),
    .Y(_05348_));
 sky130_fd_sc_hd__or3_1 _12766_ (.A(_05347_),
    .B(_05335_),
    .C(_05336_),
    .X(_05349_));
 sky130_fd_sc_hd__nand2_1 _12767_ (.A(_03434_),
    .B(_05084_),
    .Y(_05350_));
 sky130_fd_sc_hd__nand2_1 _12768_ (.A(_02935_),
    .B(_05093_),
    .Y(_05351_));
 sky130_fd_sc_hd__and2b_1 _12769_ (.A_N(_05156_),
    .B(_05155_),
    .X(_05352_));
 sky130_fd_sc_hd__xnor2_2 _12770_ (.A(_05351_),
    .B(_05352_),
    .Y(_05353_));
 sky130_fd_sc_hd__xnor2_1 _12771_ (.A(_05293_),
    .B(_05353_),
    .Y(_05354_));
 sky130_fd_sc_hd__xor2_1 _12772_ (.A(_05350_),
    .B(_05354_),
    .X(_05355_));
 sky130_fd_sc_hd__xor2_1 _12773_ (.A(_05295_),
    .B(_05355_),
    .X(_05356_));
 sky130_fd_sc_hd__a21o_1 _12774_ (.A1(_05348_),
    .A2(_05349_),
    .B1(_05356_),
    .X(_05357_));
 sky130_fd_sc_hd__nand3_2 _12775_ (.A(_05356_),
    .B(_05348_),
    .C(_05349_),
    .Y(_05358_));
 sky130_fd_sc_hd__o211a_2 _12776_ (.A1(_05299_),
    .A2(_05334_),
    .B1(_05357_),
    .C1(_05358_),
    .X(_05359_));
 sky130_fd_sc_hd__a211oi_2 _12777_ (.A1(_05358_),
    .A2(_05357_),
    .B1(_05334_),
    .C1(_05299_),
    .Y(_05360_));
 sky130_fd_sc_hd__a32o_1 _12778_ (.A1(_03945_),
    .A2(_05197_),
    .A3(_05315_),
    .B1(_05314_),
    .B2(_05163_),
    .X(_05361_));
 sky130_fd_sc_hd__nand2_1 _12779_ (.A(_03942_),
    .B(_04616_),
    .Y(_05362_));
 sky130_fd_sc_hd__xnor2_1 _12780_ (.A(_05361_),
    .B(_05362_),
    .Y(_05363_));
 sky130_fd_sc_hd__and3_1 _12781_ (.A(_03954_),
    .B(_05184_),
    .C(_05363_),
    .X(_05364_));
 sky130_fd_sc_hd__a31o_1 _12782_ (.A1(_04081_),
    .A2(_04616_),
    .A3(_05361_),
    .B1(_05364_),
    .X(_05365_));
 sky130_fd_sc_hd__a32o_1 _12783_ (.A1(_03945_),
    .A2(_05084_),
    .A3(_05328_),
    .B1(_05314_),
    .B2(_05327_),
    .X(_05366_));
 sky130_fd_sc_hd__nand2_1 _12784_ (.A(_03942_),
    .B(_04535_),
    .Y(_05367_));
 sky130_fd_sc_hd__xnor2_1 _12785_ (.A(_05366_),
    .B(_05367_),
    .Y(_05368_));
 sky130_fd_sc_hd__and3_1 _12786_ (.A(_03954_),
    .B(_05197_),
    .C(_05368_),
    .X(_05369_));
 sky130_fd_sc_hd__a21oi_1 _12787_ (.A1(_03959_),
    .A2(_05197_),
    .B1(_05368_),
    .Y(_05370_));
 sky130_fd_sc_hd__nor2_1 _12788_ (.A(_05369_),
    .B(_05370_),
    .Y(_05371_));
 sky130_fd_sc_hd__xor2_1 _12789_ (.A(_05332_),
    .B(_05371_),
    .X(_05372_));
 sky130_fd_sc_hd__xnor2_1 _12790_ (.A(_05365_),
    .B(_05372_),
    .Y(_05373_));
 sky130_fd_sc_hd__nor3_4 _12791_ (.A(_05359_),
    .B(_05360_),
    .C(_05373_),
    .Y(_05374_));
 sky130_fd_sc_hd__nand2_1 _12792_ (.A(_05295_),
    .B(_05355_),
    .Y(_05375_));
 sky130_fd_sc_hd__and2_1 _12793_ (.A(_05337_),
    .B(_05340_),
    .X(_05376_));
 sky130_fd_sc_hd__a21o_1 _12794_ (.A1(_05341_),
    .A2(_05346_),
    .B1(_05376_),
    .X(_05377_));
 sky130_fd_sc_hd__and2_1 _12795_ (.A(_05293_),
    .B(_05353_),
    .X(_05378_));
 sky130_fd_sc_hd__a21o_1 _12796_ (.A1(_05181_),
    .A2(_05182_),
    .B1(_05188_),
    .X(_05379_));
 sky130_fd_sc_hd__nand3_1 _12797_ (.A(_05189_),
    .B(_05378_),
    .C(_05379_),
    .Y(_05380_));
 sky130_fd_sc_hd__a21o_1 _12798_ (.A1(_05189_),
    .A2(_05379_),
    .B1(_05378_),
    .X(_05381_));
 sky130_fd_sc_hd__nand3_1 _12799_ (.A(_05377_),
    .B(_05380_),
    .C(_05381_),
    .Y(_05382_));
 sky130_fd_sc_hd__a21o_1 _12800_ (.A1(_05380_),
    .A2(_05381_),
    .B1(_05377_),
    .X(_05383_));
 sky130_fd_sc_hd__or2_1 _12801_ (.A(_05350_),
    .B(_05354_),
    .X(_05384_));
 sky130_fd_sc_hd__xnor2_1 _12802_ (.A(_05149_),
    .B(_05158_),
    .Y(_05385_));
 sky130_fd_sc_hd__xnor2_1 _12803_ (.A(_05384_),
    .B(_05385_),
    .Y(_05386_));
 sky130_fd_sc_hd__a21oi_1 _12804_ (.A1(_05382_),
    .A2(_05383_),
    .B1(_05386_),
    .Y(_05387_));
 sky130_fd_sc_hd__and3_1 _12805_ (.A(_05386_),
    .B(_05382_),
    .C(_05383_),
    .X(_05388_));
 sky130_fd_sc_hd__a211oi_2 _12806_ (.A1(_05375_),
    .A2(_05358_),
    .B1(_05387_),
    .C1(_05388_),
    .Y(_05389_));
 sky130_fd_sc_hd__o211a_1 _12807_ (.A1(_05388_),
    .A2(_05387_),
    .B1(_05358_),
    .C1(_05375_),
    .X(_05390_));
 sky130_fd_sc_hd__a31o_1 _12808_ (.A1(_03944_),
    .A2(_04535_),
    .A3(_05366_),
    .B1(_05369_),
    .X(_05391_));
 sky130_fd_sc_hd__a31o_1 _12809_ (.A1(_03491_),
    .A2(_04616_),
    .A3(_05345_),
    .B1(_05344_),
    .X(_05392_));
 sky130_fd_sc_hd__nand2_1 _12810_ (.A(_02887_),
    .B(_04448_),
    .Y(_05393_));
 sky130_fd_sc_hd__xnor2_1 _12811_ (.A(_05392_),
    .B(_05393_),
    .Y(_05394_));
 sky130_fd_sc_hd__and3_1 _12812_ (.A(_03947_),
    .B(_05084_),
    .C(_05394_),
    .X(_05395_));
 sky130_fd_sc_hd__a21oi_1 _12813_ (.A1(_03954_),
    .A2(_05084_),
    .B1(_05394_),
    .Y(_05396_));
 sky130_fd_sc_hd__nor2_1 _12814_ (.A(_05395_),
    .B(_05396_),
    .Y(_05397_));
 sky130_fd_sc_hd__xnor2_1 _12815_ (.A(_05348_),
    .B(_05397_),
    .Y(_05398_));
 sky130_fd_sc_hd__xnor2_1 _12816_ (.A(_05391_),
    .B(_05398_),
    .Y(_05399_));
 sky130_fd_sc_hd__o21ai_1 _12817_ (.A1(_05389_),
    .A2(_05390_),
    .B1(_05399_),
    .Y(_05400_));
 sky130_fd_sc_hd__or3_1 _12818_ (.A(_05389_),
    .B(_05390_),
    .C(_05399_),
    .X(_05401_));
 sky130_fd_sc_hd__o211ai_2 _12819_ (.A1(_05359_),
    .A2(_05374_),
    .B1(_05400_),
    .C1(_05401_),
    .Y(_05402_));
 sky130_fd_sc_hd__and2_1 _12820_ (.A(_05332_),
    .B(_05371_),
    .X(_05403_));
 sky130_fd_sc_hd__a21oi_1 _12821_ (.A1(_05365_),
    .A2(_05372_),
    .B1(_05403_),
    .Y(_05404_));
 sky130_fd_sc_hd__a211o_1 _12822_ (.A1(_05401_),
    .A2(_05400_),
    .B1(_05374_),
    .C1(_05359_),
    .X(_05405_));
 sky130_fd_sc_hd__nand2_1 _12823_ (.A(_05402_),
    .B(_05405_),
    .Y(_05406_));
 sky130_fd_sc_hd__or2_1 _12824_ (.A(_05404_),
    .B(_05406_),
    .X(_05407_));
 sky130_fd_sc_hd__or3_1 _12825_ (.A(_05395_),
    .B(_05348_),
    .C(_05396_),
    .X(_05408_));
 sky130_fd_sc_hd__nand2_1 _12826_ (.A(_05391_),
    .B(_05398_),
    .Y(_05409_));
 sky130_fd_sc_hd__nor3_1 _12827_ (.A(_05389_),
    .B(_05390_),
    .C(_05399_),
    .Y(_05410_));
 sky130_fd_sc_hd__or2b_1 _12828_ (.A(_05384_),
    .B_N(_05385_),
    .X(_05411_));
 sky130_fd_sc_hd__nand3_1 _12829_ (.A(_05386_),
    .B(_05382_),
    .C(_05383_),
    .Y(_05412_));
 sky130_fd_sc_hd__a21oi_1 _12830_ (.A1(_05207_),
    .A2(_05208_),
    .B1(_05172_),
    .Y(_05413_));
 sky130_fd_sc_hd__a211oi_2 _12831_ (.A1(_05411_),
    .A2(_05412_),
    .B1(_05413_),
    .C1(_05209_),
    .Y(_05414_));
 sky130_fd_sc_hd__o211a_1 _12832_ (.A1(_05209_),
    .A2(_05413_),
    .B1(_05412_),
    .C1(_05411_),
    .X(_05415_));
 sky130_fd_sc_hd__a31o_1 _12833_ (.A1(_03944_),
    .A2(_04448_),
    .A3(_05392_),
    .B1(_05395_),
    .X(_05416_));
 sky130_fd_sc_hd__a21bo_1 _12834_ (.A1(_05377_),
    .A2(_05381_),
    .B1_N(_05380_),
    .X(_05417_));
 sky130_fd_sc_hd__a21oi_1 _12835_ (.A1(_03959_),
    .A2(_04616_),
    .B1(_05228_),
    .Y(_05418_));
 sky130_fd_sc_hd__nor2_1 _12836_ (.A(_05229_),
    .B(_05418_),
    .Y(_05419_));
 sky130_fd_sc_hd__xor2_1 _12837_ (.A(_05417_),
    .B(_05419_),
    .X(_05420_));
 sky130_fd_sc_hd__xnor2_1 _12838_ (.A(_05416_),
    .B(_05420_),
    .Y(_05421_));
 sky130_fd_sc_hd__o21ai_1 _12839_ (.A1(_05414_),
    .A2(_05415_),
    .B1(_05421_),
    .Y(_05422_));
 sky130_fd_sc_hd__or3_1 _12840_ (.A(_05414_),
    .B(_05415_),
    .C(_05421_),
    .X(_05423_));
 sky130_fd_sc_hd__o211a_1 _12841_ (.A1(_05389_),
    .A2(_05410_),
    .B1(_05422_),
    .C1(_05423_),
    .X(_05424_));
 sky130_fd_sc_hd__a211oi_1 _12842_ (.A1(_05423_),
    .A2(_05422_),
    .B1(_05410_),
    .C1(_05389_),
    .Y(_05425_));
 sky130_fd_sc_hd__a211oi_2 _12843_ (.A1(_05408_),
    .A2(_05409_),
    .B1(_05424_),
    .C1(_05425_),
    .Y(_05426_));
 sky130_fd_sc_hd__o211a_1 _12844_ (.A1(_05424_),
    .A2(_05425_),
    .B1(_05408_),
    .C1(_05409_),
    .X(_05427_));
 sky130_fd_sc_hd__a211oi_1 _12845_ (.A1(_05402_),
    .A2(_05407_),
    .B1(_05426_),
    .C1(_05427_),
    .Y(_05428_));
 sky130_fd_sc_hd__o211a_1 _12846_ (.A1(_05426_),
    .A2(_05427_),
    .B1(_05402_),
    .C1(_05407_),
    .X(_05429_));
 sky130_fd_sc_hd__or2_1 _12847_ (.A(_05428_),
    .B(_05429_),
    .X(_05430_));
 sky130_fd_sc_hd__xnor2_1 _12848_ (.A(_05404_),
    .B(_05406_),
    .Y(_05431_));
 sky130_fd_sc_hd__o21a_1 _12849_ (.A1(_05332_),
    .A2(_05333_),
    .B1(_05301_),
    .X(_05432_));
 sky130_fd_sc_hd__a22oi_1 _12850_ (.A1(_03435_),
    .A2(_05184_),
    .B1(_05147_),
    .B2(_03142_),
    .Y(_05433_));
 sky130_fd_sc_hd__nor2_1 _12851_ (.A(_05298_),
    .B(_05433_),
    .Y(_05434_));
 sky130_fd_sc_hd__xor2_1 _12852_ (.A(_05312_),
    .B(_05317_),
    .X(_05435_));
 sky130_fd_sc_hd__a22o_1 _12853_ (.A1(_02917_),
    .A2(_05093_),
    .B1(_05302_),
    .B2(_05303_),
    .X(_05436_));
 sky130_fd_sc_hd__and4_1 _12854_ (.A(_03213_),
    .B(_02926_),
    .C(_05118_),
    .D(_04967_),
    .X(_05437_));
 sky130_fd_sc_hd__and3_1 _12855_ (.A(_05304_),
    .B(_05436_),
    .C(_05437_),
    .X(_05438_));
 sky130_fd_sc_hd__a21oi_1 _12856_ (.A1(_05304_),
    .A2(_05436_),
    .B1(_05437_),
    .Y(_05439_));
 sky130_fd_sc_hd__nand2_1 _12857_ (.A(_02892_),
    .B(_05184_),
    .Y(_05440_));
 sky130_fd_sc_hd__a22oi_1 _12858_ (.A1(_03873_),
    .A2(_04643_),
    .B1(_05092_),
    .B2(_02894_),
    .Y(_05441_));
 sky130_fd_sc_hd__and4_1 _12859_ (.A(_03633_),
    .B(_03637_),
    .C(_04643_),
    .D(_05092_),
    .X(_05442_));
 sky130_fd_sc_hd__nor2_1 _12860_ (.A(_05441_),
    .B(_05442_),
    .Y(_05443_));
 sky130_fd_sc_hd__xnor2_1 _12861_ (.A(_05440_),
    .B(_05443_),
    .Y(_05444_));
 sky130_fd_sc_hd__nor3b_1 _12862_ (.A(_05438_),
    .B(_05439_),
    .C_N(_05444_),
    .Y(_05445_));
 sky130_fd_sc_hd__nor2_1 _12863_ (.A(_05438_),
    .B(_05445_),
    .Y(_05446_));
 sky130_fd_sc_hd__xnor2_1 _12864_ (.A(_05435_),
    .B(_05446_),
    .Y(_05447_));
 sky130_fd_sc_hd__and2_1 _12865_ (.A(_05434_),
    .B(_05447_),
    .X(_05448_));
 sky130_fd_sc_hd__or3b_4 _12866_ (.A(_05334_),
    .B(_05432_),
    .C_N(_05448_),
    .X(_05449_));
 sky130_fd_sc_hd__o21bai_2 _12867_ (.A1(_05334_),
    .A2(_05432_),
    .B1_N(_05448_),
    .Y(_05450_));
 sky130_fd_sc_hd__a31o_1 _12868_ (.A1(_03491_),
    .A2(_05184_),
    .A3(_05443_),
    .B1(_05442_),
    .X(_05451_));
 sky130_fd_sc_hd__nand2_1 _12869_ (.A(_03948_),
    .B(_05084_),
    .Y(_05452_));
 sky130_fd_sc_hd__xnor2_1 _12870_ (.A(_05451_),
    .B(_05452_),
    .Y(_05453_));
 sky130_fd_sc_hd__and3_1 _12871_ (.A(_03947_),
    .B(_05327_),
    .C(_05453_),
    .X(_05454_));
 sky130_fd_sc_hd__a31oi_4 _12872_ (.A1(_04081_),
    .A2(_05084_),
    .A3(_05451_),
    .B1(_05454_),
    .Y(_05455_));
 sky130_fd_sc_hd__or2b_1 _12873_ (.A(_05446_),
    .B_N(_05435_),
    .X(_05456_));
 sky130_fd_sc_hd__a21oi_1 _12874_ (.A1(_03959_),
    .A2(_05184_),
    .B1(_05363_),
    .Y(_05457_));
 sky130_fd_sc_hd__nor2_1 _12875_ (.A(_05364_),
    .B(_05457_),
    .Y(_05458_));
 sky130_fd_sc_hd__xnor2_1 _12876_ (.A(_05456_),
    .B(_05458_),
    .Y(_05459_));
 sky130_fd_sc_hd__xnor2_2 _12877_ (.A(_05455_),
    .B(_05459_),
    .Y(_05460_));
 sky130_fd_sc_hd__nand3_4 _12878_ (.A(_05449_),
    .B(_05450_),
    .C(_05460_),
    .Y(_05461_));
 sky130_fd_sc_hd__o21a_1 _12879_ (.A1(_05359_),
    .A2(_05360_),
    .B1(_05373_),
    .X(_05462_));
 sky130_fd_sc_hd__a211oi_4 _12880_ (.A1(_05449_),
    .A2(_05461_),
    .B1(_05462_),
    .C1(_05374_),
    .Y(_05463_));
 sky130_fd_sc_hd__or3_2 _12881_ (.A(_05364_),
    .B(_05456_),
    .C(_05457_),
    .X(_05464_));
 sky130_fd_sc_hd__or2b_1 _12882_ (.A(_05455_),
    .B_N(_05459_),
    .X(_05465_));
 sky130_fd_sc_hd__o211a_1 _12883_ (.A1(_05374_),
    .A2(_05462_),
    .B1(_05461_),
    .C1(_05449_),
    .X(_05466_));
 sky130_fd_sc_hd__a211oi_4 _12884_ (.A1(_05464_),
    .A2(_05465_),
    .B1(_05463_),
    .C1(_05466_),
    .Y(_05467_));
 sky130_fd_sc_hd__nor2_1 _12885_ (.A(_05463_),
    .B(_05467_),
    .Y(_05468_));
 sky130_fd_sc_hd__nor2_1 _12886_ (.A(_05431_),
    .B(_05468_),
    .Y(_05469_));
 sky130_fd_sc_hd__and2_1 _12887_ (.A(_05431_),
    .B(_05468_),
    .X(_05470_));
 sky130_fd_sc_hd__or2_1 _12888_ (.A(_05469_),
    .B(_05470_),
    .X(_05471_));
 sky130_fd_sc_hd__o211a_1 _12889_ (.A1(_05463_),
    .A2(_05466_),
    .B1(_05464_),
    .C1(_05465_),
    .X(_05472_));
 sky130_fd_sc_hd__xnor2_2 _12890_ (.A(_05434_),
    .B(_05447_),
    .Y(_05473_));
 sky130_fd_sc_hd__o21ba_1 _12891_ (.A1(_05438_),
    .A2(_05439_),
    .B1_N(_05444_),
    .X(_05474_));
 sky130_fd_sc_hd__a22oi_1 _12892_ (.A1(_02917_),
    .A2(_05292_),
    .B1(_05145_),
    .B2(_02923_),
    .Y(_05475_));
 sky130_fd_sc_hd__nor2_1 _12893_ (.A(_05437_),
    .B(_05475_),
    .Y(_05476_));
 sky130_fd_sc_hd__nand2_1 _12894_ (.A(\wfg_stim_mem_top.cfg_gain_q[9] ),
    .B(_04524_),
    .Y(_05477_));
 sky130_fd_sc_hd__a22oi_2 _12895_ (.A1(_02899_),
    .A2(_05092_),
    .B1(_05093_),
    .B2(_03633_),
    .Y(_05478_));
 sky130_fd_sc_hd__and4_2 _12896_ (.A(\wfg_stim_mem_top.cfg_gain_q[13] ),
    .B(_02899_),
    .C(_04681_),
    .D(_04686_),
    .X(_05479_));
 sky130_fd_sc_hd__or3_1 _12897_ (.A(_05477_),
    .B(_05478_),
    .C(_05479_),
    .X(_05480_));
 sky130_fd_sc_hd__o21ai_1 _12898_ (.A1(_05478_),
    .A2(_05479_),
    .B1(_05477_),
    .Y(_05481_));
 sky130_fd_sc_hd__nand3_2 _12899_ (.A(_05476_),
    .B(_05480_),
    .C(_05481_),
    .Y(_05482_));
 sky130_fd_sc_hd__or3_2 _12900_ (.A(_05445_),
    .B(_05474_),
    .C(_05482_),
    .X(_05483_));
 sky130_fd_sc_hd__o21ai_2 _12901_ (.A1(_05445_),
    .A2(_05474_),
    .B1(_05482_),
    .Y(_05484_));
 sky130_fd_sc_hd__nand4_4 _12902_ (.A(_03435_),
    .B(_05327_),
    .C(_05483_),
    .D(_05484_),
    .Y(_05485_));
 sky130_fd_sc_hd__nor2_1 _12903_ (.A(_05473_),
    .B(_05485_),
    .Y(_05486_));
 sky130_fd_sc_hd__xor2_2 _12904_ (.A(_05473_),
    .B(_05485_),
    .X(_05487_));
 sky130_fd_sc_hd__a21oi_1 _12905_ (.A1(_02908_),
    .A2(_05327_),
    .B1(_05453_),
    .Y(_05488_));
 sky130_fd_sc_hd__nor2_1 _12906_ (.A(_05454_),
    .B(_05488_),
    .Y(_05489_));
 sky130_fd_sc_hd__xnor2_1 _12907_ (.A(_05483_),
    .B(_05489_),
    .Y(_05490_));
 sky130_fd_sc_hd__nand2_1 _12908_ (.A(_02906_),
    .B(_05077_),
    .Y(_05491_));
 sky130_fd_sc_hd__nor3_1 _12909_ (.A(_05477_),
    .B(_05478_),
    .C(_05479_),
    .Y(_05492_));
 sky130_fd_sc_hd__a211oi_1 _12910_ (.A1(_02887_),
    .A2(_05197_),
    .B1(_05479_),
    .C1(_05492_),
    .Y(_05493_));
 sky130_fd_sc_hd__o211a_1 _12911_ (.A1(_05479_),
    .A2(_05492_),
    .B1(_02886_),
    .C1(_05197_),
    .X(_05494_));
 sky130_fd_sc_hd__o21ba_1 _12912_ (.A1(_05491_),
    .A2(_05493_),
    .B1_N(_05494_),
    .X(_05495_));
 sky130_fd_sc_hd__xnor2_1 _12913_ (.A(_05490_),
    .B(_05495_),
    .Y(_05496_));
 sky130_fd_sc_hd__and2_1 _12914_ (.A(_05487_),
    .B(_05496_),
    .X(_05497_));
 sky130_fd_sc_hd__a21o_1 _12915_ (.A1(_05449_),
    .A2(_05450_),
    .B1(_05460_),
    .X(_05498_));
 sky130_fd_sc_hd__o211ai_4 _12916_ (.A1(_05486_),
    .A2(_05497_),
    .B1(_05498_),
    .C1(_05461_),
    .Y(_05499_));
 sky130_fd_sc_hd__and2b_1 _12917_ (.A_N(_05483_),
    .B(_05489_),
    .X(_05500_));
 sky130_fd_sc_hd__and2b_1 _12918_ (.A_N(_05495_),
    .B(_05490_),
    .X(_05501_));
 sky130_fd_sc_hd__a211o_1 _12919_ (.A1(_05461_),
    .A2(_05498_),
    .B1(_05497_),
    .C1(_05486_),
    .X(_05502_));
 sky130_fd_sc_hd__o211ai_4 _12920_ (.A1(_05500_),
    .A2(_05501_),
    .B1(_05499_),
    .C1(_05502_),
    .Y(_05503_));
 sky130_fd_sc_hd__o211a_2 _12921_ (.A1(_05467_),
    .A2(_05472_),
    .B1(_05499_),
    .C1(_05503_),
    .X(_05504_));
 sky130_fd_sc_hd__a211o_1 _12922_ (.A1(_05499_),
    .A2(_05502_),
    .B1(_05500_),
    .C1(_05501_),
    .X(_05505_));
 sky130_fd_sc_hd__nand2_2 _12923_ (.A(_05503_),
    .B(_05505_),
    .Y(_05506_));
 sky130_fd_sc_hd__nand2_1 _12924_ (.A(\wfg_stim_mem_top.cfg_gain_q[9] ),
    .B(_04512_),
    .Y(_05507_));
 sky130_fd_sc_hd__a22oi_2 _12925_ (.A1(_02899_),
    .A2(_05093_),
    .B1(_05118_),
    .B2(_03633_),
    .Y(_05508_));
 sky130_fd_sc_hd__and4_1 _12926_ (.A(\wfg_stim_mem_top.cfg_gain_q[13] ),
    .B(\wfg_stim_mem_top.cfg_gain_q[12] ),
    .C(_04686_),
    .D(_04944_),
    .X(_05509_));
 sky130_fd_sc_hd__or3_2 _12927_ (.A(_05507_),
    .B(_05508_),
    .C(_05509_),
    .X(_05510_));
 sky130_fd_sc_hd__o21ai_2 _12928_ (.A1(_05508_),
    .A2(_05509_),
    .B1(_05507_),
    .Y(_05511_));
 sky130_fd_sc_hd__nand4_2 _12929_ (.A(_02918_),
    .B(_05147_),
    .C(_05510_),
    .D(_05511_),
    .Y(_05512_));
 sky130_fd_sc_hd__a21o_1 _12930_ (.A1(_05480_),
    .A2(_05481_),
    .B1(_05476_),
    .X(_05513_));
 sky130_fd_sc_hd__and3b_1 _12931_ (.A_N(_05512_),
    .B(_05513_),
    .C(_05482_),
    .X(_05514_));
 sky130_fd_sc_hd__nor2_1 _12932_ (.A(_05494_),
    .B(_05493_),
    .Y(_05515_));
 sky130_fd_sc_hd__xnor2_2 _12933_ (.A(_05491_),
    .B(_05515_),
    .Y(_05516_));
 sky130_fd_sc_hd__nand2_1 _12934_ (.A(_02906_),
    .B(_05163_),
    .Y(_05517_));
 sky130_fd_sc_hd__o21bai_2 _12935_ (.A1(_05507_),
    .A2(_05508_),
    .B1_N(_05509_),
    .Y(_05518_));
 sky130_fd_sc_hd__a21oi_2 _12936_ (.A1(_03948_),
    .A2(_05184_),
    .B1(_05518_),
    .Y(_05519_));
 sky130_fd_sc_hd__and3_1 _12937_ (.A(_02887_),
    .B(_05184_),
    .C(_05518_),
    .X(_05520_));
 sky130_fd_sc_hd__o21ba_1 _12938_ (.A1(_05517_),
    .A2(_05519_),
    .B1_N(_05520_),
    .X(_05521_));
 sky130_fd_sc_hd__xor2_1 _12939_ (.A(_05514_),
    .B(_05516_),
    .X(_05522_));
 sky130_fd_sc_hd__or2b_1 _12940_ (.A(_05521_),
    .B_N(_05522_),
    .X(_05523_));
 sky130_fd_sc_hd__a21bo_1 _12941_ (.A1(_05514_),
    .A2(_05516_),
    .B1_N(_05523_),
    .X(_05524_));
 sky130_fd_sc_hd__a22o_1 _12942_ (.A1(_03435_),
    .A2(_05327_),
    .B1(_05483_),
    .B2(_05484_),
    .X(_05525_));
 sky130_fd_sc_hd__nand2_1 _12943_ (.A(_03435_),
    .B(_05077_),
    .Y(_05526_));
 sky130_fd_sc_hd__a21boi_1 _12944_ (.A1(_05482_),
    .A2(_05513_),
    .B1_N(_05512_),
    .Y(_05527_));
 sky130_fd_sc_hd__or3_1 _12945_ (.A(_05526_),
    .B(_05514_),
    .C(_05527_),
    .X(_05528_));
 sky130_fd_sc_hd__a21bo_1 _12946_ (.A1(_05485_),
    .A2(_05525_),
    .B1_N(_05528_),
    .X(_05529_));
 sky130_fd_sc_hd__xnor2_1 _12947_ (.A(_05521_),
    .B(_05522_),
    .Y(_05530_));
 sky130_fd_sc_hd__nand3b_1 _12948_ (.A_N(_05528_),
    .B(_05525_),
    .C(_05485_),
    .Y(_05531_));
 sky130_fd_sc_hd__a21bo_1 _12949_ (.A1(_05529_),
    .A2(_05530_),
    .B1_N(_05531_),
    .X(_05532_));
 sky130_fd_sc_hd__xor2_2 _12950_ (.A(_05487_),
    .B(_05496_),
    .X(_05533_));
 sky130_fd_sc_hd__or2_1 _12951_ (.A(_05532_),
    .B(_05533_),
    .X(_05534_));
 sky130_fd_sc_hd__nand2_1 _12952_ (.A(_05532_),
    .B(_05533_),
    .Y(_05535_));
 sky130_fd_sc_hd__a21bo_1 _12953_ (.A1(_05524_),
    .A2(_05534_),
    .B1_N(_05535_),
    .X(_05536_));
 sky130_fd_sc_hd__xor2_1 _12954_ (.A(_05506_),
    .B(_05536_),
    .X(_05537_));
 sky130_fd_sc_hd__xnor2_1 _12955_ (.A(_05532_),
    .B(_05533_),
    .Y(_05538_));
 sky130_fd_sc_hd__xnor2_1 _12956_ (.A(_05524_),
    .B(_05538_),
    .Y(_05539_));
 sky130_fd_sc_hd__a22o_1 _12957_ (.A1(_02918_),
    .A2(_05147_),
    .B1(_05510_),
    .B2(_05511_),
    .X(_05540_));
 sky130_fd_sc_hd__nand4_2 _12958_ (.A(_03435_),
    .B(_05163_),
    .C(_05512_),
    .D(_05540_),
    .Y(_05541_));
 sky130_fd_sc_hd__o21ai_1 _12959_ (.A1(_05514_),
    .A2(_05527_),
    .B1(_05526_),
    .Y(_05542_));
 sky130_fd_sc_hd__nand3b_1 _12960_ (.A_N(_05541_),
    .B(_05542_),
    .C(_05528_),
    .Y(_05543_));
 sky130_fd_sc_hd__a21bo_1 _12961_ (.A1(_05528_),
    .A2(_05542_),
    .B1_N(_05541_),
    .X(_05544_));
 sky130_fd_sc_hd__nor2_1 _12962_ (.A(_05520_),
    .B(_05519_),
    .Y(_05545_));
 sky130_fd_sc_hd__xnor2_1 _12963_ (.A(_05517_),
    .B(_05545_),
    .Y(_05546_));
 sky130_fd_sc_hd__and2_1 _12964_ (.A(\wfg_stim_mem_top.cfg_gain_q[9] ),
    .B(_04643_),
    .X(_05547_));
 sky130_fd_sc_hd__a22o_1 _12965_ (.A1(_02899_),
    .A2(_05118_),
    .B1(_04967_),
    .B2(_03633_),
    .X(_05548_));
 sky130_fd_sc_hd__nand4_2 _12966_ (.A(_03636_),
    .B(_03637_),
    .C(_05118_),
    .D(_04967_),
    .Y(_05549_));
 sky130_fd_sc_hd__a21bo_1 _12967_ (.A1(_05547_),
    .A2(_05548_),
    .B1_N(_05549_),
    .X(_05550_));
 sky130_fd_sc_hd__nand2_1 _12968_ (.A(_02886_),
    .B(_05327_),
    .Y(_05551_));
 sky130_fd_sc_hd__xnor2_1 _12969_ (.A(_05550_),
    .B(_05551_),
    .Y(_05552_));
 sky130_fd_sc_hd__and3_1 _12970_ (.A(_03942_),
    .B(_05327_),
    .C(_05550_),
    .X(_05553_));
 sky130_fd_sc_hd__a31oi_2 _12971_ (.A1(_03947_),
    .A2(_05167_),
    .A3(_05552_),
    .B1(_05553_),
    .Y(_05554_));
 sky130_fd_sc_hd__xnor2_1 _12972_ (.A(_05546_),
    .B(_05554_),
    .Y(_05555_));
 sky130_fd_sc_hd__nand3_1 _12973_ (.A(_05543_),
    .B(_05544_),
    .C(_05555_),
    .Y(_05556_));
 sky130_fd_sc_hd__a21oi_1 _12974_ (.A1(_05531_),
    .A2(_05529_),
    .B1(_05530_),
    .Y(_05557_));
 sky130_fd_sc_hd__and3_1 _12975_ (.A(_05531_),
    .B(_05529_),
    .C(_05530_),
    .X(_05558_));
 sky130_fd_sc_hd__a211oi_1 _12976_ (.A1(_05543_),
    .A2(_05556_),
    .B1(_05557_),
    .C1(_05558_),
    .Y(_05559_));
 sky130_fd_sc_hd__or2b_1 _12977_ (.A(_05554_),
    .B_N(_05546_),
    .X(_05560_));
 sky130_fd_sc_hd__o211a_1 _12978_ (.A1(_05558_),
    .A2(_05557_),
    .B1(_05556_),
    .C1(_05543_),
    .X(_05561_));
 sky130_fd_sc_hd__or3_1 _12979_ (.A(_05560_),
    .B(_05559_),
    .C(_05561_),
    .X(_05562_));
 sky130_fd_sc_hd__and2b_1 _12980_ (.A_N(_05559_),
    .B(_05562_),
    .X(_05563_));
 sky130_fd_sc_hd__xnor2_1 _12981_ (.A(_05539_),
    .B(_05563_),
    .Y(_05564_));
 sky130_fd_sc_hd__o21ai_1 _12982_ (.A1(_05559_),
    .A2(_05561_),
    .B1(_05560_),
    .Y(_05565_));
 sky130_fd_sc_hd__a22o_1 _12983_ (.A1(_03434_),
    .A2(_05163_),
    .B1(_05512_),
    .B2(_05540_),
    .X(_05566_));
 sky130_fd_sc_hd__nand3_1 _12984_ (.A(_05549_),
    .B(_05547_),
    .C(_05548_),
    .Y(_05567_));
 sky130_fd_sc_hd__a21o_1 _12985_ (.A1(_05549_),
    .A2(_05548_),
    .B1(_05547_),
    .X(_05568_));
 sky130_fd_sc_hd__and4_1 _12986_ (.A(_03434_),
    .B(_05167_),
    .C(_05567_),
    .D(_05568_),
    .X(_05569_));
 sky130_fd_sc_hd__nand3_1 _12987_ (.A(_05541_),
    .B(_05566_),
    .C(_05569_),
    .Y(_05570_));
 sky130_fd_sc_hd__inv_2 _12988_ (.A(_05570_),
    .Y(_05571_));
 sky130_fd_sc_hd__a21o_1 _12989_ (.A1(_05541_),
    .A2(_05566_),
    .B1(_05569_),
    .X(_05572_));
 sky130_fd_sc_hd__nand2_1 _12990_ (.A(_02906_),
    .B(_05167_),
    .Y(_05573_));
 sky130_fd_sc_hd__xnor2_1 _12991_ (.A(_05573_),
    .B(_05552_),
    .Y(_05574_));
 sky130_fd_sc_hd__clkbuf_4 _12992_ (.A(_05093_),
    .X(_05575_));
 sky130_fd_sc_hd__and4_1 _12993_ (.A(_02900_),
    .B(\wfg_stim_mem_top.cfg_gain_q[9] ),
    .C(_05092_),
    .D(_05145_),
    .X(_05576_));
 sky130_fd_sc_hd__nand2_1 _12994_ (.A(_02886_),
    .B(_05077_),
    .Y(_05577_));
 sky130_fd_sc_hd__xnor2_1 _12995_ (.A(_05576_),
    .B(_05577_),
    .Y(_05578_));
 sky130_fd_sc_hd__and3_1 _12996_ (.A(_02886_),
    .B(_05077_),
    .C(_05576_),
    .X(_05579_));
 sky130_fd_sc_hd__a31oi_2 _12997_ (.A1(_02906_),
    .A2(_05575_),
    .A3(_05578_),
    .B1(_05579_),
    .Y(_05580_));
 sky130_fd_sc_hd__xnor2_1 _12998_ (.A(_05574_),
    .B(_05580_),
    .Y(_05581_));
 sky130_fd_sc_hd__and3_1 _12999_ (.A(_05570_),
    .B(_05572_),
    .C(_05581_),
    .X(_05582_));
 sky130_fd_sc_hd__a21o_1 _13000_ (.A1(_05543_),
    .A2(_05544_),
    .B1(_05555_),
    .X(_05583_));
 sky130_fd_sc_hd__o211a_1 _13001_ (.A1(_05571_),
    .A2(_05582_),
    .B1(_05583_),
    .C1(_05556_),
    .X(_05584_));
 sky130_fd_sc_hd__or2b_1 _13002_ (.A(_05580_),
    .B_N(_05574_),
    .X(_05585_));
 sky130_fd_sc_hd__a211oi_1 _13003_ (.A1(_05556_),
    .A2(_05583_),
    .B1(_05582_),
    .C1(_05571_),
    .Y(_05586_));
 sky130_fd_sc_hd__or3_1 _13004_ (.A(_05585_),
    .B(_05584_),
    .C(_05586_),
    .X(_05587_));
 sky130_fd_sc_hd__or2b_1 _13005_ (.A(_05584_),
    .B_N(_05587_),
    .X(_05588_));
 sky130_fd_sc_hd__a21o_1 _13006_ (.A1(_05562_),
    .A2(_05565_),
    .B1(_05588_),
    .X(_05589_));
 sky130_fd_sc_hd__o21ai_1 _13007_ (.A1(_05584_),
    .A2(_05586_),
    .B1(_05585_),
    .Y(_05590_));
 sky130_fd_sc_hd__nand4_1 _13008_ (.A(_03435_),
    .B(_05167_),
    .C(_05567_),
    .D(_05568_),
    .Y(_05591_));
 sky130_fd_sc_hd__a22o_1 _13009_ (.A1(_03434_),
    .A2(_05167_),
    .B1(_05567_),
    .B2(_05568_),
    .X(_05592_));
 sky130_fd_sc_hd__nand2_1 _13010_ (.A(_03434_),
    .B(_05575_),
    .Y(_05593_));
 sky130_fd_sc_hd__a22oi_1 _13011_ (.A1(_03869_),
    .A2(_05167_),
    .B1(_05145_),
    .B2(_02897_),
    .Y(_05594_));
 sky130_fd_sc_hd__or2_1 _13012_ (.A(_05576_),
    .B(_05594_),
    .X(_05595_));
 sky130_fd_sc_hd__nor2_1 _13013_ (.A(_05593_),
    .B(_05595_),
    .Y(_05596_));
 sky130_fd_sc_hd__nand3_1 _13014_ (.A(_05591_),
    .B(_05592_),
    .C(_05596_),
    .Y(_05597_));
 sky130_fd_sc_hd__nand2_1 _13015_ (.A(_02906_),
    .B(_05575_),
    .Y(_05598_));
 sky130_fd_sc_hd__xnor2_1 _13016_ (.A(_05598_),
    .B(_05578_),
    .Y(_05599_));
 sky130_fd_sc_hd__and4_2 _13017_ (.A(\wfg_stim_mem_top.cfg_gain_q[11] ),
    .B(\wfg_stim_mem_top.cfg_gain_q[8] ),
    .C(_05163_),
    .D(_05292_),
    .X(_05600_));
 sky130_fd_sc_hd__xor2_1 _13018_ (.A(_05599_),
    .B(_05600_),
    .X(_05601_));
 sky130_fd_sc_hd__a21o_1 _13019_ (.A1(_05591_),
    .A2(_05592_),
    .B1(_05596_),
    .X(_05602_));
 sky130_fd_sc_hd__nand3_1 _13020_ (.A(_05597_),
    .B(_05601_),
    .C(_05602_),
    .Y(_05603_));
 sky130_fd_sc_hd__a21oi_1 _13021_ (.A1(_05570_),
    .A2(_05572_),
    .B1(_05581_),
    .Y(_05604_));
 sky130_fd_sc_hd__a211oi_1 _13022_ (.A1(_05597_),
    .A2(_05603_),
    .B1(_05582_),
    .C1(_05604_),
    .Y(_05605_));
 sky130_fd_sc_hd__nand2_1 _13023_ (.A(_05599_),
    .B(_05600_),
    .Y(_05606_));
 sky130_fd_sc_hd__o211a_1 _13024_ (.A1(_05582_),
    .A2(_05604_),
    .B1(_05597_),
    .C1(_05603_),
    .X(_05607_));
 sky130_fd_sc_hd__or3_1 _13025_ (.A(_05606_),
    .B(_05605_),
    .C(_05607_),
    .X(_05608_));
 sky130_fd_sc_hd__or2b_1 _13026_ (.A(_05605_),
    .B_N(_05608_),
    .X(_05609_));
 sky130_fd_sc_hd__a21o_1 _13027_ (.A1(_05587_),
    .A2(_05590_),
    .B1(_05609_),
    .X(_05610_));
 sky130_fd_sc_hd__o21ai_1 _13028_ (.A1(_05605_),
    .A2(_05607_),
    .B1(_05606_),
    .Y(_05611_));
 sky130_fd_sc_hd__a21o_1 _13029_ (.A1(_05597_),
    .A2(_05602_),
    .B1(_05601_),
    .X(_05612_));
 sky130_fd_sc_hd__and3_1 _13030_ (.A(_03069_),
    .B(\wfg_stim_mem_top.cfg_gain_q[9] ),
    .C(_05118_),
    .X(_05613_));
 sky130_fd_sc_hd__a21oi_1 _13031_ (.A1(_03492_),
    .A2(_05292_),
    .B1(_05593_),
    .Y(_05614_));
 sky130_fd_sc_hd__xnor2_1 _13032_ (.A(_05595_),
    .B(_05614_),
    .Y(_05615_));
 sky130_fd_sc_hd__a22oi_1 _13033_ (.A1(_02886_),
    .A2(_05163_),
    .B1(_05292_),
    .B2(_02906_),
    .Y(_05616_));
 sky130_fd_sc_hd__or2_1 _13034_ (.A(_05600_),
    .B(_05616_),
    .X(_05617_));
 sky130_fd_sc_hd__and4_1 _13035_ (.A(_02906_),
    .B(_02886_),
    .C(_05167_),
    .D(_05145_),
    .X(_05618_));
 sky130_fd_sc_hd__xnor2_1 _13036_ (.A(_05617_),
    .B(_05618_),
    .Y(_05619_));
 sky130_fd_sc_hd__a32o_1 _13037_ (.A1(_05575_),
    .A2(_05595_),
    .A3(_05613_),
    .B1(_05615_),
    .B2(_05619_),
    .X(_05620_));
 sky130_fd_sc_hd__nand3_1 _13038_ (.A(_05603_),
    .B(_05612_),
    .C(_05620_),
    .Y(_05621_));
 sky130_fd_sc_hd__and2b_1 _13039_ (.A_N(_05617_),
    .B(_05618_),
    .X(_05622_));
 sky130_fd_sc_hd__a21o_1 _13040_ (.A1(_05603_),
    .A2(_05612_),
    .B1(_05620_),
    .X(_05623_));
 sky130_fd_sc_hd__nand3_1 _13041_ (.A(_05622_),
    .B(_05621_),
    .C(_05623_),
    .Y(_05624_));
 sky130_fd_sc_hd__nand2_1 _13042_ (.A(_05621_),
    .B(_05624_),
    .Y(_05625_));
 sky130_fd_sc_hd__a21oi_1 _13043_ (.A1(_05608_),
    .A2(_05611_),
    .B1(_05625_),
    .Y(_05626_));
 sky130_fd_sc_hd__a21o_1 _13044_ (.A1(_05621_),
    .A2(_05623_),
    .B1(_05622_),
    .X(_05627_));
 sky130_fd_sc_hd__xnor2_1 _13045_ (.A(_05619_),
    .B(_05615_),
    .Y(_05628_));
 sky130_fd_sc_hd__nand2_1 _13046_ (.A(_05147_),
    .B(_05613_),
    .Y(_05629_));
 sky130_fd_sc_hd__a22oi_1 _13047_ (.A1(_02886_),
    .A2(_05167_),
    .B1(_05147_),
    .B2(_02906_),
    .Y(_05630_));
 sky130_fd_sc_hd__or2_1 _13048_ (.A(_05618_),
    .B(_05630_),
    .X(_05631_));
 sky130_fd_sc_hd__and3b_1 _13049_ (.A_N(_05145_),
    .B(_05613_),
    .C(_05575_),
    .X(_05632_));
 sky130_fd_sc_hd__nand2_1 _13050_ (.A(_03490_),
    .B(_05145_),
    .Y(_05633_));
 sky130_fd_sc_hd__a32o_1 _13051_ (.A1(_03069_),
    .A2(_05292_),
    .A3(_05633_),
    .B1(_03869_),
    .B2(_05575_),
    .X(_05634_));
 sky130_fd_sc_hd__and2b_1 _13052_ (.A_N(_05632_),
    .B(_05634_),
    .X(_05635_));
 sky130_fd_sc_hd__or2b_1 _13053_ (.A(_05631_),
    .B_N(_05635_),
    .X(_05636_));
 sky130_fd_sc_hd__o21a_1 _13054_ (.A1(_05575_),
    .A2(_05629_),
    .B1(_05636_),
    .X(_05637_));
 sky130_fd_sc_hd__nor2_1 _13055_ (.A(_05628_),
    .B(_05637_),
    .Y(_05638_));
 sky130_fd_sc_hd__a21o_1 _13056_ (.A1(_05624_),
    .A2(_05627_),
    .B1(_05638_),
    .X(_05639_));
 sky130_fd_sc_hd__xnor2_2 _13057_ (.A(_05631_),
    .B(_05635_),
    .Y(_05640_));
 sky130_fd_sc_hd__xnor2_1 _13058_ (.A(_05628_),
    .B(_05637_),
    .Y(_05641_));
 sky130_fd_sc_hd__a22o_1 _13059_ (.A1(_03492_),
    .A2(_05292_),
    .B1(_05147_),
    .B2(_03435_),
    .X(_05642_));
 sky130_fd_sc_hd__and4_1 _13060_ (.A(_03942_),
    .B(_05575_),
    .C(_05629_),
    .D(_05642_),
    .X(_05643_));
 sky130_fd_sc_hd__nand2_1 _13061_ (.A(_05640_),
    .B(_05643_),
    .Y(_05644_));
 sky130_fd_sc_hd__xor2_1 _13062_ (.A(_05641_),
    .B(_05644_),
    .X(_05645_));
 sky130_fd_sc_hd__nand4_1 _13063_ (.A(_03944_),
    .B(_05575_),
    .C(_05629_),
    .D(_05642_),
    .Y(_05646_));
 sky130_fd_sc_hd__a22o_1 _13064_ (.A1(_03943_),
    .A2(_05575_),
    .B1(_05629_),
    .B2(_05642_),
    .X(_05647_));
 sky130_fd_sc_hd__and4_1 _13065_ (.A(_03492_),
    .B(_03943_),
    .C(_05292_),
    .D(_05147_),
    .X(_05648_));
 sky130_fd_sc_hd__and3_1 _13066_ (.A(_05646_),
    .B(_05647_),
    .C(_05648_),
    .X(_05649_));
 sky130_fd_sc_hd__nor2_1 _13067_ (.A(_05641_),
    .B(_05644_),
    .Y(_05650_));
 sky130_fd_sc_hd__a31o_1 _13068_ (.A1(_05640_),
    .A2(_05645_),
    .A3(_05649_),
    .B1(_05650_),
    .X(_05651_));
 sky130_fd_sc_hd__and3_1 _13069_ (.A(_05624_),
    .B(_05627_),
    .C(_05638_),
    .X(_05652_));
 sky130_fd_sc_hd__a21oi_1 _13070_ (.A1(_05639_),
    .A2(_05651_),
    .B1(_05652_),
    .Y(_05653_));
 sky130_fd_sc_hd__and3_1 _13071_ (.A(_05608_),
    .B(_05611_),
    .C(_05625_),
    .X(_05654_));
 sky130_fd_sc_hd__o21bai_1 _13072_ (.A1(_05626_),
    .A2(_05653_),
    .B1_N(_05654_),
    .Y(_05655_));
 sky130_fd_sc_hd__and3_1 _13073_ (.A(_05587_),
    .B(_05590_),
    .C(_05609_),
    .X(_05656_));
 sky130_fd_sc_hd__a21o_1 _13074_ (.A1(_05610_),
    .A2(_05655_),
    .B1(_05656_),
    .X(_05657_));
 sky130_fd_sc_hd__and3_1 _13075_ (.A(_05562_),
    .B(_05565_),
    .C(_05588_),
    .X(_05658_));
 sky130_fd_sc_hd__a21o_1 _13076_ (.A1(_05589_),
    .A2(_05657_),
    .B1(_05658_),
    .X(_05659_));
 sky130_fd_sc_hd__and2b_1 _13077_ (.A_N(_05563_),
    .B(_05539_),
    .X(_05660_));
 sky130_fd_sc_hd__a21oi_1 _13078_ (.A1(_05564_),
    .A2(_05659_),
    .B1(_05660_),
    .Y(_05661_));
 sky130_fd_sc_hd__a211oi_4 _13079_ (.A1(_05499_),
    .A2(_05503_),
    .B1(_05467_),
    .C1(_05472_),
    .Y(_05662_));
 sky130_fd_sc_hd__inv_2 _13080_ (.A(_05662_),
    .Y(_05663_));
 sky130_fd_sc_hd__or2b_1 _13081_ (.A(_05506_),
    .B_N(_05536_),
    .X(_05664_));
 sky130_fd_sc_hd__o211a_1 _13082_ (.A1(_05537_),
    .A2(_05661_),
    .B1(_05663_),
    .C1(_05664_),
    .X(_05665_));
 sky130_fd_sc_hd__or4_4 _13083_ (.A(_05430_),
    .B(_05471_),
    .C(_05504_),
    .D(_05665_),
    .X(_05666_));
 sky130_fd_sc_hd__o211ai_1 _13084_ (.A1(_05253_),
    .A2(_05257_),
    .B1(_05255_),
    .C1(_05256_),
    .Y(_05667_));
 sky130_fd_sc_hd__nand2_2 _13085_ (.A(_05258_),
    .B(_05667_),
    .Y(_05668_));
 sky130_fd_sc_hd__nand2_1 _13086_ (.A(_05417_),
    .B(_05419_),
    .Y(_05669_));
 sky130_fd_sc_hd__a21bo_1 _13087_ (.A1(_05416_),
    .A2(_05420_),
    .B1_N(_05669_),
    .X(_05670_));
 sky130_fd_sc_hd__nor3_1 _13088_ (.A(_05414_),
    .B(_05415_),
    .C(_05421_),
    .Y(_05671_));
 sky130_fd_sc_hd__o21ai_1 _13089_ (.A1(_05224_),
    .A2(_05225_),
    .B1(_05239_),
    .Y(_05672_));
 sky130_fd_sc_hd__or3_1 _13090_ (.A(_05224_),
    .B(_05225_),
    .C(_05239_),
    .X(_05673_));
 sky130_fd_sc_hd__o211a_1 _13091_ (.A1(_05414_),
    .A2(_05671_),
    .B1(_05672_),
    .C1(_05673_),
    .X(_05674_));
 sky130_fd_sc_hd__a211oi_1 _13092_ (.A1(_05673_),
    .A2(_05672_),
    .B1(_05671_),
    .C1(_05414_),
    .Y(_05675_));
 sky130_fd_sc_hd__nor2_1 _13093_ (.A(_05674_),
    .B(_05675_),
    .Y(_05676_));
 sky130_fd_sc_hd__a21oi_2 _13094_ (.A1(_05670_),
    .A2(_05676_),
    .B1(_05674_),
    .Y(_05677_));
 sky130_fd_sc_hd__nor2_1 _13095_ (.A(_05668_),
    .B(_05677_),
    .Y(_05678_));
 sky130_fd_sc_hd__xnor2_1 _13096_ (.A(_05670_),
    .B(_05676_),
    .Y(_05679_));
 sky130_fd_sc_hd__nor2_1 _13097_ (.A(_05424_),
    .B(_05426_),
    .Y(_05680_));
 sky130_fd_sc_hd__nor2_1 _13098_ (.A(_05679_),
    .B(_05680_),
    .Y(_05681_));
 sky130_fd_sc_hd__nand2_1 _13099_ (.A(_05668_),
    .B(_05677_),
    .Y(_05682_));
 sky130_fd_sc_hd__o21a_1 _13100_ (.A1(_05678_),
    .A2(_05681_),
    .B1(_05682_),
    .X(_05683_));
 sky130_fd_sc_hd__o21ba_1 _13101_ (.A1(_05428_),
    .A2(_05469_),
    .B1_N(_05429_),
    .X(_05684_));
 sky130_fd_sc_hd__nor2_2 _13102_ (.A(_05683_),
    .B(_05684_),
    .Y(_05685_));
 sky130_fd_sc_hd__nand4_2 _13103_ (.A(_04760_),
    .B(_04839_),
    .C(_04919_),
    .D(_04997_),
    .Y(_05686_));
 sky130_fd_sc_hd__nor2_2 _13104_ (.A(_05266_),
    .B(_05267_),
    .Y(_05687_));
 sky130_fd_sc_hd__nand2_1 _13105_ (.A(_05254_),
    .B(_05258_),
    .Y(_05688_));
 sky130_fd_sc_hd__xor2_4 _13106_ (.A(_05687_),
    .B(_05688_),
    .X(_05689_));
 sky130_fd_sc_hd__a211oi_1 _13107_ (.A1(_05271_),
    .A2(_05270_),
    .B1(_05266_),
    .C1(_05264_),
    .Y(_05690_));
 sky130_fd_sc_hd__nor2_2 _13108_ (.A(_05690_),
    .B(_05272_),
    .Y(_05691_));
 sky130_fd_sc_hd__or4bb_1 _13109_ (.A(_05071_),
    .B(_05144_),
    .C_N(_05689_),
    .D_N(_05691_),
    .X(_05692_));
 sky130_fd_sc_hd__or2_1 _13110_ (.A(_05686_),
    .B(_05692_),
    .X(_05693_));
 sky130_fd_sc_hd__xnor2_2 _13111_ (.A(_05668_),
    .B(_05677_),
    .Y(_05694_));
 sky130_fd_sc_hd__nand2_1 _13112_ (.A(_05679_),
    .B(_05680_),
    .Y(_05695_));
 sky130_fd_sc_hd__or2b_1 _13113_ (.A(_05681_),
    .B_N(_05695_),
    .X(_05696_));
 sky130_fd_sc_hd__o21ba_2 _13114_ (.A1(_05694_),
    .A2(_05696_),
    .B1_N(_05683_),
    .X(_05697_));
 sky130_fd_sc_hd__a2111o_2 _13115_ (.A1(_05666_),
    .A2(_05685_),
    .B1(_05693_),
    .C1(_05697_),
    .D1(_04678_),
    .X(_05698_));
 sky130_fd_sc_hd__xor2_1 _13116_ (.A(_03748_),
    .B(_03746_),
    .X(_05699_));
 sky130_fd_sc_hd__xnor2_2 _13117_ (.A(_03706_),
    .B(_03726_),
    .Y(_05700_));
 sky130_fd_sc_hd__o22a_1 _13118_ (.A1(_03692_),
    .A2(_03693_),
    .B1(_03702_),
    .B2(_03703_),
    .X(_05701_));
 sky130_fd_sc_hd__a211o_1 _13119_ (.A1(_04047_),
    .A2(_04056_),
    .B1(_03704_),
    .C1(_05701_),
    .X(_05702_));
 sky130_fd_sc_hd__o211ai_2 _13120_ (.A1(_03704_),
    .A2(_05701_),
    .B1(_04047_),
    .C1(_04056_),
    .Y(_05703_));
 sky130_fd_sc_hd__a21bo_1 _13121_ (.A1(_04049_),
    .A2(_04053_),
    .B1_N(_04052_),
    .X(_05704_));
 sky130_fd_sc_hd__a21o_1 _13122_ (.A1(_03713_),
    .A2(_03714_),
    .B1(_03718_),
    .X(_05705_));
 sky130_fd_sc_hd__and3_2 _13123_ (.A(_05704_),
    .B(_03719_),
    .C(_05705_),
    .X(_05706_));
 sky130_fd_sc_hd__a21oi_2 _13124_ (.A1(_03719_),
    .A2(_05705_),
    .B1(_05704_),
    .Y(_05707_));
 sky130_fd_sc_hd__a211o_1 _13125_ (.A1(_04064_),
    .A2(_04071_),
    .B1(_05706_),
    .C1(_05707_),
    .X(_05708_));
 sky130_fd_sc_hd__o211ai_2 _13126_ (.A1(_05706_),
    .A2(_05707_),
    .B1(_04064_),
    .C1(_04071_),
    .Y(_05709_));
 sky130_fd_sc_hd__nand4_2 _13127_ (.A(_05702_),
    .B(_05703_),
    .C(_05708_),
    .D(_05709_),
    .Y(_05710_));
 sky130_fd_sc_hd__nand2_2 _13128_ (.A(_05702_),
    .B(_05710_),
    .Y(_05711_));
 sky130_fd_sc_hd__xor2_2 _13129_ (.A(_05700_),
    .B(_05711_),
    .X(_05712_));
 sky130_fd_sc_hd__a211oi_2 _13130_ (.A1(_04064_),
    .A2(_04071_),
    .B1(_05706_),
    .C1(_05707_),
    .Y(_05713_));
 sky130_fd_sc_hd__nand2_1 _13131_ (.A(_02909_),
    .B(_02953_),
    .Y(_05714_));
 sky130_fd_sc_hd__and2b_1 _13132_ (.A_N(_03739_),
    .B(_03738_),
    .X(_05715_));
 sky130_fd_sc_hd__xnor2_1 _13133_ (.A(_05714_),
    .B(_05715_),
    .Y(_05716_));
 sky130_fd_sc_hd__o21ai_1 _13134_ (.A1(_05706_),
    .A2(_05713_),
    .B1(_05716_),
    .Y(_05717_));
 sky130_fd_sc_hd__or3_1 _13135_ (.A(_05706_),
    .B(_05713_),
    .C(_05716_),
    .X(_05718_));
 sky130_fd_sc_hd__and2_1 _13136_ (.A(_05717_),
    .B(_05718_),
    .X(_05719_));
 sky130_fd_sc_hd__nor2_1 _13137_ (.A(_04066_),
    .B(_04069_),
    .Y(_05720_));
 sky130_fd_sc_hd__or3_1 _13138_ (.A(_02891_),
    .B(_04068_),
    .C(_05720_),
    .X(_05721_));
 sky130_fd_sc_hd__o21a_1 _13139_ (.A1(_04068_),
    .A2(_05720_),
    .B1(_02891_),
    .X(_05722_));
 sky130_fd_sc_hd__a31oi_2 _13140_ (.A1(_02909_),
    .A2(_03022_),
    .A3(_05721_),
    .B1(_05722_),
    .Y(_05723_));
 sky130_fd_sc_hd__xor2_2 _13141_ (.A(_05719_),
    .B(_05723_),
    .X(_05724_));
 sky130_fd_sc_hd__or2b_1 _13142_ (.A(_05700_),
    .B_N(_05711_),
    .X(_05725_));
 sky130_fd_sc_hd__o21a_1 _13143_ (.A1(_05712_),
    .A2(_05724_),
    .B1(_05725_),
    .X(_05726_));
 sky130_fd_sc_hd__xor2_1 _13144_ (.A(_03730_),
    .B(_03741_),
    .X(_05727_));
 sky130_fd_sc_hd__or2b_1 _13145_ (.A(_05726_),
    .B_N(_05727_),
    .X(_05728_));
 sky130_fd_sc_hd__xor2_1 _13146_ (.A(_05727_),
    .B(_05726_),
    .X(_05729_));
 sky130_fd_sc_hd__or2b_1 _13147_ (.A(_05723_),
    .B_N(_05719_),
    .X(_05730_));
 sky130_fd_sc_hd__nand2_1 _13148_ (.A(_05717_),
    .B(_05730_),
    .Y(_05731_));
 sky130_fd_sc_hd__or2b_1 _13149_ (.A(_05729_),
    .B_N(_05731_),
    .X(_05732_));
 sky130_fd_sc_hd__nand2_1 _13150_ (.A(_05728_),
    .B(_05732_),
    .Y(_05733_));
 sky130_fd_sc_hd__xor2_1 _13151_ (.A(_05699_),
    .B(_05733_),
    .X(_05734_));
 sky130_fd_sc_hd__xor2_1 _13152_ (.A(_05731_),
    .B(_05729_),
    .X(_05735_));
 sky130_fd_sc_hd__a31o_2 _13153_ (.A1(_02909_),
    .A2(_03029_),
    .A3(_04088_),
    .B1(_04087_),
    .X(_05736_));
 sky130_fd_sc_hd__nand2_1 _13154_ (.A(_02909_),
    .B(_03022_),
    .Y(_05737_));
 sky130_fd_sc_hd__and2b_1 _13155_ (.A_N(_05722_),
    .B(_05721_),
    .X(_05738_));
 sky130_fd_sc_hd__xnor2_2 _13156_ (.A(_05737_),
    .B(_05738_),
    .Y(_05739_));
 sky130_fd_sc_hd__o21a_1 _13157_ (.A1(_04073_),
    .A2(_04075_),
    .B1(_05739_),
    .X(_05740_));
 sky130_fd_sc_hd__nor3_1 _13158_ (.A(_04073_),
    .B(_04075_),
    .C(_05739_),
    .Y(_05741_));
 sky130_fd_sc_hd__nor2_1 _13159_ (.A(_05740_),
    .B(_05741_),
    .Y(_05742_));
 sky130_fd_sc_hd__a21oi_2 _13160_ (.A1(_05736_),
    .A2(_05742_),
    .B1(_05740_),
    .Y(_05743_));
 sky130_fd_sc_hd__o211ai_2 _13161_ (.A1(_03979_),
    .A2(_03992_),
    .B1(_04056_),
    .C1(_04057_),
    .Y(_05744_));
 sky130_fd_sc_hd__inv_2 _13162_ (.A(_05710_),
    .Y(_05745_));
 sky130_fd_sc_hd__a22oi_2 _13163_ (.A1(_05702_),
    .A2(_05703_),
    .B1(_05708_),
    .B2(_05709_),
    .Y(_05746_));
 sky130_fd_sc_hd__a211oi_2 _13164_ (.A1(_05744_),
    .A2(_04077_),
    .B1(_05745_),
    .C1(_05746_),
    .Y(_05747_));
 sky130_fd_sc_hd__o211a_1 _13165_ (.A1(_05745_),
    .A2(_05746_),
    .B1(_05744_),
    .C1(_04077_),
    .X(_05748_));
 sky130_fd_sc_hd__xnor2_1 _13166_ (.A(_05736_),
    .B(_05742_),
    .Y(_05749_));
 sky130_fd_sc_hd__nor3_1 _13167_ (.A(_05747_),
    .B(_05748_),
    .C(_05749_),
    .Y(_05750_));
 sky130_fd_sc_hd__xor2_2 _13168_ (.A(_05712_),
    .B(_05724_),
    .X(_05751_));
 sky130_fd_sc_hd__o21ai_1 _13169_ (.A1(_05747_),
    .A2(_05750_),
    .B1(_05751_),
    .Y(_05752_));
 sky130_fd_sc_hd__or3_1 _13170_ (.A(_05747_),
    .B(_05750_),
    .C(_05751_),
    .X(_05753_));
 sky130_fd_sc_hd__nand2_1 _13171_ (.A(_05752_),
    .B(_05753_),
    .Y(_05754_));
 sky130_fd_sc_hd__o21a_1 _13172_ (.A1(_05743_),
    .A2(_05754_),
    .B1(_05752_),
    .X(_05755_));
 sky130_fd_sc_hd__xnor2_1 _13173_ (.A(_05735_),
    .B(_05755_),
    .Y(_05756_));
 sky130_fd_sc_hd__or2_1 _13174_ (.A(_05734_),
    .B(_05756_),
    .X(_05757_));
 sky130_fd_sc_hd__or2b_1 _13175_ (.A(_04084_),
    .B_N(_04090_),
    .X(_05758_));
 sky130_fd_sc_hd__nand2_1 _13176_ (.A(_04082_),
    .B(_04091_),
    .Y(_05759_));
 sky130_fd_sc_hd__nor3_1 _13177_ (.A(_04079_),
    .B(_04080_),
    .C(_04092_),
    .Y(_05760_));
 sky130_fd_sc_hd__inv_2 _13178_ (.A(_05750_),
    .Y(_05761_));
 sky130_fd_sc_hd__o21ai_1 _13179_ (.A1(_05747_),
    .A2(_05748_),
    .B1(_05749_),
    .Y(_05762_));
 sky130_fd_sc_hd__o211a_1 _13180_ (.A1(_04079_),
    .A2(_05760_),
    .B1(_05761_),
    .C1(_05762_),
    .X(_05763_));
 sky130_fd_sc_hd__a211oi_2 _13181_ (.A1(_05761_),
    .A2(_05762_),
    .B1(_04079_),
    .C1(_05760_),
    .Y(_05764_));
 sky130_fd_sc_hd__a211oi_2 _13182_ (.A1(_05758_),
    .A2(_05759_),
    .B1(_05763_),
    .C1(_05764_),
    .Y(_05765_));
 sky130_fd_sc_hd__o211ai_1 _13183_ (.A1(_05763_),
    .A2(_05764_),
    .B1(_05758_),
    .C1(_05759_),
    .Y(_05766_));
 sky130_fd_sc_hd__or2b_1 _13184_ (.A(_05765_),
    .B_N(_05766_),
    .X(_05767_));
 sky130_fd_sc_hd__or2_1 _13185_ (.A(_04095_),
    .B(_04097_),
    .X(_05768_));
 sky130_fd_sc_hd__xor2_1 _13186_ (.A(_05767_),
    .B(_05768_),
    .X(_05769_));
 sky130_fd_sc_hd__xor2_2 _13187_ (.A(_05743_),
    .B(_05754_),
    .X(_05770_));
 sky130_fd_sc_hd__nor3_2 _13188_ (.A(_05763_),
    .B(_05765_),
    .C(_05770_),
    .Y(_05771_));
 sky130_fd_sc_hd__o21a_1 _13189_ (.A1(_05763_),
    .A2(_05765_),
    .B1(_05770_),
    .X(_05772_));
 sky130_fd_sc_hd__or3_1 _13190_ (.A(_05769_),
    .B(_05771_),
    .C(_05772_),
    .X(_05773_));
 sky130_fd_sc_hd__a211o_2 _13191_ (.A1(_05291_),
    .A2(_05698_),
    .B1(_05757_),
    .C1(_05773_),
    .X(_05774_));
 sky130_fd_sc_hd__and3_1 _13192_ (.A(_05699_),
    .B(_05728_),
    .C(_05732_),
    .X(_05775_));
 sky130_fd_sc_hd__or2_1 _13193_ (.A(_05735_),
    .B(_05755_),
    .X(_05776_));
 sky130_fd_sc_hd__and3b_1 _13194_ (.A_N(_05765_),
    .B(_05766_),
    .C(_05768_),
    .X(_05777_));
 sky130_fd_sc_hd__nor2_1 _13195_ (.A(_05777_),
    .B(_05772_),
    .Y(_05778_));
 sky130_fd_sc_hd__or2_1 _13196_ (.A(_05771_),
    .B(_05778_),
    .X(_05779_));
 sky130_fd_sc_hd__or2b_1 _13197_ (.A(_05699_),
    .B_N(_05733_),
    .X(_05780_));
 sky130_fd_sc_hd__o221a_2 _13198_ (.A1(_05775_),
    .A2(_05776_),
    .B1(_05757_),
    .B2(_05779_),
    .C1(_05780_),
    .X(_05781_));
 sky130_fd_sc_hd__and2b_1 _13199_ (.A_N(_03752_),
    .B(_03670_),
    .X(_05782_));
 sky130_fd_sc_hd__and3_1 _13200_ (.A(_03744_),
    .B(_03749_),
    .C(_03750_),
    .X(_05783_));
 sky130_fd_sc_hd__nor2_1 _13201_ (.A(_03751_),
    .B(_05783_),
    .Y(_05784_));
 sky130_fd_sc_hd__nand2_1 _13202_ (.A(_05782_),
    .B(_05784_),
    .Y(_05785_));
 sky130_fd_sc_hd__a211o_2 _13203_ (.A1(_05774_),
    .A2(_05781_),
    .B1(_05785_),
    .C1(_03591_),
    .X(_05786_));
 sky130_fd_sc_hd__nand2_1 _13204_ (.A(_03380_),
    .B(_03385_),
    .Y(_05787_));
 sky130_fd_sc_hd__or2b_1 _13205_ (.A(_03387_),
    .B_N(_03386_),
    .X(_05788_));
 sky130_fd_sc_hd__a21oi_1 _13206_ (.A1(_05787_),
    .A2(_05788_),
    .B1(_02932_),
    .Y(_05789_));
 sky130_fd_sc_hd__and3_1 _13207_ (.A(_02932_),
    .B(_05787_),
    .C(_05788_),
    .X(_05790_));
 sky130_fd_sc_hd__or2_1 _13208_ (.A(_05789_),
    .B(_05790_),
    .X(_05791_));
 sky130_fd_sc_hd__and2b_1 _13209_ (.A_N(_03409_),
    .B(_02916_),
    .X(_05792_));
 sky130_fd_sc_hd__or2_1 _13210_ (.A(_02925_),
    .B(_05792_),
    .X(_05793_));
 sky130_fd_sc_hd__and2b_1 _13211_ (.A_N(_05791_),
    .B(_05793_),
    .X(_05794_));
 sky130_fd_sc_hd__o21a_1 _13212_ (.A1(_05789_),
    .A2(_05794_),
    .B1(_02913_),
    .X(_05795_));
 sky130_fd_sc_hd__nor3_1 _13213_ (.A(_02913_),
    .B(_05789_),
    .C(_05794_),
    .Y(_05796_));
 sky130_fd_sc_hd__nor2_1 _13214_ (.A(_05795_),
    .B(_05796_),
    .Y(_05797_));
 sky130_fd_sc_hd__a21o_1 _13215_ (.A1(_02982_),
    .A2(_05797_),
    .B1(_05795_),
    .X(_05798_));
 sky130_fd_sc_hd__a31o_1 _13216_ (.A1(_02950_),
    .A2(_03040_),
    .A3(_03390_),
    .B1(_03389_),
    .X(_05799_));
 sky130_fd_sc_hd__and4_1 _13217_ (.A(_02969_),
    .B(_03302_),
    .C(_02952_),
    .D(_03022_),
    .X(_05800_));
 sky130_fd_sc_hd__a22oi_1 _13218_ (.A1(_03302_),
    .A2(_02952_),
    .B1(_03022_),
    .B2(_02969_),
    .Y(_05801_));
 sky130_fd_sc_hd__nor2_1 _13219_ (.A(_05800_),
    .B(_05801_),
    .Y(_05802_));
 sky130_fd_sc_hd__xnor2_1 _13220_ (.A(_02936_),
    .B(_05802_),
    .Y(_05803_));
 sky130_fd_sc_hd__xor2_1 _13221_ (.A(_05799_),
    .B(_05803_),
    .X(_05804_));
 sky130_fd_sc_hd__o21ba_1 _13222_ (.A1(_03381_),
    .A2(_03383_),
    .B1_N(_03382_),
    .X(_05805_));
 sky130_fd_sc_hd__xnor2_1 _13223_ (.A(_05804_),
    .B(_05805_),
    .Y(_05806_));
 sky130_fd_sc_hd__and4_1 _13224_ (.A(_02961_),
    .B(_02956_),
    .C(_03039_),
    .D(_03094_),
    .X(_05807_));
 sky130_fd_sc_hd__a22oi_2 _13225_ (.A1(_02956_),
    .A2(_03039_),
    .B1(_03094_),
    .B2(_02961_),
    .Y(_05808_));
 sky130_fd_sc_hd__nor2_1 _13226_ (.A(_05807_),
    .B(_05808_),
    .Y(_05809_));
 sky130_fd_sc_hd__nand2_1 _13227_ (.A(_03100_),
    .B(_03029_),
    .Y(_05810_));
 sky130_fd_sc_hd__xnor2_1 _13228_ (.A(_05809_),
    .B(_05810_),
    .Y(_05811_));
 sky130_fd_sc_hd__nand2_1 _13229_ (.A(_03021_),
    .B(_03394_),
    .Y(_05812_));
 sky130_fd_sc_hd__xor2_1 _13230_ (.A(_03130_),
    .B(_05812_),
    .X(_05813_));
 sky130_fd_sc_hd__xor2_1 _13231_ (.A(_05811_),
    .B(_05813_),
    .X(_05814_));
 sky130_fd_sc_hd__a2bb2o_1 _13232_ (.A1_N(_05812_),
    .A2_N(_03359_),
    .B1(_03396_),
    .B2(_03393_),
    .X(_05815_));
 sky130_fd_sc_hd__and2_1 _13233_ (.A(_05814_),
    .B(_05815_),
    .X(_05816_));
 sky130_fd_sc_hd__nor2_1 _13234_ (.A(_05814_),
    .B(_05815_),
    .Y(_05817_));
 sky130_fd_sc_hd__nor2_1 _13235_ (.A(_05816_),
    .B(_05817_),
    .Y(_05818_));
 sky130_fd_sc_hd__and2_1 _13236_ (.A(_05806_),
    .B(_05818_),
    .X(_05819_));
 sky130_fd_sc_hd__nor2_1 _13237_ (.A(_05806_),
    .B(_05818_),
    .Y(_05820_));
 sky130_fd_sc_hd__a211o_1 _13238_ (.A1(_03399_),
    .A2(_03402_),
    .B1(_05819_),
    .C1(_05820_),
    .X(_05821_));
 sky130_fd_sc_hd__xnor2_1 _13239_ (.A(_05791_),
    .B(_05793_),
    .Y(_05822_));
 sky130_fd_sc_hd__o211ai_1 _13240_ (.A1(_05819_),
    .A2(_05820_),
    .B1(_03399_),
    .C1(_03402_),
    .Y(_05823_));
 sky130_fd_sc_hd__and3_1 _13241_ (.A(_05822_),
    .B(_05821_),
    .C(_05823_),
    .X(_05824_));
 sky130_fd_sc_hd__inv_2 _13242_ (.A(_05824_),
    .Y(_05825_));
 sky130_fd_sc_hd__nand2_1 _13243_ (.A(_05799_),
    .B(_05803_),
    .Y(_05826_));
 sky130_fd_sc_hd__or2b_1 _13244_ (.A(_05805_),
    .B_N(_05804_),
    .X(_05827_));
 sky130_fd_sc_hd__a21o_1 _13245_ (.A1(_05826_),
    .A2(_05827_),
    .B1(_02932_),
    .X(_05828_));
 sky130_fd_sc_hd__nand3_1 _13246_ (.A(_02932_),
    .B(_05826_),
    .C(_05827_),
    .Y(_05829_));
 sky130_fd_sc_hd__nand2_1 _13247_ (.A(_05828_),
    .B(_05829_),
    .Y(_05830_));
 sky130_fd_sc_hd__xnor2_1 _13248_ (.A(_02975_),
    .B(_05830_),
    .Y(_05831_));
 sky130_fd_sc_hd__o21ba_1 _13249_ (.A1(_05808_),
    .A2(_05810_),
    .B1_N(_05807_),
    .X(_05832_));
 sky130_fd_sc_hd__and2b_1 _13250_ (.A_N(_03147_),
    .B(_03146_),
    .X(_05833_));
 sky130_fd_sc_hd__xnor2_1 _13251_ (.A(_02936_),
    .B(_05833_),
    .Y(_05834_));
 sky130_fd_sc_hd__xnor2_1 _13252_ (.A(_05832_),
    .B(_05834_),
    .Y(_05835_));
 sky130_fd_sc_hd__o21ba_1 _13253_ (.A1(_02936_),
    .A2(_05801_),
    .B1_N(_05800_),
    .X(_05836_));
 sky130_fd_sc_hd__xor2_1 _13254_ (.A(_05835_),
    .B(_05836_),
    .X(_05837_));
 sky130_fd_sc_hd__xnor2_1 _13255_ (.A(_03137_),
    .B(_03132_),
    .Y(_05838_));
 sky130_fd_sc_hd__a2bb2o_1 _13256_ (.A1_N(_03131_),
    .A2_N(_03394_),
    .B1(_05813_),
    .B2(_05811_),
    .X(_05839_));
 sky130_fd_sc_hd__xor2_1 _13257_ (.A(_05838_),
    .B(_05839_),
    .X(_05840_));
 sky130_fd_sc_hd__or2_1 _13258_ (.A(_05837_),
    .B(_05840_),
    .X(_05841_));
 sky130_fd_sc_hd__nand2_1 _13259_ (.A(_05837_),
    .B(_05840_),
    .Y(_05842_));
 sky130_fd_sc_hd__o211a_1 _13260_ (.A1(_05816_),
    .A2(_05819_),
    .B1(_05841_),
    .C1(_05842_),
    .X(_05843_));
 sky130_fd_sc_hd__a211oi_1 _13261_ (.A1(_05841_),
    .A2(_05842_),
    .B1(_05816_),
    .C1(_05819_),
    .Y(_05844_));
 sky130_fd_sc_hd__or3_1 _13262_ (.A(_05831_),
    .B(_05843_),
    .C(_05844_),
    .X(_05845_));
 sky130_fd_sc_hd__o21ai_1 _13263_ (.A1(_05843_),
    .A2(_05844_),
    .B1(_05831_),
    .Y(_05846_));
 sky130_fd_sc_hd__nand2_1 _13264_ (.A(_05845_),
    .B(_05846_),
    .Y(_05847_));
 sky130_fd_sc_hd__a21oi_4 _13265_ (.A1(_05821_),
    .A2(_05825_),
    .B1(_05847_),
    .Y(_05848_));
 sky130_fd_sc_hd__xnor2_1 _13266_ (.A(_02981_),
    .B(_05797_),
    .Y(_05849_));
 sky130_fd_sc_hd__and3_1 _13267_ (.A(_05821_),
    .B(_05825_),
    .C(_05847_),
    .X(_05850_));
 sky130_fd_sc_hd__nor3_4 _13268_ (.A(_05849_),
    .B(_05848_),
    .C(_05850_),
    .Y(_05851_));
 sky130_fd_sc_hd__o21ai_1 _13269_ (.A1(_02975_),
    .A2(_05830_),
    .B1(_05828_),
    .Y(_05852_));
 sky130_fd_sc_hd__xor2_1 _13270_ (.A(_02913_),
    .B(_05852_),
    .X(_05853_));
 sky130_fd_sc_hd__nand2_1 _13271_ (.A(_02981_),
    .B(_05853_),
    .Y(_05854_));
 sky130_fd_sc_hd__or2_1 _13272_ (.A(_02981_),
    .B(_05853_),
    .X(_05855_));
 sky130_fd_sc_hd__nand2_1 _13273_ (.A(_05854_),
    .B(_05855_),
    .Y(_05856_));
 sky130_fd_sc_hd__inv_2 _13274_ (.A(_05843_),
    .Y(_05857_));
 sky130_fd_sc_hd__or2b_1 _13275_ (.A(_05832_),
    .B_N(_05834_),
    .X(_05858_));
 sky130_fd_sc_hd__or2b_1 _13276_ (.A(_05836_),
    .B_N(_05835_),
    .X(_05859_));
 sky130_fd_sc_hd__a21o_1 _13277_ (.A1(_05858_),
    .A2(_05859_),
    .B1(_02932_),
    .X(_05860_));
 sky130_fd_sc_hd__nand3_1 _13278_ (.A(_02932_),
    .B(_05858_),
    .C(_05859_),
    .Y(_05861_));
 sky130_fd_sc_hd__nand2_1 _13279_ (.A(_05860_),
    .B(_05861_),
    .Y(_05862_));
 sky130_fd_sc_hd__xnor2_1 _13280_ (.A(_02975_),
    .B(_05862_),
    .Y(_05863_));
 sky130_fd_sc_hd__or2b_1 _13281_ (.A(_05838_),
    .B_N(_05839_),
    .X(_05864_));
 sky130_fd_sc_hd__xnor2_1 _13282_ (.A(_03149_),
    .B(_03150_),
    .Y(_05865_));
 sky130_fd_sc_hd__a21oi_1 _13283_ (.A1(_05864_),
    .A2(_05841_),
    .B1(_05865_),
    .Y(_05866_));
 sky130_fd_sc_hd__and3_1 _13284_ (.A(_05864_),
    .B(_05841_),
    .C(_05865_),
    .X(_05867_));
 sky130_fd_sc_hd__or2_1 _13285_ (.A(_05866_),
    .B(_05867_),
    .X(_05868_));
 sky130_fd_sc_hd__nor2_1 _13286_ (.A(_05863_),
    .B(_05868_),
    .Y(_05869_));
 sky130_fd_sc_hd__and2_1 _13287_ (.A(_05863_),
    .B(_05868_),
    .X(_05870_));
 sky130_fd_sc_hd__or2_1 _13288_ (.A(_05869_),
    .B(_05870_),
    .X(_05871_));
 sky130_fd_sc_hd__a21oi_1 _13289_ (.A1(_05857_),
    .A2(_05845_),
    .B1(_05871_),
    .Y(_05872_));
 sky130_fd_sc_hd__and3_1 _13290_ (.A(_05857_),
    .B(_05845_),
    .C(_05871_),
    .X(_05873_));
 sky130_fd_sc_hd__or3_2 _13291_ (.A(_05856_),
    .B(_05872_),
    .C(_05873_),
    .X(_05874_));
 sky130_fd_sc_hd__o21ai_2 _13292_ (.A1(_05872_),
    .A2(_05873_),
    .B1(_05856_),
    .Y(_05875_));
 sky130_fd_sc_hd__o211ai_4 _13293_ (.A1(_05848_),
    .A2(_05851_),
    .B1(_05874_),
    .C1(_05875_),
    .Y(_05876_));
 sky130_fd_sc_hd__a211o_1 _13294_ (.A1(_05874_),
    .A2(_05875_),
    .B1(_05848_),
    .C1(_05851_),
    .X(_05877_));
 sky130_fd_sc_hd__nand3_1 _13295_ (.A(_05798_),
    .B(_05876_),
    .C(_05877_),
    .Y(_05878_));
 sky130_fd_sc_hd__a21o_1 _13296_ (.A1(_05876_),
    .A2(_05877_),
    .B1(_05798_),
    .X(_05879_));
 sky130_fd_sc_hd__nand2_1 _13297_ (.A(_05878_),
    .B(_05879_),
    .Y(_05880_));
 sky130_fd_sc_hd__a21oi_1 _13298_ (.A1(_05821_),
    .A2(_05823_),
    .B1(_05822_),
    .Y(_05881_));
 sky130_fd_sc_hd__a211o_1 _13299_ (.A1(_03404_),
    .A2(_03418_),
    .B1(_05824_),
    .C1(_05881_),
    .X(_05882_));
 sky130_fd_sc_hd__or2b_1 _13300_ (.A(_03415_),
    .B_N(_03413_),
    .X(_05883_));
 sky130_fd_sc_hd__nand2_1 _13301_ (.A(_03411_),
    .B(_05883_),
    .Y(_05884_));
 sky130_fd_sc_hd__xor2_1 _13302_ (.A(_02913_),
    .B(_05884_),
    .X(_05885_));
 sky130_fd_sc_hd__xor2_1 _13303_ (.A(_02981_),
    .B(_05885_),
    .X(_05886_));
 sky130_fd_sc_hd__o211ai_2 _13304_ (.A1(_05824_),
    .A2(_05881_),
    .B1(_03404_),
    .C1(_03418_),
    .Y(_05887_));
 sky130_fd_sc_hd__nand3_2 _13305_ (.A(_05886_),
    .B(_05882_),
    .C(_05887_),
    .Y(_05888_));
 sky130_fd_sc_hd__o21a_1 _13306_ (.A1(_05848_),
    .A2(_05850_),
    .B1(_05849_),
    .X(_05889_));
 sky130_fd_sc_hd__a211oi_2 _13307_ (.A1(_05882_),
    .A2(_05888_),
    .B1(_05851_),
    .C1(_05889_),
    .Y(_05890_));
 sky130_fd_sc_hd__nand2_1 _13308_ (.A(_02914_),
    .B(_05884_),
    .Y(_05891_));
 sky130_fd_sc_hd__nand2_1 _13309_ (.A(_02982_),
    .B(_05885_),
    .Y(_05892_));
 sky130_fd_sc_hd__o211a_1 _13310_ (.A1(_05851_),
    .A2(_05889_),
    .B1(_05882_),
    .C1(_05888_),
    .X(_05893_));
 sky130_fd_sc_hd__a211oi_2 _13311_ (.A1(_05891_),
    .A2(_05892_),
    .B1(_05890_),
    .C1(_05893_),
    .Y(_05894_));
 sky130_fd_sc_hd__nor2_1 _13312_ (.A(_05890_),
    .B(_05894_),
    .Y(_05895_));
 sky130_fd_sc_hd__or2_1 _13313_ (.A(_05880_),
    .B(_05895_),
    .X(_05896_));
 sky130_fd_sc_hd__nand2_1 _13314_ (.A(_05880_),
    .B(_05895_),
    .Y(_05897_));
 sky130_fd_sc_hd__nand2_1 _13315_ (.A(_05896_),
    .B(_05897_),
    .Y(_05898_));
 sky130_fd_sc_hd__nand2_1 _13316_ (.A(_02914_),
    .B(_05852_),
    .Y(_05899_));
 sky130_fd_sc_hd__o21ai_1 _13317_ (.A1(_02976_),
    .A2(_05862_),
    .B1(_05860_),
    .Y(_05900_));
 sky130_fd_sc_hd__xor2_1 _13318_ (.A(_02913_),
    .B(_05900_),
    .X(_05901_));
 sky130_fd_sc_hd__nand2_1 _13319_ (.A(_02981_),
    .B(_05901_),
    .Y(_05902_));
 sky130_fd_sc_hd__or2_1 _13320_ (.A(_02981_),
    .B(_05901_),
    .X(_05903_));
 sky130_fd_sc_hd__nand2_1 _13321_ (.A(_05902_),
    .B(_05903_),
    .Y(_05904_));
 sky130_fd_sc_hd__o21ai_1 _13322_ (.A1(_03154_),
    .A2(_03162_),
    .B1(_03161_),
    .Y(_05905_));
 sky130_fd_sc_hd__o211a_1 _13323_ (.A1(_05866_),
    .A2(_05869_),
    .B1(_05905_),
    .C1(_03163_),
    .X(_05906_));
 sky130_fd_sc_hd__a211oi_1 _13324_ (.A1(_03163_),
    .A2(_05905_),
    .B1(_05869_),
    .C1(_05866_),
    .Y(_05907_));
 sky130_fd_sc_hd__nor3_1 _13325_ (.A(_05904_),
    .B(_05906_),
    .C(_05907_),
    .Y(_05908_));
 sky130_fd_sc_hd__o21a_1 _13326_ (.A1(_05906_),
    .A2(_05907_),
    .B1(_05904_),
    .X(_05909_));
 sky130_fd_sc_hd__or2_1 _13327_ (.A(_05908_),
    .B(_05909_),
    .X(_05910_));
 sky130_fd_sc_hd__and2b_1 _13328_ (.A_N(_05872_),
    .B(_05874_),
    .X(_05911_));
 sky130_fd_sc_hd__nor2_1 _13329_ (.A(_05910_),
    .B(_05911_),
    .Y(_05912_));
 sky130_fd_sc_hd__and2_1 _13330_ (.A(_05910_),
    .B(_05911_),
    .X(_05913_));
 sky130_fd_sc_hd__a211oi_2 _13331_ (.A1(_05899_),
    .A2(_05854_),
    .B1(_05912_),
    .C1(_05913_),
    .Y(_05914_));
 sky130_fd_sc_hd__o211a_1 _13332_ (.A1(_05912_),
    .A2(_05913_),
    .B1(_05899_),
    .C1(_05854_),
    .X(_05915_));
 sky130_fd_sc_hd__a211o_1 _13333_ (.A1(_05876_),
    .A2(_05878_),
    .B1(_05914_),
    .C1(_05915_),
    .X(_05916_));
 sky130_fd_sc_hd__o211ai_1 _13334_ (.A1(_05914_),
    .A2(_05915_),
    .B1(_05876_),
    .C1(_05878_),
    .Y(_05917_));
 sky130_fd_sc_hd__nand2_1 _13335_ (.A(_05916_),
    .B(_05917_),
    .Y(_05918_));
 sky130_fd_sc_hd__or2_1 _13336_ (.A(_05898_),
    .B(_05918_),
    .X(_05919_));
 sky130_fd_sc_hd__a21o_1 _13337_ (.A1(_02982_),
    .A2(_03424_),
    .B1(_03422_),
    .X(_05920_));
 sky130_fd_sc_hd__a21o_1 _13338_ (.A1(_05882_),
    .A2(_05887_),
    .B1(_05886_),
    .X(_05921_));
 sky130_fd_sc_hd__o211ai_2 _13339_ (.A1(_03421_),
    .A2(_03427_),
    .B1(_05888_),
    .C1(_05921_),
    .Y(_05922_));
 sky130_fd_sc_hd__a211o_1 _13340_ (.A1(_05888_),
    .A2(_05921_),
    .B1(_03421_),
    .C1(_03427_),
    .X(_05923_));
 sky130_fd_sc_hd__nand3_1 _13341_ (.A(_05920_),
    .B(_05922_),
    .C(_05923_),
    .Y(_05924_));
 sky130_fd_sc_hd__a21o_1 _13342_ (.A1(_05922_),
    .A2(_05923_),
    .B1(_05920_),
    .X(_05925_));
 sky130_fd_sc_hd__and2_1 _13343_ (.A(_05924_),
    .B(_05925_),
    .X(_05926_));
 sky130_fd_sc_hd__o21ai_2 _13344_ (.A1(_03429_),
    .A2(_03431_),
    .B1(_05926_),
    .Y(_05927_));
 sky130_fd_sc_hd__or3_1 _13345_ (.A(_05926_),
    .B(_03429_),
    .C(_03431_),
    .X(_05928_));
 sky130_fd_sc_hd__and2_1 _13346_ (.A(_05927_),
    .B(_05928_),
    .X(_05929_));
 sky130_fd_sc_hd__o211a_1 _13347_ (.A1(_05890_),
    .A2(_05893_),
    .B1(_05891_),
    .C1(_05892_),
    .X(_05930_));
 sky130_fd_sc_hd__o211a_1 _13348_ (.A1(_05894_),
    .A2(_05930_),
    .B1(_05922_),
    .C1(_05924_),
    .X(_05931_));
 sky130_fd_sc_hd__a211o_1 _13349_ (.A1(_05922_),
    .A2(_05924_),
    .B1(_05894_),
    .C1(_05930_),
    .X(_05932_));
 sky130_fd_sc_hd__or2b_1 _13350_ (.A(_05931_),
    .B_N(_05932_),
    .X(_05933_));
 sky130_fd_sc_hd__inv_2 _13351_ (.A(_05933_),
    .Y(_05934_));
 sky130_fd_sc_hd__nand2_1 _13352_ (.A(_05929_),
    .B(_05934_),
    .Y(_05935_));
 sky130_fd_sc_hd__a211o_1 _13353_ (.A1(_03755_),
    .A2(_05786_),
    .B1(_05919_),
    .C1(_05935_),
    .X(_05936_));
 sky130_fd_sc_hd__o211a_1 _13354_ (.A1(_05914_),
    .A2(_05915_),
    .B1(_05876_),
    .C1(_05878_),
    .X(_05937_));
 sky130_fd_sc_hd__a21o_1 _13355_ (.A1(_05927_),
    .A2(_05932_),
    .B1(_05931_),
    .X(_05938_));
 sky130_fd_sc_hd__o221a_1 _13356_ (.A1(_05896_),
    .A2(_05937_),
    .B1(_05919_),
    .B2(_05938_),
    .C1(_05916_),
    .X(_05939_));
 sky130_fd_sc_hd__a21bo_1 _13357_ (.A1(_02914_),
    .A2(_05900_),
    .B1_N(_05902_),
    .X(_05940_));
 sky130_fd_sc_hd__o21ai_1 _13358_ (.A1(_03165_),
    .A2(_03171_),
    .B1(_03170_),
    .Y(_05941_));
 sky130_fd_sc_hd__o211a_1 _13359_ (.A1(_05906_),
    .A2(_05908_),
    .B1(_05941_),
    .C1(_03172_),
    .X(_05942_));
 sky130_fd_sc_hd__a211oi_1 _13360_ (.A1(_03172_),
    .A2(_05941_),
    .B1(_05908_),
    .C1(_05906_),
    .Y(_05943_));
 sky130_fd_sc_hd__nor2_1 _13361_ (.A(_05942_),
    .B(_05943_),
    .Y(_05944_));
 sky130_fd_sc_hd__xnor2_1 _13362_ (.A(_05940_),
    .B(_05944_),
    .Y(_05945_));
 sky130_fd_sc_hd__or2_1 _13363_ (.A(_05912_),
    .B(_05914_),
    .X(_05946_));
 sky130_fd_sc_hd__xnor2_1 _13364_ (.A(_05945_),
    .B(_05946_),
    .Y(_05947_));
 sky130_fd_sc_hd__inv_2 _13365_ (.A(_05947_),
    .Y(_05948_));
 sky130_fd_sc_hd__and2_1 _13366_ (.A(_05940_),
    .B(_05944_),
    .X(_05949_));
 sky130_fd_sc_hd__xnor2_1 _13367_ (.A(_03175_),
    .B(_03174_),
    .Y(_05950_));
 sky130_fd_sc_hd__o21a_1 _13368_ (.A1(_05942_),
    .A2(_05949_),
    .B1(_05950_),
    .X(_05951_));
 sky130_fd_sc_hd__or3_1 _13369_ (.A(_05942_),
    .B(_05949_),
    .C(_05950_),
    .X(_05952_));
 sky130_fd_sc_hd__and2b_1 _13370_ (.A_N(_05951_),
    .B(_05952_),
    .X(_05953_));
 sky130_fd_sc_hd__inv_2 _13371_ (.A(_05953_),
    .Y(_05954_));
 sky130_fd_sc_hd__a211o_1 _13372_ (.A1(_05936_),
    .A2(_05939_),
    .B1(_05948_),
    .C1(_05954_),
    .X(_05955_));
 sky130_fd_sc_hd__and2b_1 _13373_ (.A_N(_05945_),
    .B(_05946_),
    .X(_05956_));
 sky130_fd_sc_hd__o21ai_1 _13374_ (.A1(_05956_),
    .A2(_05951_),
    .B1(_05952_),
    .Y(_05957_));
 sky130_fd_sc_hd__o22a_1 _13375_ (.A1(_03203_),
    .A2(_03204_),
    .B1(_03207_),
    .B2(_05957_),
    .X(_05958_));
 sky130_fd_sc_hd__o21ai_2 _13376_ (.A1(_03207_),
    .A2(_05955_),
    .B1(_05958_),
    .Y(_05959_));
 sky130_fd_sc_hd__a21o_1 _13377_ (.A1(_03179_),
    .A2(_03202_),
    .B1(_03200_),
    .X(_05960_));
 sky130_fd_sc_hd__inv_2 _13378_ (.A(_03197_),
    .Y(_05961_));
 sky130_fd_sc_hd__a21o_1 _13379_ (.A1(_03191_),
    .A2(_05961_),
    .B1(_03189_),
    .X(_05962_));
 sky130_fd_sc_hd__or2_1 _13380_ (.A(_02933_),
    .B(_03181_),
    .X(_05963_));
 sky130_fd_sc_hd__o21a_1 _13381_ (.A1(_02976_),
    .A2(_03182_),
    .B1(_05963_),
    .X(_05964_));
 sky130_fd_sc_hd__inv_2 _13382_ (.A(_03194_),
    .Y(_05965_));
 sky130_fd_sc_hd__o21a_1 _13383_ (.A1(_02982_),
    .A2(_05965_),
    .B1(_03195_),
    .X(_05966_));
 sky130_fd_sc_hd__xnor2_1 _13384_ (.A(_05964_),
    .B(_05966_),
    .Y(_05967_));
 sky130_fd_sc_hd__o21ai_1 _13385_ (.A1(_03183_),
    .A2(_03187_),
    .B1(_03185_),
    .Y(_05968_));
 sky130_fd_sc_hd__or3b_1 _13386_ (.A(_03074_),
    .B(_03067_),
    .C_N(_03068_),
    .X(_05969_));
 sky130_fd_sc_hd__mux2_1 _13387_ (.A0(_03185_),
    .A1(_05969_),
    .S(_03183_),
    .X(_05970_));
 sky130_fd_sc_hd__nand2_1 _13388_ (.A(_05968_),
    .B(_05970_),
    .Y(_05971_));
 sky130_fd_sc_hd__xnor2_1 _13389_ (.A(_05967_),
    .B(_05971_),
    .Y(_05972_));
 sky130_fd_sc_hd__xnor2_2 _13390_ (.A(_05962_),
    .B(_05972_),
    .Y(_05973_));
 sky130_fd_sc_hd__xnor2_4 _13391_ (.A(_05960_),
    .B(_05973_),
    .Y(_05974_));
 sky130_fd_sc_hd__and2_1 _13392_ (.A(\wfg_stim_mem_top.ctrl_en_q ),
    .B(\wfg_stim_mem_top.wfg_stim_mem.cur_state[0] ),
    .X(_05975_));
 sky130_fd_sc_hd__clkbuf_2 _13393_ (.A(_05975_),
    .X(_00000_));
 sky130_fd_sc_hd__or3b_2 _13394_ (.A(\wfg_interconnect_top.driver1_select_q[1] ),
    .B(\wfg_drive_pat_top.wfg_axis_tready_o ),
    .C_N(\wfg_interconnect_top.driver1_select_q[0] ),
    .X(_05976_));
 sky130_fd_sc_hd__and2b_1 _13395_ (.A_N(\wfg_interconnect_top.driver1_select_q[1] ),
    .B(\wfg_interconnect_top.driver1_select_q[0] ),
    .X(_05977_));
 sky130_fd_sc_hd__mux2_1 _13396_ (.A0(_05977_),
    .A1(\wfg_drive_spi_top.wfg_axis_tready_o ),
    .S(_02798_),
    .X(_05978_));
 sky130_fd_sc_hd__nand2_1 _13397_ (.A(_05976_),
    .B(_05978_),
    .Y(_05979_));
 sky130_fd_sc_hd__a21o_1 _13398_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.cur_state[3] ),
    .A2(_05979_),
    .B1(\wfg_stim_mem_top.wfg_stim_mem.cur_state[1] ),
    .X(_00002_));
 sky130_fd_sc_hd__or3b_4 _13399_ (.A(_00000_),
    .B(_00002_),
    .C_N(\wfg_stim_mem_top.wfg_stim_mem.cur_state[2] ),
    .X(_05980_));
 sky130_fd_sc_hd__buf_2 _13400_ (.A(_05980_),
    .X(_05981_));
 sky130_fd_sc_hd__inv_2 _13401_ (.A(_05981_),
    .Y(_05982_));
 sky130_fd_sc_hd__o21ai_1 _13402_ (.A1(_05959_),
    .A2(_05974_),
    .B1(_05982_),
    .Y(_05983_));
 sky130_fd_sc_hd__a21oi_4 _13403_ (.A1(_05959_),
    .A2(_05974_),
    .B1(_05983_),
    .Y(_05984_));
 sky130_fd_sc_hd__buf_2 _13404_ (.A(_05984_),
    .X(_05985_));
 sky130_fd_sc_hd__a21o_1 _13405_ (.A1(_05936_),
    .A2(_05939_),
    .B1(_05948_),
    .X(_05986_));
 sky130_fd_sc_hd__or3b_1 _13406_ (.A(_05956_),
    .B(_05953_),
    .C_N(_05986_),
    .X(_05987_));
 sky130_fd_sc_hd__inv_2 _13407_ (.A(_05956_),
    .Y(_05988_));
 sky130_fd_sc_hd__a21o_1 _13408_ (.A1(_05988_),
    .A2(_05986_),
    .B1(_05954_),
    .X(_05989_));
 sky130_fd_sc_hd__a21bo_1 _13409_ (.A1(_03755_),
    .A2(_05786_),
    .B1_N(_05929_),
    .X(_05990_));
 sky130_fd_sc_hd__nand2_1 _13410_ (.A(_05927_),
    .B(_05990_),
    .Y(_05991_));
 sky130_fd_sc_hd__xnor2_1 _13411_ (.A(_05933_),
    .B(_05991_),
    .Y(_05992_));
 sky130_fd_sc_hd__a21o_1 _13412_ (.A1(_05774_),
    .A2(_05781_),
    .B1(_05785_),
    .X(_05993_));
 sky130_fd_sc_hd__a21oi_1 _13413_ (.A1(_05993_),
    .A2(_03753_),
    .B1(_03590_),
    .Y(_05994_));
 sky130_fd_sc_hd__nor2_1 _13414_ (.A(_03588_),
    .B(_03507_),
    .Y(_05995_));
 sky130_fd_sc_hd__o21a_1 _13415_ (.A1(_03586_),
    .A2(_05994_),
    .B1(_05995_),
    .X(_05996_));
 sky130_fd_sc_hd__nor3_1 _13416_ (.A(_03586_),
    .B(_05995_),
    .C(_05994_),
    .Y(_05997_));
 sky130_fd_sc_hd__nand2_1 _13417_ (.A(_03755_),
    .B(_05786_),
    .Y(_05998_));
 sky130_fd_sc_hd__xnor2_1 _13418_ (.A(_05929_),
    .B(_05998_),
    .Y(_05999_));
 sky130_fd_sc_hd__a21o_1 _13419_ (.A1(_05291_),
    .A2(_05698_),
    .B1(_05769_),
    .X(_06000_));
 sky130_fd_sc_hd__a211o_1 _13420_ (.A1(_06000_),
    .A2(_05778_),
    .B1(_05756_),
    .C1(_05771_),
    .X(_06001_));
 sky130_fd_sc_hd__and3_1 _13421_ (.A(_05734_),
    .B(_05776_),
    .C(_06001_),
    .X(_06002_));
 sky130_fd_sc_hd__a21oi_2 _13422_ (.A1(_05776_),
    .A2(_06001_),
    .B1(_05734_),
    .Y(_06003_));
 sky130_fd_sc_hd__and3_1 _13423_ (.A(_05993_),
    .B(_03753_),
    .C(_03590_),
    .X(_06004_));
 sky130_fd_sc_hd__o22a_1 _13424_ (.A1(_06002_),
    .A2(_06003_),
    .B1(_05994_),
    .B2(_06004_),
    .X(_06005_));
 sky130_fd_sc_hd__a21boi_1 _13425_ (.A1(_05774_),
    .A2(_05781_),
    .B1_N(_05784_),
    .Y(_06006_));
 sky130_fd_sc_hd__o21bai_1 _13426_ (.A1(_03751_),
    .A2(_06006_),
    .B1_N(_05782_),
    .Y(_06007_));
 sky130_fd_sc_hd__and2b_1 _13427_ (.A_N(_03751_),
    .B(_05782_),
    .X(_06008_));
 sky130_fd_sc_hd__nor2_1 _13428_ (.A(_05784_),
    .B(_06008_),
    .Y(_06009_));
 sky130_fd_sc_hd__a31o_1 _13429_ (.A1(_05774_),
    .A2(_05781_),
    .A3(_06009_),
    .B1(_06006_),
    .X(_06010_));
 sky130_fd_sc_hd__o211ai_1 _13430_ (.A1(_06000_),
    .A2(_05771_),
    .B1(_05756_),
    .C1(_05779_),
    .Y(_06011_));
 sky130_fd_sc_hd__nand2_1 _13431_ (.A(_06001_),
    .B(_06011_),
    .Y(_06012_));
 sky130_fd_sc_hd__inv_2 _13432_ (.A(_05777_),
    .Y(_06013_));
 sky130_fd_sc_hd__nor2_1 _13433_ (.A(_05771_),
    .B(_05772_),
    .Y(_06014_));
 sky130_fd_sc_hd__a21oi_1 _13434_ (.A1(_06013_),
    .A2(_06000_),
    .B1(_06014_),
    .Y(_06015_));
 sky130_fd_sc_hd__nand2_1 _13435_ (.A(_05291_),
    .B(_05698_),
    .Y(_06016_));
 sky130_fd_sc_hd__a21bo_1 _13436_ (.A1(_06013_),
    .A2(_06014_),
    .B1_N(_05769_),
    .X(_06017_));
 sky130_fd_sc_hd__o21a_1 _13437_ (.A1(_06016_),
    .A2(_06017_),
    .B1(_06000_),
    .X(_06018_));
 sky130_fd_sc_hd__nor2_1 _13438_ (.A(_06015_),
    .B(_06018_),
    .Y(_06019_));
 sky130_fd_sc_hd__and4_1 _13439_ (.A(_06007_),
    .B(_06010_),
    .C(_06012_),
    .D(_06019_),
    .X(_06020_));
 sky130_fd_sc_hd__o2111ai_4 _13440_ (.A1(_05996_),
    .A2(_05997_),
    .B1(_05999_),
    .C1(_06005_),
    .D1(_06020_),
    .Y(_06021_));
 sky130_fd_sc_hd__a311o_1 _13441_ (.A1(_05927_),
    .A2(_05990_),
    .A3(_05932_),
    .B1(_05898_),
    .C1(_05931_),
    .X(_06022_));
 sky130_fd_sc_hd__o211ai_1 _13442_ (.A1(_05990_),
    .A2(_05933_),
    .B1(_05898_),
    .C1(_05938_),
    .Y(_06023_));
 sky130_fd_sc_hd__nand3_1 _13443_ (.A(_05936_),
    .B(_05939_),
    .C(_05948_),
    .Y(_06024_));
 sky130_fd_sc_hd__a22o_1 _13444_ (.A1(_06022_),
    .A2(_06023_),
    .B1(_05986_),
    .B2(_06024_),
    .X(_06025_));
 sky130_fd_sc_hd__a2111o_1 _13445_ (.A1(_05987_),
    .A2(_05989_),
    .B1(_05992_),
    .C1(_06021_),
    .D1(_06025_),
    .X(_06026_));
 sky130_fd_sc_hd__or2_1 _13446_ (.A(_03123_),
    .B(_03177_),
    .X(_06027_));
 sky130_fd_sc_hd__a21o_1 _13447_ (.A1(_05955_),
    .A2(_05957_),
    .B1(_03178_),
    .X(_06028_));
 sky130_fd_sc_hd__and3_1 _13448_ (.A(_06027_),
    .B(_03205_),
    .C(_06028_),
    .X(_06029_));
 sky130_fd_sc_hd__a21o_1 _13449_ (.A1(_06027_),
    .A2(_06028_),
    .B1(_03205_),
    .X(_06030_));
 sky130_fd_sc_hd__nand3_1 _13450_ (.A(_03178_),
    .B(_05955_),
    .C(_05957_),
    .Y(_06031_));
 sky130_fd_sc_hd__and3_1 _13451_ (.A(_05896_),
    .B(_05918_),
    .C(_06022_),
    .X(_06032_));
 sky130_fd_sc_hd__a21oi_1 _13452_ (.A1(_05896_),
    .A2(_06022_),
    .B1(_05918_),
    .Y(_06033_));
 sky130_fd_sc_hd__o2bb2a_1 _13453_ (.A1_N(_06028_),
    .A2_N(_06031_),
    .B1(_06032_),
    .B2(_06033_),
    .X(_06034_));
 sky130_fd_sc_hd__and4bb_2 _13454_ (.A_N(_06026_),
    .B_N(_06029_),
    .C(_06030_),
    .D(_06034_),
    .X(_06035_));
 sky130_fd_sc_hd__buf_2 _13455_ (.A(_06035_),
    .X(_06036_));
 sky130_fd_sc_hd__a21oi_4 _13456_ (.A1(_05666_),
    .A2(_05685_),
    .B1(_05697_),
    .Y(_06037_));
 sky130_fd_sc_hd__or2b_1 _13457_ (.A(_05692_),
    .B_N(_06037_),
    .X(_06038_));
 sky130_fd_sc_hd__o21ai_2 _13458_ (.A1(_05686_),
    .A2(_06038_),
    .B1(_05280_),
    .Y(_06039_));
 sky130_fd_sc_hd__or2b_1 _13459_ (.A(_04677_),
    .B_N(_06039_),
    .X(_06040_));
 sky130_fd_sc_hd__a21oi_4 _13460_ (.A1(_05285_),
    .A2(_06040_),
    .B1(_04345_),
    .Y(_06041_));
 sky130_fd_sc_hd__o31a_2 _13461_ (.A1(_04262_),
    .A2(_05287_),
    .A3(_06041_),
    .B1(_04261_),
    .X(_06042_));
 sky130_fd_sc_hd__a21oi_2 _13462_ (.A1(_04182_),
    .A2(_06042_),
    .B1(_04180_),
    .Y(_06043_));
 sky130_fd_sc_hd__xnor2_4 _13463_ (.A(_04101_),
    .B(_06043_),
    .Y(_06044_));
 sky130_fd_sc_hd__nand2_1 _13464_ (.A(_06036_),
    .B(_06044_),
    .Y(_06045_));
 sky130_fd_sc_hd__o2bb2a_1 _13465_ (.A1_N(_05985_),
    .A2_N(_06045_),
    .B1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[31] ),
    .B2(_05982_),
    .X(_01133_));
 sky130_fd_sc_hd__buf_2 _13466_ (.A(_05981_),
    .X(_06046_));
 sky130_fd_sc_hd__xnor2_4 _13467_ (.A(_04182_),
    .B(_06042_),
    .Y(_06047_));
 sky130_fd_sc_hd__nand2_1 _13468_ (.A(_06036_),
    .B(_06047_),
    .Y(_06048_));
 sky130_fd_sc_hd__a22o_1 _13469_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[30] ),
    .A2(_06046_),
    .B1(_05985_),
    .B2(_06048_),
    .X(_01132_));
 sky130_fd_sc_hd__nor2_2 _13470_ (.A(_05287_),
    .B(_06041_),
    .Y(_06049_));
 sky130_fd_sc_hd__xnor2_4 _13471_ (.A(_04264_),
    .B(_06049_),
    .Y(_06050_));
 sky130_fd_sc_hd__nand2_1 _13472_ (.A(_06036_),
    .B(_06050_),
    .Y(_06051_));
 sky130_fd_sc_hd__a22o_1 _13473_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[29] ),
    .A2(_06046_),
    .B1(_05985_),
    .B2(_06051_),
    .X(_01131_));
 sky130_fd_sc_hd__and3_2 _13474_ (.A(_04345_),
    .B(_05285_),
    .C(_06040_),
    .X(_06052_));
 sky130_fd_sc_hd__clkbuf_4 _13475_ (.A(_06035_),
    .X(_06053_));
 sky130_fd_sc_hd__o21ai_1 _13476_ (.A1(_06041_),
    .A2(_06052_),
    .B1(_06053_),
    .Y(_06054_));
 sky130_fd_sc_hd__a22o_1 _13477_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[28] ),
    .A2(_06046_),
    .B1(_05985_),
    .B2(_06054_),
    .X(_01130_));
 sky130_fd_sc_hd__and2_4 _13478_ (.A(_04676_),
    .B(_06039_),
    .X(_06055_));
 sky130_fd_sc_hd__o2bb2a_2 _13479_ (.A1_N(_04597_),
    .A2_N(_06055_),
    .B1(_05283_),
    .B2(_05281_),
    .X(_06056_));
 sky130_fd_sc_hd__o21ba_1 _13480_ (.A1(_04509_),
    .A2(_06056_),
    .B1_N(_04507_),
    .X(_06057_));
 sky130_fd_sc_hd__xnor2_4 _13481_ (.A(_04425_),
    .B(_06057_),
    .Y(_06058_));
 sky130_fd_sc_hd__nand2_1 _13482_ (.A(_06036_),
    .B(_06058_),
    .Y(_06059_));
 sky130_fd_sc_hd__a22o_1 _13483_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[27] ),
    .A2(_06046_),
    .B1(_05985_),
    .B2(_06059_),
    .X(_01129_));
 sky130_fd_sc_hd__xnor2_4 _13484_ (.A(_04509_),
    .B(_06056_),
    .Y(_06060_));
 sky130_fd_sc_hd__nand2_1 _13485_ (.A(_06036_),
    .B(_06060_),
    .Y(_06061_));
 sky130_fd_sc_hd__a22o_1 _13486_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[26] ),
    .A2(_06046_),
    .B1(_05985_),
    .B2(_06061_),
    .X(_01128_));
 sky130_fd_sc_hd__or3_4 _13487_ (.A(_04597_),
    .B(_05282_),
    .C(_06055_),
    .X(_06062_));
 sky130_fd_sc_hd__o21ai_4 _13488_ (.A1(_05282_),
    .A2(_06055_),
    .B1(_04597_),
    .Y(_06063_));
 sky130_fd_sc_hd__buf_2 _13489_ (.A(_06035_),
    .X(_06064_));
 sky130_fd_sc_hd__a21bo_1 _13490_ (.A1(_06062_),
    .A2(_06063_),
    .B1_N(_06064_),
    .X(_06065_));
 sky130_fd_sc_hd__a22o_1 _13491_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[25] ),
    .A2(_06046_),
    .B1(_05985_),
    .B2(_06065_),
    .X(_01127_));
 sky130_fd_sc_hd__nor2_2 _13492_ (.A(_04676_),
    .B(_06039_),
    .Y(_06066_));
 sky130_fd_sc_hd__o21ai_1 _13493_ (.A1(_06055_),
    .A2(_06066_),
    .B1(_06064_),
    .Y(_06067_));
 sky130_fd_sc_hd__a22o_1 _13494_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[24] ),
    .A2(_06046_),
    .B1(_05985_),
    .B2(_06067_),
    .X(_01126_));
 sky130_fd_sc_hd__or2b_2 _13495_ (.A(_05276_),
    .B_N(_06038_),
    .X(_06068_));
 sky130_fd_sc_hd__a31o_2 _13496_ (.A1(_04919_),
    .A2(_04997_),
    .A3(_06068_),
    .B1(_05277_),
    .X(_06069_));
 sky130_fd_sc_hd__a21oi_2 _13497_ (.A1(_04839_),
    .A2(_06069_),
    .B1(_04837_),
    .Y(_06070_));
 sky130_fd_sc_hd__xnor2_4 _13498_ (.A(_04760_),
    .B(_06070_),
    .Y(_06071_));
 sky130_fd_sc_hd__or2b_1 _13499_ (.A(_06071_),
    .B_N(_06064_),
    .X(_06072_));
 sky130_fd_sc_hd__a22o_1 _13500_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[23] ),
    .A2(_06046_),
    .B1(_05985_),
    .B2(_06072_),
    .X(_01125_));
 sky130_fd_sc_hd__xnor2_4 _13501_ (.A(_04839_),
    .B(_06069_),
    .Y(_06073_));
 sky130_fd_sc_hd__nand2_1 _13502_ (.A(_06036_),
    .B(_06073_),
    .Y(_06074_));
 sky130_fd_sc_hd__a22o_1 _13503_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[22] ),
    .A2(_06046_),
    .B1(_05985_),
    .B2(_06074_),
    .X(_01124_));
 sky130_fd_sc_hd__clkbuf_4 _13504_ (.A(_05984_),
    .X(_06075_));
 sky130_fd_sc_hd__and2_1 _13505_ (.A(_04997_),
    .B(_06068_),
    .X(_06076_));
 sky130_fd_sc_hd__nor2_2 _13506_ (.A(_04995_),
    .B(_06076_),
    .Y(_06077_));
 sky130_fd_sc_hd__xor2_4 _13507_ (.A(_04919_),
    .B(_06077_),
    .X(_06078_));
 sky130_fd_sc_hd__nand2_1 _13508_ (.A(_06036_),
    .B(_06078_),
    .Y(_06079_));
 sky130_fd_sc_hd__a22o_1 _13509_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[21] ),
    .A2(_06046_),
    .B1(_06075_),
    .B2(_06079_),
    .X(_01123_));
 sky130_fd_sc_hd__clkbuf_4 _13510_ (.A(_05981_),
    .X(_06080_));
 sky130_fd_sc_hd__xnor2_4 _13511_ (.A(_04997_),
    .B(_06068_),
    .Y(_06081_));
 sky130_fd_sc_hd__nand2_1 _13512_ (.A(_06036_),
    .B(_06081_),
    .Y(_06082_));
 sky130_fd_sc_hd__a22o_1 _13513_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[20] ),
    .A2(_06080_),
    .B1(_06075_),
    .B2(_06082_),
    .X(_01122_));
 sky130_fd_sc_hd__nor2_2 _13514_ (.A(_05142_),
    .B(_05143_),
    .Y(_06083_));
 sky130_fd_sc_hd__and3_1 _13515_ (.A(_05689_),
    .B(_05691_),
    .C(_06037_),
    .X(_06084_));
 sky130_fd_sc_hd__or2b_2 _13516_ (.A(_06084_),
    .B_N(_05274_),
    .X(_06085_));
 sky130_fd_sc_hd__a21oi_2 _13517_ (.A1(_06083_),
    .A2(_06085_),
    .B1(_05142_),
    .Y(_06086_));
 sky130_fd_sc_hd__xnor2_4 _13518_ (.A(_05071_),
    .B(_06086_),
    .Y(_06087_));
 sky130_fd_sc_hd__nand2_1 _13519_ (.A(_06036_),
    .B(_06087_),
    .Y(_06088_));
 sky130_fd_sc_hd__a22o_1 _13520_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[19] ),
    .A2(_06080_),
    .B1(_06075_),
    .B2(_06088_),
    .X(_01121_));
 sky130_fd_sc_hd__xnor2_4 _13521_ (.A(_06083_),
    .B(_06085_),
    .Y(_06089_));
 sky130_fd_sc_hd__nand2_1 _13522_ (.A(_06036_),
    .B(_06089_),
    .Y(_06090_));
 sky130_fd_sc_hd__a22o_1 _13523_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[18] ),
    .A2(_06080_),
    .B1(_06075_),
    .B2(_06090_),
    .X(_01120_));
 sky130_fd_sc_hd__a21o_1 _13524_ (.A1(_05689_),
    .A2(_06037_),
    .B1(_05268_),
    .X(_06091_));
 sky130_fd_sc_hd__xnor2_4 _13525_ (.A(_05691_),
    .B(_06091_),
    .Y(_06092_));
 sky130_fd_sc_hd__nand2_1 _13526_ (.A(_06053_),
    .B(_06092_),
    .Y(_06093_));
 sky130_fd_sc_hd__a22o_1 _13527_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[17] ),
    .A2(_06080_),
    .B1(_06075_),
    .B2(_06093_),
    .X(_01119_));
 sky130_fd_sc_hd__xnor2_4 _13528_ (.A(_05689_),
    .B(_06037_),
    .Y(_06094_));
 sky130_fd_sc_hd__nand2_1 _13529_ (.A(_06053_),
    .B(_06094_),
    .Y(_06095_));
 sky130_fd_sc_hd__a22o_1 _13530_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[16] ),
    .A2(_06080_),
    .B1(_06075_),
    .B2(_06095_),
    .X(_01118_));
 sky130_fd_sc_hd__and2b_1 _13531_ (.A_N(_05684_),
    .B(_05666_),
    .X(_06096_));
 sky130_fd_sc_hd__o21ba_1 _13532_ (.A1(_05696_),
    .A2(_06096_),
    .B1_N(_05681_),
    .X(_06097_));
 sky130_fd_sc_hd__xnor2_2 _13533_ (.A(_05694_),
    .B(_06097_),
    .Y(_06098_));
 sky130_fd_sc_hd__nand2_1 _13534_ (.A(_06053_),
    .B(_06098_),
    .Y(_06099_));
 sky130_fd_sc_hd__a22o_1 _13535_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[15] ),
    .A2(_06080_),
    .B1(_06075_),
    .B2(_06099_),
    .X(_01117_));
 sky130_fd_sc_hd__xnor2_2 _13536_ (.A(_05696_),
    .B(_06096_),
    .Y(_06100_));
 sky130_fd_sc_hd__nand2_1 _13537_ (.A(_06053_),
    .B(_06100_),
    .Y(_06101_));
 sky130_fd_sc_hd__a22o_1 _13538_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[14] ),
    .A2(_06080_),
    .B1(_06075_),
    .B2(_06101_),
    .X(_01116_));
 sky130_fd_sc_hd__or2_1 _13539_ (.A(_05504_),
    .B(_05665_),
    .X(_06102_));
 sky130_fd_sc_hd__o21bai_1 _13540_ (.A1(_05471_),
    .A2(_06102_),
    .B1_N(_05469_),
    .Y(_06103_));
 sky130_fd_sc_hd__xor2_2 _13541_ (.A(_05430_),
    .B(_06103_),
    .X(_06104_));
 sky130_fd_sc_hd__nand2_1 _13542_ (.A(_06053_),
    .B(_06104_),
    .Y(_06105_));
 sky130_fd_sc_hd__a22o_1 _13543_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[13] ),
    .A2(_06080_),
    .B1(_06075_),
    .B2(_06105_),
    .X(_01115_));
 sky130_fd_sc_hd__xor2_2 _13544_ (.A(_05471_),
    .B(_06102_),
    .X(_06106_));
 sky130_fd_sc_hd__or2b_1 _13545_ (.A(_06106_),
    .B_N(_06064_),
    .X(_06107_));
 sky130_fd_sc_hd__a22o_1 _13546_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[12] ),
    .A2(_06080_),
    .B1(_06075_),
    .B2(_06107_),
    .X(_01114_));
 sky130_fd_sc_hd__clkbuf_4 _13547_ (.A(_05984_),
    .X(_06108_));
 sky130_fd_sc_hd__or2_1 _13548_ (.A(_05537_),
    .B(_05661_),
    .X(_06109_));
 sky130_fd_sc_hd__nor2_1 _13549_ (.A(_05504_),
    .B(_05662_),
    .Y(_06110_));
 sky130_fd_sc_hd__and3_1 _13550_ (.A(_05664_),
    .B(_06109_),
    .C(_06110_),
    .X(_06111_));
 sky130_fd_sc_hd__a21oi_1 _13551_ (.A1(_05664_),
    .A2(_06109_),
    .B1(_06110_),
    .Y(_06112_));
 sky130_fd_sc_hd__or3b_1 _13552_ (.A(_06111_),
    .B(_06112_),
    .C_N(_06035_),
    .X(_06113_));
 sky130_fd_sc_hd__a22o_1 _13553_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[11] ),
    .A2(_06080_),
    .B1(_06108_),
    .B2(_06113_),
    .X(_01113_));
 sky130_fd_sc_hd__clkbuf_4 _13554_ (.A(_05981_),
    .X(_06114_));
 sky130_fd_sc_hd__nand2_1 _13555_ (.A(_05537_),
    .B(_05661_),
    .Y(_06115_));
 sky130_fd_sc_hd__a21bo_1 _13556_ (.A1(_06109_),
    .A2(_06115_),
    .B1_N(_06064_),
    .X(_06116_));
 sky130_fd_sc_hd__a22o_1 _13557_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[10] ),
    .A2(_06114_),
    .B1(_06108_),
    .B2(_06116_),
    .X(_01112_));
 sky130_fd_sc_hd__xnor2_1 _13558_ (.A(_05564_),
    .B(_05659_),
    .Y(_06117_));
 sky130_fd_sc_hd__nand2_1 _13559_ (.A(_06053_),
    .B(_06117_),
    .Y(_06118_));
 sky130_fd_sc_hd__a22o_1 _13560_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[9] ),
    .A2(_06114_),
    .B1(_06108_),
    .B2(_06118_),
    .X(_01111_));
 sky130_fd_sc_hd__and2b_1 _13561_ (.A_N(_05658_),
    .B(_05589_),
    .X(_06119_));
 sky130_fd_sc_hd__xnor2_1 _13562_ (.A(_06119_),
    .B(_05657_),
    .Y(_06120_));
 sky130_fd_sc_hd__nand2_1 _13563_ (.A(_06053_),
    .B(_06120_),
    .Y(_06121_));
 sky130_fd_sc_hd__a22o_1 _13564_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[8] ),
    .A2(_06114_),
    .B1(_06108_),
    .B2(_06121_),
    .X(_01110_));
 sky130_fd_sc_hd__and2b_1 _13565_ (.A_N(_05656_),
    .B(_05610_),
    .X(_06122_));
 sky130_fd_sc_hd__xnor2_1 _13566_ (.A(_06122_),
    .B(_05655_),
    .Y(_06123_));
 sky130_fd_sc_hd__nand2_1 _13567_ (.A(_06053_),
    .B(_06123_),
    .Y(_06124_));
 sky130_fd_sc_hd__a22o_1 _13568_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[7] ),
    .A2(_06114_),
    .B1(_06108_),
    .B2(_06124_),
    .X(_01109_));
 sky130_fd_sc_hd__or3_1 _13569_ (.A(_05654_),
    .B(_05626_),
    .C(_05653_),
    .X(_06125_));
 sky130_fd_sc_hd__o21ai_1 _13570_ (.A1(_05654_),
    .A2(_05626_),
    .B1(_05653_),
    .Y(_06126_));
 sky130_fd_sc_hd__a21bo_1 _13571_ (.A1(_06125_),
    .A2(_06126_),
    .B1_N(_06064_),
    .X(_06127_));
 sky130_fd_sc_hd__a22o_1 _13572_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[6] ),
    .A2(_06114_),
    .B1(_06108_),
    .B2(_06127_),
    .X(_01108_));
 sky130_fd_sc_hd__and2b_1 _13573_ (.A_N(_05652_),
    .B(_05639_),
    .X(_06128_));
 sky130_fd_sc_hd__xnor2_1 _13574_ (.A(_06128_),
    .B(_05651_),
    .Y(_06129_));
 sky130_fd_sc_hd__nand2_1 _13575_ (.A(_06053_),
    .B(_06129_),
    .Y(_06130_));
 sky130_fd_sc_hd__a22o_1 _13576_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[5] ),
    .A2(_06114_),
    .B1(_06108_),
    .B2(_06130_),
    .X(_01107_));
 sky130_fd_sc_hd__and3_1 _13577_ (.A(_05640_),
    .B(_05645_),
    .C(_05649_),
    .X(_06131_));
 sky130_fd_sc_hd__a21oi_1 _13578_ (.A1(_05640_),
    .A2(_05649_),
    .B1(_05645_),
    .Y(_06132_));
 sky130_fd_sc_hd__o21ai_1 _13579_ (.A1(_06131_),
    .A2(_06132_),
    .B1(_06064_),
    .Y(_06133_));
 sky130_fd_sc_hd__a22o_1 _13580_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[4] ),
    .A2(_06114_),
    .B1(_06108_),
    .B2(_06133_),
    .X(_01106_));
 sky130_fd_sc_hd__or3_1 _13581_ (.A(_05640_),
    .B(_05643_),
    .C(_05649_),
    .X(_06134_));
 sky130_fd_sc_hd__o21ai_1 _13582_ (.A1(_05643_),
    .A2(_05649_),
    .B1(_05640_),
    .Y(_06135_));
 sky130_fd_sc_hd__a21bo_1 _13583_ (.A1(_06134_),
    .A2(_06135_),
    .B1_N(_06064_),
    .X(_06136_));
 sky130_fd_sc_hd__a22o_1 _13584_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[3] ),
    .A2(_06114_),
    .B1(_06108_),
    .B2(_06136_),
    .X(_01105_));
 sky130_fd_sc_hd__a21oi_1 _13585_ (.A1(_05646_),
    .A2(_05647_),
    .B1(_05648_),
    .Y(_06137_));
 sky130_fd_sc_hd__o21ai_1 _13586_ (.A1(_05649_),
    .A2(_06137_),
    .B1(_06064_),
    .Y(_06138_));
 sky130_fd_sc_hd__a22o_1 _13587_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[2] ),
    .A2(_06114_),
    .B1(_06108_),
    .B2(_06138_),
    .X(_01104_));
 sky130_fd_sc_hd__a21boi_1 _13588_ (.A1(_04081_),
    .A2(_05292_),
    .B1_N(_05633_),
    .Y(_06139_));
 sky130_fd_sc_hd__o21ai_1 _13589_ (.A1(_05648_),
    .A2(_06139_),
    .B1(_06064_),
    .Y(_06140_));
 sky130_fd_sc_hd__a22o_1 _13590_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[1] ),
    .A2(_06114_),
    .B1(_05984_),
    .B2(_06140_),
    .X(_01103_));
 sky130_fd_sc_hd__a21bo_1 _13591_ (.A1(_04081_),
    .A2(_05147_),
    .B1_N(_06035_),
    .X(_06141_));
 sky130_fd_sc_hd__a22o_1 _13592_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[0] ),
    .A2(_05981_),
    .B1(_05984_),
    .B2(_06141_),
    .X(_01102_));
 sky130_fd_sc_hd__clkbuf_4 _13593_ (.A(\wfg_stim_mem_top.wfg_stim_mem.cur_state[1] ),
    .X(_06142_));
 sky130_fd_sc_hd__mux2_1 _13594_ (.A0(\wfg_interconnect_top.stimulus_1[31] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[31] ),
    .S(_06142_),
    .X(_06143_));
 sky130_fd_sc_hd__clkbuf_1 _13595_ (.A(_06143_),
    .X(_01101_));
 sky130_fd_sc_hd__mux2_1 _13596_ (.A0(\wfg_interconnect_top.stimulus_1[30] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[30] ),
    .S(_06142_),
    .X(_06144_));
 sky130_fd_sc_hd__clkbuf_1 _13597_ (.A(_06144_),
    .X(_01100_));
 sky130_fd_sc_hd__mux2_1 _13598_ (.A0(\wfg_interconnect_top.stimulus_1[29] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[29] ),
    .S(_06142_),
    .X(_06145_));
 sky130_fd_sc_hd__clkbuf_1 _13599_ (.A(_06145_),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_1 _13600_ (.A0(\wfg_interconnect_top.stimulus_1[28] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[28] ),
    .S(_06142_),
    .X(_06146_));
 sky130_fd_sc_hd__clkbuf_1 _13601_ (.A(_06146_),
    .X(_01098_));
 sky130_fd_sc_hd__mux2_1 _13602_ (.A0(\wfg_interconnect_top.stimulus_1[27] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[27] ),
    .S(_06142_),
    .X(_06147_));
 sky130_fd_sc_hd__clkbuf_1 _13603_ (.A(_06147_),
    .X(_01097_));
 sky130_fd_sc_hd__mux2_1 _13604_ (.A0(\wfg_interconnect_top.stimulus_1[26] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[26] ),
    .S(_06142_),
    .X(_06148_));
 sky130_fd_sc_hd__clkbuf_1 _13605_ (.A(_06148_),
    .X(_01096_));
 sky130_fd_sc_hd__mux2_1 _13606_ (.A0(\wfg_interconnect_top.stimulus_1[25] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[25] ),
    .S(_06142_),
    .X(_06149_));
 sky130_fd_sc_hd__clkbuf_1 _13607_ (.A(_06149_),
    .X(_01095_));
 sky130_fd_sc_hd__mux2_1 _13608_ (.A0(\wfg_interconnect_top.stimulus_1[24] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[24] ),
    .S(_06142_),
    .X(_06150_));
 sky130_fd_sc_hd__clkbuf_1 _13609_ (.A(_06150_),
    .X(_01094_));
 sky130_fd_sc_hd__mux2_1 _13610_ (.A0(\wfg_interconnect_top.stimulus_1[23] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[23] ),
    .S(_06142_),
    .X(_06151_));
 sky130_fd_sc_hd__clkbuf_1 _13611_ (.A(_06151_),
    .X(_01093_));
 sky130_fd_sc_hd__mux2_1 _13612_ (.A0(\wfg_interconnect_top.stimulus_1[22] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[22] ),
    .S(_06142_),
    .X(_06152_));
 sky130_fd_sc_hd__clkbuf_1 _13613_ (.A(_06152_),
    .X(_01092_));
 sky130_fd_sc_hd__buf_4 _13614_ (.A(\wfg_stim_mem_top.wfg_stim_mem.cur_state[1] ),
    .X(_06153_));
 sky130_fd_sc_hd__mux2_1 _13615_ (.A0(\wfg_interconnect_top.stimulus_1[21] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[21] ),
    .S(_06153_),
    .X(_06154_));
 sky130_fd_sc_hd__clkbuf_1 _13616_ (.A(_06154_),
    .X(_01091_));
 sky130_fd_sc_hd__mux2_1 _13617_ (.A0(\wfg_interconnect_top.stimulus_1[20] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[20] ),
    .S(_06153_),
    .X(_06155_));
 sky130_fd_sc_hd__clkbuf_1 _13618_ (.A(_06155_),
    .X(_01090_));
 sky130_fd_sc_hd__mux2_1 _13619_ (.A0(\wfg_interconnect_top.stimulus_1[19] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[19] ),
    .S(_06153_),
    .X(_06156_));
 sky130_fd_sc_hd__clkbuf_1 _13620_ (.A(_06156_),
    .X(_01089_));
 sky130_fd_sc_hd__mux2_1 _13621_ (.A0(\wfg_interconnect_top.stimulus_1[18] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[18] ),
    .S(_06153_),
    .X(_06157_));
 sky130_fd_sc_hd__clkbuf_1 _13622_ (.A(_06157_),
    .X(_01088_));
 sky130_fd_sc_hd__mux2_1 _13623_ (.A0(\wfg_interconnect_top.stimulus_1[17] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[17] ),
    .S(_06153_),
    .X(_06158_));
 sky130_fd_sc_hd__clkbuf_1 _13624_ (.A(_06158_),
    .X(_01087_));
 sky130_fd_sc_hd__mux2_1 _13625_ (.A0(\wfg_interconnect_top.stimulus_1[16] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[16] ),
    .S(_06153_),
    .X(_06159_));
 sky130_fd_sc_hd__clkbuf_1 _13626_ (.A(_06159_),
    .X(_01086_));
 sky130_fd_sc_hd__mux2_1 _13627_ (.A0(\wfg_interconnect_top.stimulus_1[15] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[15] ),
    .S(_06153_),
    .X(_06160_));
 sky130_fd_sc_hd__clkbuf_1 _13628_ (.A(_06160_),
    .X(_01085_));
 sky130_fd_sc_hd__mux2_1 _13629_ (.A0(\wfg_interconnect_top.stimulus_1[14] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[14] ),
    .S(_06153_),
    .X(_06161_));
 sky130_fd_sc_hd__clkbuf_1 _13630_ (.A(_06161_),
    .X(_01084_));
 sky130_fd_sc_hd__mux2_1 _13631_ (.A0(\wfg_interconnect_top.stimulus_1[13] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[13] ),
    .S(_06153_),
    .X(_06162_));
 sky130_fd_sc_hd__clkbuf_1 _13632_ (.A(_06162_),
    .X(_01083_));
 sky130_fd_sc_hd__mux2_1 _13633_ (.A0(\wfg_interconnect_top.stimulus_1[12] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[12] ),
    .S(_06153_),
    .X(_06163_));
 sky130_fd_sc_hd__clkbuf_1 _13634_ (.A(_06163_),
    .X(_01082_));
 sky130_fd_sc_hd__clkbuf_4 _13635_ (.A(\wfg_stim_mem_top.wfg_stim_mem.cur_state[1] ),
    .X(_06164_));
 sky130_fd_sc_hd__mux2_1 _13636_ (.A0(\wfg_interconnect_top.stimulus_1[11] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[11] ),
    .S(_06164_),
    .X(_06165_));
 sky130_fd_sc_hd__clkbuf_1 _13637_ (.A(_06165_),
    .X(_01081_));
 sky130_fd_sc_hd__mux2_1 _13638_ (.A0(\wfg_interconnect_top.stimulus_1[10] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[10] ),
    .S(_06164_),
    .X(_06166_));
 sky130_fd_sc_hd__clkbuf_1 _13639_ (.A(_06166_),
    .X(_01080_));
 sky130_fd_sc_hd__mux2_1 _13640_ (.A0(\wfg_interconnect_top.stimulus_1[9] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[9] ),
    .S(_06164_),
    .X(_06167_));
 sky130_fd_sc_hd__clkbuf_1 _13641_ (.A(_06167_),
    .X(_01079_));
 sky130_fd_sc_hd__mux2_1 _13642_ (.A0(\wfg_interconnect_top.stimulus_1[8] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[8] ),
    .S(_06164_),
    .X(_06168_));
 sky130_fd_sc_hd__clkbuf_1 _13643_ (.A(_06168_),
    .X(_01078_));
 sky130_fd_sc_hd__mux2_1 _13644_ (.A0(\wfg_interconnect_top.stimulus_1[7] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[7] ),
    .S(_06164_),
    .X(_06169_));
 sky130_fd_sc_hd__clkbuf_1 _13645_ (.A(_06169_),
    .X(_01077_));
 sky130_fd_sc_hd__mux2_1 _13646_ (.A0(\wfg_interconnect_top.stimulus_1[6] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[6] ),
    .S(_06164_),
    .X(_06170_));
 sky130_fd_sc_hd__clkbuf_1 _13647_ (.A(_06170_),
    .X(_01076_));
 sky130_fd_sc_hd__mux2_1 _13648_ (.A0(\wfg_interconnect_top.stimulus_1[5] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[5] ),
    .S(_06164_),
    .X(_06171_));
 sky130_fd_sc_hd__clkbuf_1 _13649_ (.A(_06171_),
    .X(_01075_));
 sky130_fd_sc_hd__mux2_1 _13650_ (.A0(\wfg_interconnect_top.stimulus_1[4] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[4] ),
    .S(_06164_),
    .X(_06172_));
 sky130_fd_sc_hd__clkbuf_1 _13651_ (.A(_06172_),
    .X(_01074_));
 sky130_fd_sc_hd__mux2_1 _13652_ (.A0(\wfg_interconnect_top.stimulus_1[3] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[3] ),
    .S(_06164_),
    .X(_06173_));
 sky130_fd_sc_hd__clkbuf_1 _13653_ (.A(_06173_),
    .X(_01073_));
 sky130_fd_sc_hd__mux2_1 _13654_ (.A0(\wfg_interconnect_top.stimulus_1[2] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[2] ),
    .S(_06164_),
    .X(_06174_));
 sky130_fd_sc_hd__clkbuf_1 _13655_ (.A(_06174_),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_1 _13656_ (.A0(\wfg_interconnect_top.stimulus_1[1] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[1] ),
    .S(\wfg_stim_mem_top.wfg_stim_mem.cur_state[1] ),
    .X(_06175_));
 sky130_fd_sc_hd__clkbuf_1 _13657_ (.A(_06175_),
    .X(_01071_));
 sky130_fd_sc_hd__mux2_1 _13658_ (.A0(\wfg_interconnect_top.stimulus_1[0] ),
    .A1(\wfg_stim_mem_top.wfg_stim_mem.data_calc[0] ),
    .S(\wfg_stim_mem_top.wfg_stim_mem.cur_state[1] ),
    .X(_06176_));
 sky130_fd_sc_hd__clkbuf_1 _13659_ (.A(_06176_),
    .X(_01070_));
 sky130_fd_sc_hd__inv_2 _13660_ (.A(net110),
    .Y(_06177_));
 sky130_fd_sc_hd__nor2_1 _13661_ (.A(\wfg_stim_mem_top.cfg_inc_q[7] ),
    .B(net108),
    .Y(_06178_));
 sky130_fd_sc_hd__nor2_1 _13662_ (.A(\wfg_stim_mem_top.cfg_inc_q[6] ),
    .B(net107),
    .Y(_06179_));
 sky130_fd_sc_hd__nand2_1 _13663_ (.A(\wfg_stim_mem_top.cfg_inc_q[5] ),
    .B(net106),
    .Y(_06180_));
 sky130_fd_sc_hd__or2_1 _13664_ (.A(\wfg_stim_mem_top.cfg_inc_q[5] ),
    .B(net106),
    .X(_06181_));
 sky130_fd_sc_hd__nand2_1 _13665_ (.A(_06180_),
    .B(_06181_),
    .Y(_06182_));
 sky130_fd_sc_hd__nand2_1 _13666_ (.A(\wfg_stim_mem_top.cfg_inc_q[4] ),
    .B(net105),
    .Y(_06183_));
 sky130_fd_sc_hd__or2_1 _13667_ (.A(\wfg_stim_mem_top.cfg_inc_q[4] ),
    .B(net105),
    .X(_06184_));
 sky130_fd_sc_hd__nand2_1 _13668_ (.A(_06183_),
    .B(_06184_),
    .Y(_06185_));
 sky130_fd_sc_hd__nor2_1 _13669_ (.A(\wfg_stim_mem_top.cfg_inc_q[2] ),
    .B(net103),
    .Y(_06186_));
 sky130_fd_sc_hd__nand2_1 _13670_ (.A(\wfg_stim_mem_top.cfg_inc_q[1] ),
    .B(net102),
    .Y(_06187_));
 sky130_fd_sc_hd__or2_1 _13671_ (.A(\wfg_stim_mem_top.cfg_inc_q[1] ),
    .B(net102),
    .X(_06188_));
 sky130_fd_sc_hd__nand2_1 _13672_ (.A(_06187_),
    .B(_06188_),
    .Y(_06189_));
 sky130_fd_sc_hd__nand2_1 _13673_ (.A(\wfg_stim_mem_top.cfg_inc_q[0] ),
    .B(net101),
    .Y(_06190_));
 sky130_fd_sc_hd__o21a_1 _13674_ (.A1(_06189_),
    .A2(_06190_),
    .B1(_06187_),
    .X(_06191_));
 sky130_fd_sc_hd__nand2_1 _13675_ (.A(\wfg_stim_mem_top.cfg_inc_q[2] ),
    .B(net103),
    .Y(_06192_));
 sky130_fd_sc_hd__o21ai_2 _13676_ (.A1(_06186_),
    .A2(_06191_),
    .B1(_06192_),
    .Y(_06193_));
 sky130_fd_sc_hd__a21o_1 _13677_ (.A1(\wfg_stim_mem_top.cfg_inc_q[3] ),
    .A2(net104),
    .B1(_06193_),
    .X(_06194_));
 sky130_fd_sc_hd__o21ai_2 _13678_ (.A1(\wfg_stim_mem_top.cfg_inc_q[3] ),
    .A2(net104),
    .B1(_06194_),
    .Y(_06195_));
 sky130_fd_sc_hd__o21a_1 _13679_ (.A1(_06185_),
    .A2(_06195_),
    .B1(_06183_),
    .X(_06196_));
 sky130_fd_sc_hd__o21a_1 _13680_ (.A1(_06182_),
    .A2(_06196_),
    .B1(_06180_),
    .X(_06197_));
 sky130_fd_sc_hd__nand2_1 _13681_ (.A(\wfg_stim_mem_top.cfg_inc_q[6] ),
    .B(net107),
    .Y(_06198_));
 sky130_fd_sc_hd__o21a_1 _13682_ (.A1(_06179_),
    .A2(_06197_),
    .B1(_06198_),
    .X(_06199_));
 sky130_fd_sc_hd__nand2_1 _13683_ (.A(\wfg_stim_mem_top.cfg_inc_q[7] ),
    .B(net108),
    .Y(_06200_));
 sky130_fd_sc_hd__o21ai_1 _13684_ (.A1(_06178_),
    .A2(_06199_),
    .B1(_06200_),
    .Y(_06201_));
 sky130_fd_sc_hd__nand2_1 _13685_ (.A(net109),
    .B(_06201_),
    .Y(_06202_));
 sky130_fd_sc_hd__nor2_1 _13686_ (.A(_06177_),
    .B(_06202_),
    .Y(_06203_));
 sky130_fd_sc_hd__and2_1 _13687_ (.A(\wfg_stim_mem_top.wfg_stim_mem.cur_address[10] ),
    .B(_06203_),
    .X(_06204_));
 sky130_fd_sc_hd__and3_1 _13688_ (.A(\wfg_stim_mem_top.wfg_stim_mem.cur_address[12] ),
    .B(\wfg_stim_mem_top.wfg_stim_mem.cur_address[11] ),
    .C(_06204_),
    .X(_06205_));
 sky130_fd_sc_hd__and2_1 _13689_ (.A(\wfg_stim_mem_top.wfg_stim_mem.cur_address[13] ),
    .B(_06205_),
    .X(_06206_));
 sky130_fd_sc_hd__nand2_1 _13690_ (.A(\wfg_stim_mem_top.wfg_stim_mem.cur_address[14] ),
    .B(_06206_),
    .Y(_06207_));
 sky130_fd_sc_hd__xor2_2 _13691_ (.A(\wfg_stim_mem_top.wfg_stim_mem.cur_address[15] ),
    .B(_06207_),
    .X(_06208_));
 sky130_fd_sc_hd__nor2_1 _13692_ (.A(\wfg_stim_mem_top.wfg_stim_mem.cur_address[13] ),
    .B(_06205_),
    .Y(_06209_));
 sky130_fd_sc_hd__or2_1 _13693_ (.A(_06206_),
    .B(_06209_),
    .X(_06210_));
 sky130_fd_sc_hd__or2_1 _13694_ (.A(\wfg_stim_mem_top.wfg_stim_mem.cur_address[14] ),
    .B(_06206_),
    .X(_06211_));
 sky130_fd_sc_hd__nand2_1 _13695_ (.A(_06207_),
    .B(_06211_),
    .Y(_06212_));
 sky130_fd_sc_hd__a21oi_1 _13696_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.cur_address[11] ),
    .A2(_06204_),
    .B1(\wfg_stim_mem_top.wfg_stim_mem.cur_address[12] ),
    .Y(_06213_));
 sky130_fd_sc_hd__or2_1 _13697_ (.A(_06205_),
    .B(_06213_),
    .X(_06214_));
 sky130_fd_sc_hd__xnor2_2 _13698_ (.A(\wfg_stim_mem_top.wfg_stim_mem.cur_address[11] ),
    .B(_06204_),
    .Y(_06215_));
 sky130_fd_sc_hd__nor2_1 _13699_ (.A(\wfg_stim_mem_top.wfg_stim_mem.cur_address[10] ),
    .B(_06203_),
    .Y(_06216_));
 sky130_fd_sc_hd__or2_1 _13700_ (.A(_06204_),
    .B(_06216_),
    .X(_06217_));
 sky130_fd_sc_hd__or2_1 _13701_ (.A(\wfg_stim_mem_top.end_val_q[10] ),
    .B(_06217_),
    .X(_06218_));
 sky130_fd_sc_hd__and2_1 _13702_ (.A(_06177_),
    .B(_06202_),
    .X(_06219_));
 sky130_fd_sc_hd__or2_1 _13703_ (.A(_06203_),
    .B(_06219_),
    .X(_06220_));
 sky130_fd_sc_hd__or2_1 _13704_ (.A(net109),
    .B(_06201_),
    .X(_06221_));
 sky130_fd_sc_hd__nand2_1 _13705_ (.A(_06202_),
    .B(_06221_),
    .Y(_06222_));
 sky130_fd_sc_hd__or2b_1 _13706_ (.A(_06178_),
    .B_N(_06200_),
    .X(_06223_));
 sky130_fd_sc_hd__xnor2_2 _13707_ (.A(_06199_),
    .B(_06223_),
    .Y(_06224_));
 sky130_fd_sc_hd__or2b_1 _13708_ (.A(_06179_),
    .B_N(_06198_),
    .X(_06225_));
 sky130_fd_sc_hd__xnor2_2 _13709_ (.A(_06197_),
    .B(_06225_),
    .Y(_06226_));
 sky130_fd_sc_hd__xnor2_1 _13710_ (.A(_06182_),
    .B(_06196_),
    .Y(_06227_));
 sky130_fd_sc_hd__and2_1 _13711_ (.A(\wfg_stim_mem_top.end_val_q[5] ),
    .B(_06227_),
    .X(_06228_));
 sky130_fd_sc_hd__xnor2_2 _13712_ (.A(_06185_),
    .B(_06195_),
    .Y(_06229_));
 sky130_fd_sc_hd__xor2_1 _13713_ (.A(\wfg_stim_mem_top.cfg_inc_q[3] ),
    .B(net104),
    .X(_06230_));
 sky130_fd_sc_hd__xnor2_2 _13714_ (.A(_06193_),
    .B(_06230_),
    .Y(_06231_));
 sky130_fd_sc_hd__or2b_1 _13715_ (.A(_06186_),
    .B_N(_06192_),
    .X(_06232_));
 sky130_fd_sc_hd__xnor2_2 _13716_ (.A(_06191_),
    .B(_06232_),
    .Y(_06233_));
 sky130_fd_sc_hd__xnor2_1 _13717_ (.A(_06189_),
    .B(_06190_),
    .Y(_06234_));
 sky130_fd_sc_hd__or2_1 _13718_ (.A(\wfg_stim_mem_top.cfg_inc_q[0] ),
    .B(net101),
    .X(_06235_));
 sky130_fd_sc_hd__nand2_1 _13719_ (.A(_06190_),
    .B(_06235_),
    .Y(_06236_));
 sky130_fd_sc_hd__a211o_1 _13720_ (.A1(\wfg_stim_mem_top.end_val_q[1] ),
    .A2(_06234_),
    .B1(_06236_),
    .C1(\wfg_stim_mem_top.end_val_q[0] ),
    .X(_06237_));
 sky130_fd_sc_hd__o22a_1 _13721_ (.A1(\wfg_stim_mem_top.end_val_q[2] ),
    .A2(_06233_),
    .B1(_06234_),
    .B2(\wfg_stim_mem_top.end_val_q[1] ),
    .X(_06238_));
 sky130_fd_sc_hd__a22o_1 _13722_ (.A1(\wfg_stim_mem_top.end_val_q[2] ),
    .A2(_06233_),
    .B1(_06237_),
    .B2(_06238_),
    .X(_06239_));
 sky130_fd_sc_hd__o21a_1 _13723_ (.A1(\wfg_stim_mem_top.end_val_q[3] ),
    .A2(_06231_),
    .B1(_06239_),
    .X(_06240_));
 sky130_fd_sc_hd__a221o_1 _13724_ (.A1(\wfg_stim_mem_top.end_val_q[4] ),
    .A2(_06229_),
    .B1(_06231_),
    .B2(\wfg_stim_mem_top.end_val_q[3] ),
    .C1(_06240_),
    .X(_06241_));
 sky130_fd_sc_hd__o221a_1 _13725_ (.A1(\wfg_stim_mem_top.end_val_q[5] ),
    .A2(_06227_),
    .B1(_06229_),
    .B2(\wfg_stim_mem_top.end_val_q[4] ),
    .C1(_06241_),
    .X(_06242_));
 sky130_fd_sc_hd__o22a_1 _13726_ (.A1(\wfg_stim_mem_top.end_val_q[6] ),
    .A2(_06226_),
    .B1(_06228_),
    .B2(_06242_),
    .X(_06243_));
 sky130_fd_sc_hd__a221o_1 _13727_ (.A1(\wfg_stim_mem_top.end_val_q[7] ),
    .A2(_06224_),
    .B1(_06226_),
    .B2(\wfg_stim_mem_top.end_val_q[6] ),
    .C1(_06243_),
    .X(_06244_));
 sky130_fd_sc_hd__o221a_1 _13728_ (.A1(\wfg_stim_mem_top.end_val_q[8] ),
    .A2(_06222_),
    .B1(_06224_),
    .B2(\wfg_stim_mem_top.end_val_q[7] ),
    .C1(_06244_),
    .X(_06245_));
 sky130_fd_sc_hd__a21o_1 _13729_ (.A1(\wfg_stim_mem_top.end_val_q[8] ),
    .A2(_06222_),
    .B1(_06245_),
    .X(_06246_));
 sky130_fd_sc_hd__o21a_1 _13730_ (.A1(\wfg_stim_mem_top.end_val_q[9] ),
    .A2(_06220_),
    .B1(_06246_),
    .X(_06247_));
 sky130_fd_sc_hd__a221o_1 _13731_ (.A1(\wfg_stim_mem_top.end_val_q[10] ),
    .A2(_06217_),
    .B1(_06220_),
    .B2(\wfg_stim_mem_top.end_val_q[9] ),
    .C1(_06247_),
    .X(_06248_));
 sky130_fd_sc_hd__a22o_1 _13732_ (.A1(_06218_),
    .A2(_06248_),
    .B1(_06215_),
    .B2(\wfg_stim_mem_top.end_val_q[11] ),
    .X(_06249_));
 sky130_fd_sc_hd__o221a_1 _13733_ (.A1(\wfg_stim_mem_top.end_val_q[11] ),
    .A2(_06215_),
    .B1(_06214_),
    .B2(\wfg_stim_mem_top.end_val_q[12] ),
    .C1(_06249_),
    .X(_06250_));
 sky130_fd_sc_hd__a221o_1 _13734_ (.A1(\wfg_stim_mem_top.end_val_q[12] ),
    .A2(_06214_),
    .B1(_06210_),
    .B2(\wfg_stim_mem_top.end_val_q[13] ),
    .C1(_06250_),
    .X(_06251_));
 sky130_fd_sc_hd__o221a_1 _13735_ (.A1(\wfg_stim_mem_top.end_val_q[13] ),
    .A2(_06210_),
    .B1(_06212_),
    .B2(\wfg_stim_mem_top.end_val_q[14] ),
    .C1(_06251_),
    .X(_06252_));
 sky130_fd_sc_hd__a22o_1 _13736_ (.A1(\wfg_stim_mem_top.end_val_q[14] ),
    .A2(_06212_),
    .B1(_06208_),
    .B2(\wfg_stim_mem_top.end_val_q[15] ),
    .X(_06253_));
 sky130_fd_sc_hd__o21a_1 _13737_ (.A1(_06252_),
    .A2(_06253_),
    .B1(\wfg_stim_mem_top.wfg_stim_mem.cur_state[2] ),
    .X(_06254_));
 sky130_fd_sc_hd__o21ai_4 _13738_ (.A1(\wfg_stim_mem_top.end_val_q[15] ),
    .A2(_06208_),
    .B1(_06254_),
    .Y(_06255_));
 sky130_fd_sc_hd__clkinv_2 _13739_ (.A(_06255_),
    .Y(_06256_));
 sky130_fd_sc_hd__o2bb2a_1 _13740_ (.A1_N(_06208_),
    .A2_N(_06254_),
    .B1(_06256_),
    .B2(\wfg_stim_mem_top.start_val_q[15] ),
    .X(_06257_));
 sky130_fd_sc_hd__o21ba_4 _13741_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.cur_state[2] ),
    .A2(\wfg_stim_mem_top.wfg_stim_mem.cur_state[0] ),
    .B1_N(_00000_),
    .X(_06258_));
 sky130_fd_sc_hd__buf_4 _13742_ (.A(_06258_),
    .X(_06259_));
 sky130_fd_sc_hd__mux2_1 _13743_ (.A0(\wfg_stim_mem_top.wfg_stim_mem.cur_address[15] ),
    .A1(_06257_),
    .S(_06259_),
    .X(_06260_));
 sky130_fd_sc_hd__clkbuf_1 _13744_ (.A(_06260_),
    .X(_01069_));
 sky130_fd_sc_hd__clkinv_2 _13745_ (.A(_06212_),
    .Y(_06261_));
 sky130_fd_sc_hd__buf_4 _13746_ (.A(_06255_),
    .X(_06262_));
 sky130_fd_sc_hd__mux2_1 _13747_ (.A0(_06261_),
    .A1(\wfg_stim_mem_top.start_val_q[14] ),
    .S(_06262_),
    .X(_06263_));
 sky130_fd_sc_hd__mux2_1 _13748_ (.A0(\wfg_stim_mem_top.wfg_stim_mem.cur_address[14] ),
    .A1(_06263_),
    .S(_06259_),
    .X(_06264_));
 sky130_fd_sc_hd__clkbuf_1 _13749_ (.A(_06264_),
    .X(_01068_));
 sky130_fd_sc_hd__clkinv_2 _13750_ (.A(_06210_),
    .Y(_06265_));
 sky130_fd_sc_hd__mux2_1 _13751_ (.A0(_06265_),
    .A1(\wfg_stim_mem_top.start_val_q[13] ),
    .S(_06262_),
    .X(_06266_));
 sky130_fd_sc_hd__mux2_1 _13752_ (.A0(\wfg_stim_mem_top.wfg_stim_mem.cur_address[13] ),
    .A1(_06266_),
    .S(_06259_),
    .X(_06267_));
 sky130_fd_sc_hd__clkbuf_1 _13753_ (.A(_06267_),
    .X(_01067_));
 sky130_fd_sc_hd__and2_1 _13754_ (.A(\wfg_stim_mem_top.start_val_q[12] ),
    .B(_06262_),
    .X(_06268_));
 sky130_fd_sc_hd__o21ai_1 _13755_ (.A1(_06214_),
    .A2(_06262_),
    .B1(_06259_),
    .Y(_06269_));
 sky130_fd_sc_hd__o22a_1 _13756_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.cur_address[12] ),
    .A2(_06259_),
    .B1(_06268_),
    .B2(_06269_),
    .X(_01066_));
 sky130_fd_sc_hd__clkinv_2 _13757_ (.A(_06215_),
    .Y(_06270_));
 sky130_fd_sc_hd__mux2_1 _13758_ (.A0(_06270_),
    .A1(\wfg_stim_mem_top.start_val_q[11] ),
    .S(_06262_),
    .X(_06271_));
 sky130_fd_sc_hd__mux2_1 _13759_ (.A0(\wfg_stim_mem_top.wfg_stim_mem.cur_address[11] ),
    .A1(_06271_),
    .S(_06259_),
    .X(_06272_));
 sky130_fd_sc_hd__clkbuf_1 _13760_ (.A(_06272_),
    .X(_01065_));
 sky130_fd_sc_hd__clkinv_2 _13761_ (.A(_06217_),
    .Y(_06273_));
 sky130_fd_sc_hd__mux2_1 _13762_ (.A0(_06273_),
    .A1(\wfg_stim_mem_top.start_val_q[10] ),
    .S(_06262_),
    .X(_06274_));
 sky130_fd_sc_hd__mux2_1 _13763_ (.A0(\wfg_stim_mem_top.wfg_stim_mem.cur_address[10] ),
    .A1(_06274_),
    .S(_06259_),
    .X(_06275_));
 sky130_fd_sc_hd__clkbuf_1 _13764_ (.A(_06275_),
    .X(_01064_));
 sky130_fd_sc_hd__clkinv_2 _13765_ (.A(_06220_),
    .Y(_06276_));
 sky130_fd_sc_hd__mux2_1 _13766_ (.A0(_06276_),
    .A1(\wfg_stim_mem_top.start_val_q[9] ),
    .S(_06262_),
    .X(_06277_));
 sky130_fd_sc_hd__mux2_1 _13767_ (.A0(net110),
    .A1(_06277_),
    .S(_06259_),
    .X(_06278_));
 sky130_fd_sc_hd__clkbuf_1 _13768_ (.A(_06278_),
    .X(_01063_));
 sky130_fd_sc_hd__clkinv_2 _13769_ (.A(_06222_),
    .Y(_06279_));
 sky130_fd_sc_hd__mux2_1 _13770_ (.A0(_06279_),
    .A1(\wfg_stim_mem_top.start_val_q[8] ),
    .S(_06262_),
    .X(_06280_));
 sky130_fd_sc_hd__mux2_1 _13771_ (.A0(net109),
    .A1(_06280_),
    .S(_06259_),
    .X(_06281_));
 sky130_fd_sc_hd__clkbuf_1 _13772_ (.A(_06281_),
    .X(_01062_));
 sky130_fd_sc_hd__clkinv_2 _13773_ (.A(_06224_),
    .Y(_06282_));
 sky130_fd_sc_hd__mux2_1 _13774_ (.A0(_06282_),
    .A1(\wfg_stim_mem_top.start_val_q[7] ),
    .S(_06255_),
    .X(_06283_));
 sky130_fd_sc_hd__mux2_1 _13775_ (.A0(net108),
    .A1(_06283_),
    .S(_06259_),
    .X(_06284_));
 sky130_fd_sc_hd__clkbuf_1 _13776_ (.A(_06284_),
    .X(_01061_));
 sky130_fd_sc_hd__clkinv_2 _13777_ (.A(_06226_),
    .Y(_06285_));
 sky130_fd_sc_hd__mux2_1 _13778_ (.A0(_06285_),
    .A1(\wfg_stim_mem_top.start_val_q[6] ),
    .S(_06255_),
    .X(_06286_));
 sky130_fd_sc_hd__mux2_1 _13779_ (.A0(net107),
    .A1(_06286_),
    .S(_06258_),
    .X(_06287_));
 sky130_fd_sc_hd__clkbuf_1 _13780_ (.A(_06287_),
    .X(_01060_));
 sky130_fd_sc_hd__clkinv_2 _13781_ (.A(_06227_),
    .Y(_06288_));
 sky130_fd_sc_hd__mux2_1 _13782_ (.A0(_06288_),
    .A1(\wfg_stim_mem_top.start_val_q[5] ),
    .S(_06255_),
    .X(_06289_));
 sky130_fd_sc_hd__mux2_1 _13783_ (.A0(net106),
    .A1(_06289_),
    .S(_06258_),
    .X(_06290_));
 sky130_fd_sc_hd__clkbuf_1 _13784_ (.A(_06290_),
    .X(_01059_));
 sky130_fd_sc_hd__clkinv_2 _13785_ (.A(_06229_),
    .Y(_06291_));
 sky130_fd_sc_hd__mux2_1 _13786_ (.A0(_06291_),
    .A1(\wfg_stim_mem_top.start_val_q[4] ),
    .S(_06255_),
    .X(_06292_));
 sky130_fd_sc_hd__mux2_1 _13787_ (.A0(net105),
    .A1(_06292_),
    .S(_06258_),
    .X(_06293_));
 sky130_fd_sc_hd__clkbuf_1 _13788_ (.A(_06293_),
    .X(_01058_));
 sky130_fd_sc_hd__clkinv_2 _13789_ (.A(_06231_),
    .Y(_06294_));
 sky130_fd_sc_hd__mux2_1 _13790_ (.A0(_06294_),
    .A1(\wfg_stim_mem_top.start_val_q[3] ),
    .S(_06255_),
    .X(_06295_));
 sky130_fd_sc_hd__mux2_1 _13791_ (.A0(net104),
    .A1(_06295_),
    .S(_06258_),
    .X(_06296_));
 sky130_fd_sc_hd__clkbuf_1 _13792_ (.A(_06296_),
    .X(_01057_));
 sky130_fd_sc_hd__clkinv_2 _13793_ (.A(_06233_),
    .Y(_06297_));
 sky130_fd_sc_hd__mux2_1 _13794_ (.A0(_06297_),
    .A1(\wfg_stim_mem_top.start_val_q[2] ),
    .S(_06255_),
    .X(_06298_));
 sky130_fd_sc_hd__mux2_1 _13795_ (.A0(net103),
    .A1(_06298_),
    .S(_06258_),
    .X(_06299_));
 sky130_fd_sc_hd__clkbuf_1 _13796_ (.A(_06299_),
    .X(_01056_));
 sky130_fd_sc_hd__inv_2 _13797_ (.A(\wfg_stim_mem_top.start_val_q[1] ),
    .Y(_06300_));
 sky130_fd_sc_hd__mux2_1 _13798_ (.A0(_06234_),
    .A1(_06300_),
    .S(_06255_),
    .X(_06301_));
 sky130_fd_sc_hd__inv_2 _13799_ (.A(_06301_),
    .Y(_06302_));
 sky130_fd_sc_hd__mux2_1 _13800_ (.A0(net102),
    .A1(_06302_),
    .S(_06258_),
    .X(_06303_));
 sky130_fd_sc_hd__clkbuf_1 _13801_ (.A(_06303_),
    .X(_01055_));
 sky130_fd_sc_hd__nand2_1 _13802_ (.A(\wfg_stim_mem_top.start_val_q[0] ),
    .B(_06262_),
    .Y(_06304_));
 sky130_fd_sc_hd__o21ai_1 _13803_ (.A1(_06236_),
    .A2(_06262_),
    .B1(_06304_),
    .Y(_06305_));
 sky130_fd_sc_hd__mux2_1 _13804_ (.A0(net101),
    .A1(_06305_),
    .S(_06258_),
    .X(_06306_));
 sky130_fd_sc_hd__clkbuf_1 _13805_ (.A(_06306_),
    .X(_01054_));
 sky130_fd_sc_hd__inv_2 _13806_ (.A(\wfg_stim_sine_top.inc_val_q[15] ),
    .Y(_06307_));
 sky130_fd_sc_hd__nand2_1 _13807_ (.A(\wfg_stim_sine_top.inc_val_q[14] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[14] ),
    .Y(_06308_));
 sky130_fd_sc_hd__or2_1 _13808_ (.A(\wfg_stim_sine_top.inc_val_q[14] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[14] ),
    .X(_06309_));
 sky130_fd_sc_hd__nand2_1 _13809_ (.A(_06308_),
    .B(_06309_),
    .Y(_06310_));
 sky130_fd_sc_hd__nor2_1 _13810_ (.A(\wfg_stim_sine_top.inc_val_q[12] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[12] ),
    .Y(_06311_));
 sky130_fd_sc_hd__nor2_1 _13811_ (.A(\wfg_stim_sine_top.inc_val_q[11] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[11] ),
    .Y(_06312_));
 sky130_fd_sc_hd__nor2_1 _13812_ (.A(\wfg_stim_sine_top.inc_val_q[10] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[10] ),
    .Y(_06313_));
 sky130_fd_sc_hd__and2_1 _13813_ (.A(\wfg_stim_sine_top.inc_val_q[9] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[9] ),
    .X(_06314_));
 sky130_fd_sc_hd__nand2_1 _13814_ (.A(\wfg_stim_sine_top.inc_val_q[8] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[8] ),
    .Y(_06315_));
 sky130_fd_sc_hd__inv_2 _13815_ (.A(_06315_),
    .Y(_06316_));
 sky130_fd_sc_hd__nor2_1 _13816_ (.A(\wfg_stim_sine_top.inc_val_q[8] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[8] ),
    .Y(_06317_));
 sky130_fd_sc_hd__nor2_1 _13817_ (.A(\wfg_stim_sine_top.inc_val_q[7] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[7] ),
    .Y(_06318_));
 sky130_fd_sc_hd__nor2_1 _13818_ (.A(\wfg_stim_sine_top.inc_val_q[6] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[6] ),
    .Y(_06319_));
 sky130_fd_sc_hd__and2_1 _13819_ (.A(\wfg_stim_sine_top.inc_val_q[5] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[5] ),
    .X(_06320_));
 sky130_fd_sc_hd__nand2_1 _13820_ (.A(\wfg_stim_sine_top.inc_val_q[4] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[4] ),
    .Y(_06321_));
 sky130_fd_sc_hd__or2_1 _13821_ (.A(\wfg_stim_sine_top.inc_val_q[4] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[4] ),
    .X(_06322_));
 sky130_fd_sc_hd__or2_1 _13822_ (.A(\wfg_stim_sine_top.inc_val_q[3] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[3] ),
    .X(_06323_));
 sky130_fd_sc_hd__nor2_1 _13823_ (.A(\wfg_stim_sine_top.inc_val_q[2] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[2] ),
    .Y(_06324_));
 sky130_fd_sc_hd__nand2_1 _13824_ (.A(\wfg_stim_sine_top.inc_val_q[0] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[0] ),
    .Y(_06325_));
 sky130_fd_sc_hd__nand2_1 _13825_ (.A(\wfg_stim_sine_top.inc_val_q[1] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[1] ),
    .Y(_06326_));
 sky130_fd_sc_hd__or2_1 _13826_ (.A(\wfg_stim_sine_top.inc_val_q[1] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[1] ),
    .X(_06327_));
 sky130_fd_sc_hd__nand2_1 _13827_ (.A(_06326_),
    .B(_06327_),
    .Y(_06328_));
 sky130_fd_sc_hd__o21a_1 _13828_ (.A1(_06325_),
    .A2(_06328_),
    .B1(_06326_),
    .X(_06329_));
 sky130_fd_sc_hd__nand2_1 _13829_ (.A(\wfg_stim_sine_top.inc_val_q[2] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[2] ),
    .Y(_06330_));
 sky130_fd_sc_hd__o21ai_1 _13830_ (.A1(_06324_),
    .A2(_06329_),
    .B1(_06330_),
    .Y(_06331_));
 sky130_fd_sc_hd__a21o_1 _13831_ (.A1(\wfg_stim_sine_top.inc_val_q[3] ),
    .A2(\wfg_stim_sine_top.wfg_stim_sine.phase_in[3] ),
    .B1(_06331_),
    .X(_06332_));
 sky130_fd_sc_hd__nand4_1 _13832_ (.A(_06321_),
    .B(_06322_),
    .C(_06323_),
    .D(_06332_),
    .Y(_06333_));
 sky130_fd_sc_hd__nor2_1 _13833_ (.A(\wfg_stim_sine_top.inc_val_q[5] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[5] ),
    .Y(_06334_));
 sky130_fd_sc_hd__or2_1 _13834_ (.A(_06320_),
    .B(_06334_),
    .X(_06335_));
 sky130_fd_sc_hd__a21oi_1 _13835_ (.A1(_06321_),
    .A2(_06333_),
    .B1(_06335_),
    .Y(_06336_));
 sky130_fd_sc_hd__nor2_1 _13836_ (.A(_06320_),
    .B(_06336_),
    .Y(_06337_));
 sky130_fd_sc_hd__nand2_1 _13837_ (.A(\wfg_stim_sine_top.inc_val_q[6] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[6] ),
    .Y(_06338_));
 sky130_fd_sc_hd__o21a_1 _13838_ (.A1(_06319_),
    .A2(_06337_),
    .B1(_06338_),
    .X(_06339_));
 sky130_fd_sc_hd__nand2_1 _13839_ (.A(\wfg_stim_sine_top.inc_val_q[7] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[7] ),
    .Y(_06340_));
 sky130_fd_sc_hd__o21a_1 _13840_ (.A1(_06318_),
    .A2(_06339_),
    .B1(_06340_),
    .X(_06341_));
 sky130_fd_sc_hd__or3_1 _13841_ (.A(_06316_),
    .B(_06317_),
    .C(_06341_),
    .X(_06342_));
 sky130_fd_sc_hd__nor2_1 _13842_ (.A(\wfg_stim_sine_top.inc_val_q[9] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[9] ),
    .Y(_06343_));
 sky130_fd_sc_hd__or2_1 _13843_ (.A(_06314_),
    .B(_06343_),
    .X(_06344_));
 sky130_fd_sc_hd__a21oi_1 _13844_ (.A1(_06315_),
    .A2(_06342_),
    .B1(_06344_),
    .Y(_06345_));
 sky130_fd_sc_hd__nor2_1 _13845_ (.A(_06314_),
    .B(_06345_),
    .Y(_06346_));
 sky130_fd_sc_hd__nand2_1 _13846_ (.A(\wfg_stim_sine_top.inc_val_q[10] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[10] ),
    .Y(_06347_));
 sky130_fd_sc_hd__o21a_1 _13847_ (.A1(_06313_),
    .A2(_06346_),
    .B1(_06347_),
    .X(_06348_));
 sky130_fd_sc_hd__nand2_1 _13848_ (.A(\wfg_stim_sine_top.inc_val_q[11] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[11] ),
    .Y(_06349_));
 sky130_fd_sc_hd__o21a_1 _13849_ (.A1(_06312_),
    .A2(_06348_),
    .B1(_06349_),
    .X(_06350_));
 sky130_fd_sc_hd__nand2_1 _13850_ (.A(\wfg_stim_sine_top.inc_val_q[12] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[12] ),
    .Y(_06351_));
 sky130_fd_sc_hd__o21ai_1 _13851_ (.A1(_06311_),
    .A2(_06350_),
    .B1(_06351_),
    .Y(_06352_));
 sky130_fd_sc_hd__a21o_1 _13852_ (.A1(\wfg_stim_sine_top.inc_val_q[13] ),
    .A2(\wfg_stim_sine_top.wfg_stim_sine.phase_in[13] ),
    .B1(_06352_),
    .X(_06353_));
 sky130_fd_sc_hd__o21a_1 _13853_ (.A1(\wfg_stim_sine_top.inc_val_q[13] ),
    .A2(\wfg_stim_sine_top.wfg_stim_sine.phase_in[13] ),
    .B1(_06353_),
    .X(_06354_));
 sky130_fd_sc_hd__or2b_1 _13854_ (.A(_06310_),
    .B_N(_06354_),
    .X(_06355_));
 sky130_fd_sc_hd__nand3b_4 _13855_ (.A_N(\wfg_stim_sine_top.wfg_stim_sine.cur_state[1] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.cur_state[0] ),
    .C(\wfg_stim_sine_top.wfg_stim_sine.cur_state[2] ),
    .Y(_06356_));
 sky130_fd_sc_hd__inv_4 _13856_ (.A(_06356_),
    .Y(_00023_));
 sky130_fd_sc_hd__or2_4 _13857_ (.A(\wfg_interconnect_top.driver1_select_q[1] ),
    .B(\wfg_interconnect_top.driver1_select_q[0] ),
    .X(_06357_));
 sky130_fd_sc_hd__nor2_1 _13858_ (.A(\wfg_interconnect_top.driver1_select_q[1] ),
    .B(\wfg_interconnect_top.driver1_select_q[0] ),
    .Y(_06358_));
 sky130_fd_sc_hd__mux2_1 _13859_ (.A0(_06358_),
    .A1(\wfg_drive_spi_top.wfg_axis_tready_o ),
    .S(_02796_),
    .X(_06359_));
 sky130_fd_sc_hd__o21a_4 _13860_ (.A1(\wfg_drive_pat_top.wfg_axis_tready_o ),
    .A2(_06357_),
    .B1(_06359_),
    .X(_06360_));
 sky130_fd_sc_hd__nand2_4 _13861_ (.A(_00023_),
    .B(_06360_),
    .Y(_06361_));
 sky130_fd_sc_hd__a21oi_1 _13862_ (.A1(_06308_),
    .A2(_06355_),
    .B1(_06307_),
    .Y(_06362_));
 sky130_fd_sc_hd__a311oi_2 _13863_ (.A1(_06307_),
    .A2(_06308_),
    .A3(_06355_),
    .B1(_06361_),
    .C1(_06362_),
    .Y(_06363_));
 sky130_fd_sc_hd__xor2_1 _13864_ (.A(\wfg_stim_sine_top.wfg_stim_sine.phase_in[15] ),
    .B(_06363_),
    .X(_00977_));
 sky130_fd_sc_hd__xnor2_1 _13865_ (.A(_06310_),
    .B(_06354_),
    .Y(_06364_));
 sky130_fd_sc_hd__clkbuf_4 _13866_ (.A(_06361_),
    .X(_06365_));
 sky130_fd_sc_hd__mux2_1 _13867_ (.A0(_06364_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.phase_in[14] ),
    .S(_06365_),
    .X(_06366_));
 sky130_fd_sc_hd__clkbuf_1 _13868_ (.A(_06366_),
    .X(_00976_));
 sky130_fd_sc_hd__xnor2_1 _13869_ (.A(\wfg_stim_sine_top.inc_val_q[13] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[13] ),
    .Y(_06367_));
 sky130_fd_sc_hd__xnor2_1 _13870_ (.A(_06352_),
    .B(_06367_),
    .Y(_06368_));
 sky130_fd_sc_hd__mux2_1 _13871_ (.A0(_06368_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.phase_in[13] ),
    .S(_06365_),
    .X(_06369_));
 sky130_fd_sc_hd__clkbuf_1 _13872_ (.A(_06369_),
    .X(_00975_));
 sky130_fd_sc_hd__or2b_1 _13873_ (.A(_06311_),
    .B_N(_06351_),
    .X(_06370_));
 sky130_fd_sc_hd__xor2_1 _13874_ (.A(_06350_),
    .B(_06370_),
    .X(_06371_));
 sky130_fd_sc_hd__mux2_1 _13875_ (.A0(_06371_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.phase_in[12] ),
    .S(_06365_),
    .X(_06372_));
 sky130_fd_sc_hd__clkbuf_1 _13876_ (.A(_06372_),
    .X(_00974_));
 sky130_fd_sc_hd__and2b_1 _13877_ (.A_N(_06312_),
    .B(_06349_),
    .X(_06373_));
 sky130_fd_sc_hd__xnor2_1 _13878_ (.A(_06348_),
    .B(_06373_),
    .Y(_06374_));
 sky130_fd_sc_hd__mux2_1 _13879_ (.A0(_06374_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.phase_in[11] ),
    .S(_06365_),
    .X(_06375_));
 sky130_fd_sc_hd__clkbuf_1 _13880_ (.A(_06375_),
    .X(_00973_));
 sky130_fd_sc_hd__and2b_1 _13881_ (.A_N(_06313_),
    .B(_06347_),
    .X(_06376_));
 sky130_fd_sc_hd__xnor2_1 _13882_ (.A(_06346_),
    .B(_06376_),
    .Y(_06377_));
 sky130_fd_sc_hd__mux2_1 _13883_ (.A0(_06377_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.phase_in[10] ),
    .S(_06361_),
    .X(_06378_));
 sky130_fd_sc_hd__clkbuf_1 _13884_ (.A(_06378_),
    .X(_00972_));
 sky130_fd_sc_hd__a31o_1 _13885_ (.A1(_06344_),
    .A2(_06315_),
    .A3(_06342_),
    .B1(_06365_),
    .X(_06379_));
 sky130_fd_sc_hd__a2bb2o_1 _13886_ (.A1_N(_06345_),
    .A2_N(_06379_),
    .B1(_06365_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.phase_in[9] ),
    .X(_00971_));
 sky130_fd_sc_hd__o21a_1 _13887_ (.A1(_06316_),
    .A2(_06317_),
    .B1(_06341_),
    .X(_06380_));
 sky130_fd_sc_hd__nor2_1 _13888_ (.A(_06365_),
    .B(_06380_),
    .Y(_06381_));
 sky130_fd_sc_hd__a22o_1 _13889_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.phase_in[8] ),
    .A2(_06365_),
    .B1(_06381_),
    .B2(_06342_),
    .X(_00970_));
 sky130_fd_sc_hd__and2b_1 _13890_ (.A_N(_06318_),
    .B(_06340_),
    .X(_06382_));
 sky130_fd_sc_hd__xnor2_1 _13891_ (.A(_06339_),
    .B(_06382_),
    .Y(_06383_));
 sky130_fd_sc_hd__mux2_1 _13892_ (.A0(_06383_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.phase_in[7] ),
    .S(_06361_),
    .X(_06384_));
 sky130_fd_sc_hd__clkbuf_1 _13893_ (.A(_06384_),
    .X(_00969_));
 sky130_fd_sc_hd__or2b_1 _13894_ (.A(_06319_),
    .B_N(_06338_),
    .X(_06385_));
 sky130_fd_sc_hd__xor2_1 _13895_ (.A(_06337_),
    .B(_06385_),
    .X(_06386_));
 sky130_fd_sc_hd__mux2_1 _13896_ (.A0(_06386_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.phase_in[6] ),
    .S(_06361_),
    .X(_06387_));
 sky130_fd_sc_hd__clkbuf_1 _13897_ (.A(_06387_),
    .X(_00968_));
 sky130_fd_sc_hd__a31o_1 _13898_ (.A1(_06335_),
    .A2(_06321_),
    .A3(_06333_),
    .B1(_06365_),
    .X(_06388_));
 sky130_fd_sc_hd__a2bb2o_1 _13899_ (.A1_N(_06336_),
    .A2_N(_06388_),
    .B1(_06365_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.phase_in[5] ),
    .X(_00967_));
 sky130_fd_sc_hd__a22o_1 _13900_ (.A1(_06321_),
    .A2(_06322_),
    .B1(_06323_),
    .B2(_06332_),
    .X(_06389_));
 sky130_fd_sc_hd__and2_1 _13901_ (.A(\wfg_stim_sine_top.wfg_stim_sine.phase_in[4] ),
    .B(_06361_),
    .X(_06390_));
 sky130_fd_sc_hd__a41o_1 _13902_ (.A1(_06333_),
    .A2(_00023_),
    .A3(_06360_),
    .A4(_06389_),
    .B1(_06390_),
    .X(_00966_));
 sky130_fd_sc_hd__nand2_1 _13903_ (.A(\wfg_stim_sine_top.inc_val_q[3] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.phase_in[3] ),
    .Y(_06391_));
 sky130_fd_sc_hd__and3_1 _13904_ (.A(_06323_),
    .B(_06391_),
    .C(_06331_),
    .X(_06392_));
 sky130_fd_sc_hd__a21oi_1 _13905_ (.A1(_06323_),
    .A2(_06391_),
    .B1(_06331_),
    .Y(_06393_));
 sky130_fd_sc_hd__nor2_1 _13906_ (.A(_06392_),
    .B(_06393_),
    .Y(_06394_));
 sky130_fd_sc_hd__mux2_1 _13907_ (.A0(_06394_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.phase_in[3] ),
    .S(_06361_),
    .X(_06395_));
 sky130_fd_sc_hd__clkbuf_1 _13908_ (.A(_06395_),
    .X(_00965_));
 sky130_fd_sc_hd__or2b_1 _13909_ (.A(_06324_),
    .B_N(_06330_),
    .X(_06396_));
 sky130_fd_sc_hd__xor2_1 _13910_ (.A(_06329_),
    .B(_06396_),
    .X(_06397_));
 sky130_fd_sc_hd__mux2_1 _13911_ (.A0(_06397_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.phase_in[2] ),
    .S(_06361_),
    .X(_06398_));
 sky130_fd_sc_hd__clkbuf_1 _13912_ (.A(_06398_),
    .X(_00964_));
 sky130_fd_sc_hd__xor2_1 _13913_ (.A(_06325_),
    .B(_06328_),
    .X(_06399_));
 sky130_fd_sc_hd__mux2_1 _13914_ (.A0(_06399_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.phase_in[1] ),
    .S(_06361_),
    .X(_06400_));
 sky130_fd_sc_hd__clkbuf_1 _13915_ (.A(_06400_),
    .X(_00963_));
 sky130_fd_sc_hd__nand3_1 _13916_ (.A(\wfg_stim_sine_top.inc_val_q[0] ),
    .B(_00023_),
    .C(_06360_),
    .Y(_06401_));
 sky130_fd_sc_hd__xnor2_1 _13917_ (.A(\wfg_stim_sine_top.wfg_stim_sine.phase_in[0] ),
    .B(_06401_),
    .Y(_00962_));
 sky130_fd_sc_hd__and3b_1 _13918_ (.A_N(\wfg_stim_sine_top.wfg_stim_sine.cur_state[2] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.cur_state[1] ),
    .C(\wfg_stim_sine_top.wfg_stim_sine.cur_state[0] ),
    .X(_06402_));
 sky130_fd_sc_hd__buf_2 _13919_ (.A(_06402_),
    .X(_06403_));
 sky130_fd_sc_hd__clkbuf_8 _13920_ (.A(_06403_),
    .X(_06404_));
 sky130_fd_sc_hd__buf_2 _13921_ (.A(\wfg_stim_sine_top.gain_val_q[15] ),
    .X(_06405_));
 sky130_fd_sc_hd__buf_4 _13922_ (.A(_06405_),
    .X(_06406_));
 sky130_fd_sc_hd__inv_6 _13923_ (.A(_06406_),
    .Y(_06407_));
 sky130_fd_sc_hd__buf_6 _13924_ (.A(_06407_),
    .X(_06408_));
 sky130_fd_sc_hd__buf_4 _13925_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[16] ),
    .X(_06409_));
 sky130_fd_sc_hd__inv_4 _13926_ (.A(_06409_),
    .Y(_06410_));
 sky130_fd_sc_hd__o21ai_1 _13927_ (.A1(_06408_),
    .A2(_06410_),
    .B1(_06404_),
    .Y(_06411_));
 sky130_fd_sc_hd__clkbuf_4 _13928_ (.A(\wfg_stim_sine_top.gain_val_q[14] ),
    .X(_06412_));
 sky130_fd_sc_hd__clkbuf_8 _13929_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[11] ),
    .X(_06413_));
 sky130_fd_sc_hd__buf_4 _13930_ (.A(_06413_),
    .X(_06414_));
 sky130_fd_sc_hd__buf_4 _13931_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[10] ),
    .X(_06415_));
 sky130_fd_sc_hd__buf_2 _13932_ (.A(_06415_),
    .X(_06416_));
 sky130_fd_sc_hd__and4_1 _13933_ (.A(_06405_),
    .B(_06412_),
    .C(_06414_),
    .D(_06416_),
    .X(_06417_));
 sky130_fd_sc_hd__a22oi_1 _13934_ (.A1(_06412_),
    .A2(_06414_),
    .B1(_06416_),
    .B2(_06405_),
    .Y(_06418_));
 sky130_fd_sc_hd__buf_2 _13935_ (.A(\wfg_stim_sine_top.gain_val_q[13] ),
    .X(_06419_));
 sky130_fd_sc_hd__clkbuf_4 _13936_ (.A(_06419_),
    .X(_06420_));
 sky130_fd_sc_hd__clkbuf_8 _13937_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[12] ),
    .X(_06421_));
 sky130_fd_sc_hd__buf_4 _13938_ (.A(_06421_),
    .X(_06422_));
 sky130_fd_sc_hd__buf_6 _13939_ (.A(_06422_),
    .X(_06423_));
 sky130_fd_sc_hd__and4bb_1 _13940_ (.A_N(_06417_),
    .B_N(_06418_),
    .C(_06420_),
    .D(_06423_),
    .X(_06424_));
 sky130_fd_sc_hd__o2bb2a_1 _13941_ (.A1_N(_06420_),
    .A2_N(_06423_),
    .B1(_06417_),
    .B2(_06418_),
    .X(_06425_));
 sky130_fd_sc_hd__buf_6 _13942_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[9] ),
    .X(_06426_));
 sky130_fd_sc_hd__buf_4 _13943_ (.A(_06426_),
    .X(_06427_));
 sky130_fd_sc_hd__clkbuf_8 _13944_ (.A(_06427_),
    .X(_06428_));
 sky130_fd_sc_hd__and4_1 _13945_ (.A(_06405_),
    .B(_06412_),
    .C(_06416_),
    .D(_06428_),
    .X(_06429_));
 sky130_fd_sc_hd__buf_6 _13946_ (.A(_06428_),
    .X(_06430_));
 sky130_fd_sc_hd__a22oi_1 _13947_ (.A1(_06412_),
    .A2(_06416_),
    .B1(_06430_),
    .B2(_06405_),
    .Y(_06431_));
 sky130_fd_sc_hd__buf_6 _13948_ (.A(_06414_),
    .X(_06432_));
 sky130_fd_sc_hd__and4bb_1 _13949_ (.A_N(_06429_),
    .B_N(_06431_),
    .C(_06420_),
    .D(_06432_),
    .X(_06433_));
 sky130_fd_sc_hd__nor2_1 _13950_ (.A(_06429_),
    .B(_06433_),
    .Y(_06434_));
 sky130_fd_sc_hd__or3_1 _13951_ (.A(_06424_),
    .B(_06425_),
    .C(_06434_),
    .X(_06435_));
 sky130_fd_sc_hd__nor2_1 _13952_ (.A(_06424_),
    .B(_06425_),
    .Y(_06436_));
 sky130_fd_sc_hd__xnor2_1 _13953_ (.A(_06436_),
    .B(_06434_),
    .Y(_06437_));
 sky130_fd_sc_hd__buf_2 _13954_ (.A(\wfg_stim_sine_top.gain_val_q[11] ),
    .X(_06438_));
 sky130_fd_sc_hd__clkbuf_4 _13955_ (.A(_06438_),
    .X(_06439_));
 sky130_fd_sc_hd__clkbuf_4 _13956_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[14] ),
    .X(_06440_));
 sky130_fd_sc_hd__clkbuf_4 _13957_ (.A(_06440_),
    .X(_06441_));
 sky130_fd_sc_hd__buf_4 _13958_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[13] ),
    .X(_06442_));
 sky130_fd_sc_hd__buf_4 _13959_ (.A(_06442_),
    .X(_06443_));
 sky130_fd_sc_hd__clkbuf_4 _13960_ (.A(\wfg_stim_sine_top.gain_val_q[12] ),
    .X(_06444_));
 sky130_fd_sc_hd__a22oi_1 _13961_ (.A1(_06439_),
    .A2(_06441_),
    .B1(_06443_),
    .B2(_06444_),
    .Y(_06445_));
 sky130_fd_sc_hd__buf_2 _13962_ (.A(\wfg_stim_sine_top.gain_val_q[12] ),
    .X(_06446_));
 sky130_fd_sc_hd__buf_2 _13963_ (.A(_06438_),
    .X(_06447_));
 sky130_fd_sc_hd__and4_1 _13964_ (.A(_06446_),
    .B(_06447_),
    .C(_06440_),
    .D(_06442_),
    .X(_06448_));
 sky130_fd_sc_hd__nor2_1 _13965_ (.A(_06445_),
    .B(_06448_),
    .Y(_06449_));
 sky130_fd_sc_hd__clkbuf_4 _13966_ (.A(\wfg_stim_sine_top.gain_val_q[10] ),
    .X(_06450_));
 sky130_fd_sc_hd__clkbuf_8 _13967_ (.A(_06450_),
    .X(_06451_));
 sky130_fd_sc_hd__buf_4 _13968_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[15] ),
    .X(_06452_));
 sky130_fd_sc_hd__buf_4 _13969_ (.A(_06452_),
    .X(_06453_));
 sky130_fd_sc_hd__buf_4 _13970_ (.A(_06453_),
    .X(_06454_));
 sky130_fd_sc_hd__nand2_1 _13971_ (.A(_06451_),
    .B(_06454_),
    .Y(_06455_));
 sky130_fd_sc_hd__xnor2_1 _13972_ (.A(_06449_),
    .B(_06455_),
    .Y(_06456_));
 sky130_fd_sc_hd__nand2_1 _13973_ (.A(_06437_),
    .B(_06456_),
    .Y(_06457_));
 sky130_fd_sc_hd__buf_2 _13974_ (.A(\wfg_stim_sine_top.gain_val_q[15] ),
    .X(_06458_));
 sky130_fd_sc_hd__buf_2 _13975_ (.A(\wfg_stim_sine_top.gain_val_q[14] ),
    .X(_06459_));
 sky130_fd_sc_hd__and4_1 _13976_ (.A(_06458_),
    .B(_06459_),
    .C(_06421_),
    .D(_06413_),
    .X(_06460_));
 sky130_fd_sc_hd__a22o_1 _13977_ (.A1(_06412_),
    .A2(_06421_),
    .B1(_06413_),
    .B2(_06405_),
    .X(_06461_));
 sky130_fd_sc_hd__and2b_1 _13978_ (.A_N(_06460_),
    .B(_06461_),
    .X(_06462_));
 sky130_fd_sc_hd__buf_4 _13979_ (.A(_06443_),
    .X(_06463_));
 sky130_fd_sc_hd__nand2_1 _13980_ (.A(_06420_),
    .B(_06463_),
    .Y(_06464_));
 sky130_fd_sc_hd__xnor2_1 _13981_ (.A(_06462_),
    .B(_06464_),
    .Y(_06465_));
 sky130_fd_sc_hd__nor2_1 _13982_ (.A(_06417_),
    .B(_06424_),
    .Y(_06466_));
 sky130_fd_sc_hd__xnor2_1 _13983_ (.A(_06465_),
    .B(_06466_),
    .Y(_06467_));
 sky130_fd_sc_hd__buf_4 _13984_ (.A(_06450_),
    .X(_06468_));
 sky130_fd_sc_hd__buf_4 _13985_ (.A(_06409_),
    .X(_06469_));
 sky130_fd_sc_hd__nand2_4 _13986_ (.A(_06468_),
    .B(_06469_),
    .Y(_06470_));
 sky130_fd_sc_hd__buf_4 _13987_ (.A(_06439_),
    .X(_06471_));
 sky130_fd_sc_hd__buf_6 _13988_ (.A(_06453_),
    .X(_06472_));
 sky130_fd_sc_hd__clkbuf_4 _13989_ (.A(_06441_),
    .X(_06473_));
 sky130_fd_sc_hd__buf_4 _13990_ (.A(_06444_),
    .X(_06474_));
 sky130_fd_sc_hd__a22oi_1 _13991_ (.A1(_06471_),
    .A2(_06472_),
    .B1(_06473_),
    .B2(_06474_),
    .Y(_06475_));
 sky130_fd_sc_hd__and4_1 _13992_ (.A(_06444_),
    .B(_06471_),
    .C(_06453_),
    .D(_06473_),
    .X(_06476_));
 sky130_fd_sc_hd__nor2_1 _13993_ (.A(_06475_),
    .B(_06476_),
    .Y(_06477_));
 sky130_fd_sc_hd__xnor2_1 _13994_ (.A(_06470_),
    .B(_06477_),
    .Y(_06478_));
 sky130_fd_sc_hd__nand2_1 _13995_ (.A(_06467_),
    .B(_06478_),
    .Y(_06479_));
 sky130_fd_sc_hd__or2_1 _13996_ (.A(_06467_),
    .B(_06478_),
    .X(_06480_));
 sky130_fd_sc_hd__nand2_1 _13997_ (.A(_06479_),
    .B(_06480_),
    .Y(_06481_));
 sky130_fd_sc_hd__a21o_1 _13998_ (.A1(_06435_),
    .A2(_06457_),
    .B1(_06481_),
    .X(_06482_));
 sky130_fd_sc_hd__nand3_1 _13999_ (.A(_06481_),
    .B(_06435_),
    .C(_06457_),
    .Y(_06483_));
 sky130_fd_sc_hd__buf_2 _14000_ (.A(\wfg_stim_sine_top.gain_val_q[7] ),
    .X(_06484_));
 sky130_fd_sc_hd__buf_4 _14001_ (.A(_06484_),
    .X(_06485_));
 sky130_fd_sc_hd__buf_6 _14002_ (.A(_06485_),
    .X(_06486_));
 sky130_fd_sc_hd__clkbuf_4 _14003_ (.A(\wfg_stim_sine_top.gain_val_q[9] ),
    .X(_06487_));
 sky130_fd_sc_hd__clkbuf_4 _14004_ (.A(\wfg_stim_sine_top.gain_val_q[8] ),
    .X(_06488_));
 sky130_fd_sc_hd__and3_2 _14005_ (.A(_06487_),
    .B(_06488_),
    .C(_06409_),
    .X(_06489_));
 sky130_fd_sc_hd__clkbuf_4 _14006_ (.A(\wfg_stim_sine_top.gain_val_q[8] ),
    .X(_06490_));
 sky130_fd_sc_hd__o21ai_2 _14007_ (.A1(_06487_),
    .A2(_06490_),
    .B1(_06409_),
    .Y(_06491_));
 sky130_fd_sc_hd__nor2_4 _14008_ (.A(_06489_),
    .B(_06491_),
    .Y(_06492_));
 sky130_fd_sc_hd__a21oi_4 _14009_ (.A1(_06486_),
    .A2(_06492_),
    .B1(_06489_),
    .Y(_06493_));
 sky130_fd_sc_hd__nand2_2 _14010_ (.A(_06485_),
    .B(_06469_),
    .Y(_06494_));
 sky130_fd_sc_hd__xnor2_4 _14011_ (.A(_06492_),
    .B(_06494_),
    .Y(_06495_));
 sky130_fd_sc_hd__a31o_1 _14012_ (.A1(_06468_),
    .A2(_06472_),
    .A3(_06449_),
    .B1(_06448_),
    .X(_06496_));
 sky130_fd_sc_hd__nand2_1 _14013_ (.A(_06495_),
    .B(_06496_),
    .Y(_06497_));
 sky130_fd_sc_hd__or2_1 _14014_ (.A(_06495_),
    .B(_06496_),
    .X(_06498_));
 sky130_fd_sc_hd__nand2_1 _14015_ (.A(_06497_),
    .B(_06498_),
    .Y(_06499_));
 sky130_fd_sc_hd__or2_1 _14016_ (.A(_06493_),
    .B(_06499_),
    .X(_06500_));
 sky130_fd_sc_hd__nand2_1 _14017_ (.A(_06493_),
    .B(_06499_),
    .Y(_06501_));
 sky130_fd_sc_hd__and2_1 _14018_ (.A(_06500_),
    .B(_06501_),
    .X(_06502_));
 sky130_fd_sc_hd__nand3_1 _14019_ (.A(_06482_),
    .B(_06483_),
    .C(_06502_),
    .Y(_06503_));
 sky130_fd_sc_hd__or2b_1 _14020_ (.A(_06466_),
    .B_N(_06465_),
    .X(_06504_));
 sky130_fd_sc_hd__buf_4 _14021_ (.A(_06412_),
    .X(_06505_));
 sky130_fd_sc_hd__and4_1 _14022_ (.A(_06405_),
    .B(_06505_),
    .C(_06443_),
    .D(_06422_),
    .X(_06506_));
 sky130_fd_sc_hd__a22oi_1 _14023_ (.A1(_06505_),
    .A2(_06463_),
    .B1(_06423_),
    .B2(_06406_),
    .Y(_06507_));
 sky130_fd_sc_hd__and4bb_1 _14024_ (.A_N(_06506_),
    .B_N(_06507_),
    .C(_06420_),
    .D(_06473_),
    .X(_06508_));
 sky130_fd_sc_hd__clkbuf_8 _14025_ (.A(_06420_),
    .X(_06509_));
 sky130_fd_sc_hd__clkbuf_8 _14026_ (.A(_06473_),
    .X(_06510_));
 sky130_fd_sc_hd__o2bb2a_1 _14027_ (.A1_N(_06509_),
    .A2_N(_06510_),
    .B1(_06506_),
    .B2(_06507_),
    .X(_06511_));
 sky130_fd_sc_hd__nor2_1 _14028_ (.A(_06508_),
    .B(_06511_),
    .Y(_06512_));
 sky130_fd_sc_hd__buf_4 _14029_ (.A(_06463_),
    .X(_06513_));
 sky130_fd_sc_hd__a31o_1 _14030_ (.A1(_06509_),
    .A2(_06513_),
    .A3(_06461_),
    .B1(_06460_),
    .X(_06514_));
 sky130_fd_sc_hd__xor2_1 _14031_ (.A(_06512_),
    .B(_06514_),
    .X(_06515_));
 sky130_fd_sc_hd__and3_1 _14032_ (.A(_06471_),
    .B(_06469_),
    .C(_06472_),
    .X(_06516_));
 sky130_fd_sc_hd__a22o_1 _14033_ (.A1(_06471_),
    .A2(_06469_),
    .B1(_06472_),
    .B2(_06474_),
    .X(_06517_));
 sky130_fd_sc_hd__a21bo_1 _14034_ (.A1(_06474_),
    .A2(_06516_),
    .B1_N(_06517_),
    .X(_06518_));
 sky130_fd_sc_hd__xor2_1 _14035_ (.A(_06470_),
    .B(_06518_),
    .X(_06519_));
 sky130_fd_sc_hd__and2_1 _14036_ (.A(_06515_),
    .B(_06519_),
    .X(_06520_));
 sky130_fd_sc_hd__nor2_1 _14037_ (.A(_06515_),
    .B(_06519_),
    .Y(_06521_));
 sky130_fd_sc_hd__or2_1 _14038_ (.A(_06520_),
    .B(_06521_),
    .X(_06522_));
 sky130_fd_sc_hd__a21o_1 _14039_ (.A1(_06504_),
    .A2(_06479_),
    .B1(_06522_),
    .X(_06523_));
 sky130_fd_sc_hd__nand3_1 _14040_ (.A(_06522_),
    .B(_06504_),
    .C(_06479_),
    .Y(_06524_));
 sky130_fd_sc_hd__buf_4 _14041_ (.A(_06469_),
    .X(_06525_));
 sky130_fd_sc_hd__a31o_1 _14042_ (.A1(_06451_),
    .A2(_06525_),
    .A3(_06477_),
    .B1(_06476_),
    .X(_06526_));
 sky130_fd_sc_hd__xnor2_1 _14043_ (.A(_06495_),
    .B(_06526_),
    .Y(_06527_));
 sky130_fd_sc_hd__or2_1 _14044_ (.A(_06493_),
    .B(_06527_),
    .X(_06528_));
 sky130_fd_sc_hd__nand2_1 _14045_ (.A(_06493_),
    .B(_06527_),
    .Y(_06529_));
 sky130_fd_sc_hd__and2_1 _14046_ (.A(_06528_),
    .B(_06529_),
    .X(_06530_));
 sky130_fd_sc_hd__and3_1 _14047_ (.A(_06523_),
    .B(_06524_),
    .C(_06530_),
    .X(_06531_));
 sky130_fd_sc_hd__a21oi_1 _14048_ (.A1(_06523_),
    .A2(_06524_),
    .B1(_06530_),
    .Y(_06532_));
 sky130_fd_sc_hd__a211oi_2 _14049_ (.A1(_06482_),
    .A2(_06503_),
    .B1(_06531_),
    .C1(_06532_),
    .Y(_06533_));
 sky130_fd_sc_hd__inv_2 _14050_ (.A(_06533_),
    .Y(_06534_));
 sky130_fd_sc_hd__o211a_1 _14051_ (.A1(_06531_),
    .A2(_06532_),
    .B1(_06482_),
    .C1(_06503_),
    .X(_06535_));
 sky130_fd_sc_hd__and3_1 _14052_ (.A(\wfg_stim_sine_top.gain_val_q[1] ),
    .B(\wfg_stim_sine_top.gain_val_q[0] ),
    .C(\wfg_stim_sine_top.wfg_stim_sine.sin_17[16] ),
    .X(_06536_));
 sky130_fd_sc_hd__buf_2 _14053_ (.A(_06536_),
    .X(_06537_));
 sky130_fd_sc_hd__clkbuf_4 _14054_ (.A(\wfg_stim_sine_top.gain_val_q[1] ),
    .X(_06538_));
 sky130_fd_sc_hd__clkbuf_4 _14055_ (.A(\wfg_stim_sine_top.gain_val_q[0] ),
    .X(_06539_));
 sky130_fd_sc_hd__o21ai_2 _14056_ (.A1(_06538_),
    .A2(_06539_),
    .B1(_06409_),
    .Y(_06540_));
 sky130_fd_sc_hd__nor2_8 _14057_ (.A(_06537_),
    .B(_06540_),
    .Y(_06541_));
 sky130_fd_sc_hd__nand2_4 _14058_ (.A(\wfg_stim_sine_top.gain_val_q[2] ),
    .B(_06469_),
    .Y(_06542_));
 sky130_fd_sc_hd__xor2_4 _14059_ (.A(_06541_),
    .B(_06542_),
    .X(_06543_));
 sky130_fd_sc_hd__clkbuf_4 _14060_ (.A(\wfg_stim_sine_top.gain_val_q[4] ),
    .X(_06544_));
 sky130_fd_sc_hd__nand2_2 _14061_ (.A(_06544_),
    .B(_06409_),
    .Y(_06545_));
 sky130_fd_sc_hd__clkbuf_4 _14062_ (.A(\wfg_stim_sine_top.gain_val_q[6] ),
    .X(_06546_));
 sky130_fd_sc_hd__buf_4 _14063_ (.A(_06546_),
    .X(_06547_));
 sky130_fd_sc_hd__clkbuf_4 _14064_ (.A(\wfg_stim_sine_top.gain_val_q[5] ),
    .X(_06548_));
 sky130_fd_sc_hd__buf_4 _14065_ (.A(_06548_),
    .X(_06549_));
 sky130_fd_sc_hd__o21ai_1 _14066_ (.A1(_06547_),
    .A2(_06549_),
    .B1(_06469_),
    .Y(_06550_));
 sky130_fd_sc_hd__buf_4 _14067_ (.A(_06544_),
    .X(_06551_));
 sky130_fd_sc_hd__and3_1 _14068_ (.A(_06547_),
    .B(_06549_),
    .C(_06409_),
    .X(_06552_));
 sky130_fd_sc_hd__and2_1 _14069_ (.A(_06551_),
    .B(_06552_),
    .X(_06553_));
 sky130_fd_sc_hd__a21o_4 _14070_ (.A1(_06545_),
    .A2(_06550_),
    .B1(_06553_),
    .X(_06554_));
 sky130_fd_sc_hd__o21bai_4 _14071_ (.A1(_06543_),
    .A2(_06554_),
    .B1_N(_06553_),
    .Y(_06555_));
 sky130_fd_sc_hd__buf_4 _14072_ (.A(_06555_),
    .X(_06556_));
 sky130_fd_sc_hd__xnor2_4 _14073_ (.A(_06543_),
    .B(_06554_),
    .Y(_06557_));
 sky130_fd_sc_hd__a21oi_1 _14074_ (.A1(_06497_),
    .A2(_06500_),
    .B1(_06557_),
    .Y(_06558_));
 sky130_fd_sc_hd__and3_1 _14075_ (.A(_06557_),
    .B(_06497_),
    .C(_06500_),
    .X(_06559_));
 sky130_fd_sc_hd__nor2_1 _14076_ (.A(_06558_),
    .B(_06559_),
    .Y(_06560_));
 sky130_fd_sc_hd__xnor2_1 _14077_ (.A(_06556_),
    .B(_06560_),
    .Y(_06561_));
 sky130_fd_sc_hd__or3_2 _14078_ (.A(_06533_),
    .B(_06535_),
    .C(_06561_),
    .X(_06562_));
 sky130_fd_sc_hd__a21oi_1 _14079_ (.A1(_06504_),
    .A2(_06479_),
    .B1(_06522_),
    .Y(_06563_));
 sky130_fd_sc_hd__and2_1 _14080_ (.A(_06512_),
    .B(_06514_),
    .X(_06564_));
 sky130_fd_sc_hd__and3_1 _14081_ (.A(_06474_),
    .B(_06471_),
    .C(_06469_),
    .X(_06565_));
 sky130_fd_sc_hd__o21ai_1 _14082_ (.A1(_06474_),
    .A2(_06471_),
    .B1(_06525_),
    .Y(_06566_));
 sky130_fd_sc_hd__nor2_2 _14083_ (.A(_06565_),
    .B(_06566_),
    .Y(_06567_));
 sky130_fd_sc_hd__xnor2_4 _14084_ (.A(_06470_),
    .B(_06567_),
    .Y(_06568_));
 sky130_fd_sc_hd__and4_1 _14085_ (.A(_06406_),
    .B(_06505_),
    .C(_06441_),
    .D(_06443_),
    .X(_06569_));
 sky130_fd_sc_hd__a22oi_1 _14086_ (.A1(_06505_),
    .A2(_06473_),
    .B1(_06463_),
    .B2(_06406_),
    .Y(_06570_));
 sky130_fd_sc_hd__and4bb_1 _14087_ (.A_N(_06569_),
    .B_N(_06570_),
    .C(_06509_),
    .D(_06454_),
    .X(_06571_));
 sky130_fd_sc_hd__o2bb2a_1 _14088_ (.A1_N(_06509_),
    .A2_N(_06454_),
    .B1(_06569_),
    .B2(_06570_),
    .X(_06572_));
 sky130_fd_sc_hd__nor2_1 _14089_ (.A(_06571_),
    .B(_06572_),
    .Y(_06573_));
 sky130_fd_sc_hd__nor2_1 _14090_ (.A(_06506_),
    .B(_06508_),
    .Y(_06574_));
 sky130_fd_sc_hd__xnor2_1 _14091_ (.A(_06573_),
    .B(_06574_),
    .Y(_06575_));
 sky130_fd_sc_hd__xor2_1 _14092_ (.A(_06568_),
    .B(_06575_),
    .X(_06576_));
 sky130_fd_sc_hd__o21ai_2 _14093_ (.A1(_06564_),
    .A2(_06520_),
    .B1(_06576_),
    .Y(_06577_));
 sky130_fd_sc_hd__or3_1 _14094_ (.A(_06576_),
    .B(_06564_),
    .C(_06520_),
    .X(_06578_));
 sky130_fd_sc_hd__nand2_1 _14095_ (.A(_06577_),
    .B(_06578_),
    .Y(_06579_));
 sky130_fd_sc_hd__and2_1 _14096_ (.A(_06474_),
    .B(_06516_),
    .X(_06580_));
 sky130_fd_sc_hd__a31o_1 _14097_ (.A1(_06451_),
    .A2(_06525_),
    .A3(_06517_),
    .B1(_06580_),
    .X(_06581_));
 sky130_fd_sc_hd__nand2_1 _14098_ (.A(_06495_),
    .B(_06581_),
    .Y(_06582_));
 sky130_fd_sc_hd__or2_1 _14099_ (.A(_06495_),
    .B(_06581_),
    .X(_06583_));
 sky130_fd_sc_hd__nand2_1 _14100_ (.A(_06582_),
    .B(_06583_),
    .Y(_06584_));
 sky130_fd_sc_hd__or2_1 _14101_ (.A(_06493_),
    .B(_06584_),
    .X(_06585_));
 sky130_fd_sc_hd__nand2_1 _14102_ (.A(_06493_),
    .B(_06584_),
    .Y(_06586_));
 sky130_fd_sc_hd__nand2_1 _14103_ (.A(_06585_),
    .B(_06586_),
    .Y(_06587_));
 sky130_fd_sc_hd__xor2_1 _14104_ (.A(_06579_),
    .B(_06587_),
    .X(_06588_));
 sky130_fd_sc_hd__o21a_1 _14105_ (.A1(_06563_),
    .A2(_06531_),
    .B1(_06588_),
    .X(_06589_));
 sky130_fd_sc_hd__nor3_1 _14106_ (.A(_06588_),
    .B(_06563_),
    .C(_06531_),
    .Y(_06590_));
 sky130_fd_sc_hd__a21bo_1 _14107_ (.A1(_06495_),
    .A2(_06526_),
    .B1_N(_06528_),
    .X(_06591_));
 sky130_fd_sc_hd__xnor2_1 _14108_ (.A(_06557_),
    .B(_06591_),
    .Y(_06592_));
 sky130_fd_sc_hd__xnor2_1 _14109_ (.A(_06556_),
    .B(_06592_),
    .Y(_06593_));
 sky130_fd_sc_hd__nor3_1 _14110_ (.A(_06589_),
    .B(_06590_),
    .C(_06593_),
    .Y(_06594_));
 sky130_fd_sc_hd__o21a_1 _14111_ (.A1(_06589_),
    .A2(_06590_),
    .B1(_06593_),
    .X(_06595_));
 sky130_fd_sc_hd__or2_1 _14112_ (.A(_06594_),
    .B(_06595_),
    .X(_06596_));
 sky130_fd_sc_hd__a21oi_2 _14113_ (.A1(_06534_),
    .A2(_06562_),
    .B1(_06596_),
    .Y(_06597_));
 sky130_fd_sc_hd__and3_1 _14114_ (.A(_06596_),
    .B(_06534_),
    .C(_06562_),
    .X(_06598_));
 sky130_fd_sc_hd__buf_8 _14115_ (.A(\wfg_stim_sine_top.gain_val_q[3] ),
    .X(_06599_));
 sky130_fd_sc_hd__buf_6 _14116_ (.A(_06525_),
    .X(_06600_));
 sky130_fd_sc_hd__nand2_8 _14117_ (.A(_06599_),
    .B(_06600_),
    .Y(_06601_));
 sky130_fd_sc_hd__clkbuf_4 _14118_ (.A(_06601_),
    .X(_06602_));
 sky130_fd_sc_hd__buf_4 _14119_ (.A(_06602_),
    .X(_06603_));
 sky130_fd_sc_hd__buf_4 _14120_ (.A(\wfg_stim_sine_top.gain_val_q[2] ),
    .X(_06604_));
 sky130_fd_sc_hd__clkbuf_8 _14121_ (.A(_06604_),
    .X(_06605_));
 sky130_fd_sc_hd__a21oi_4 _14122_ (.A1(_06605_),
    .A2(_06541_),
    .B1(_06537_),
    .Y(_06606_));
 sky130_fd_sc_hd__buf_4 _14123_ (.A(_06606_),
    .X(_06607_));
 sky130_fd_sc_hd__a21oi_1 _14124_ (.A1(_06556_),
    .A2(_06560_),
    .B1(_06558_),
    .Y(_06608_));
 sky130_fd_sc_hd__or2_1 _14125_ (.A(_06607_),
    .B(_06608_),
    .X(_06609_));
 sky130_fd_sc_hd__nand2_1 _14126_ (.A(_06607_),
    .B(_06608_),
    .Y(_06610_));
 sky130_fd_sc_hd__nand2_1 _14127_ (.A(_06609_),
    .B(_06610_),
    .Y(_06611_));
 sky130_fd_sc_hd__xnor2_1 _14128_ (.A(_06603_),
    .B(_06611_),
    .Y(_06612_));
 sky130_fd_sc_hd__nor3_1 _14129_ (.A(_06597_),
    .B(_06598_),
    .C(_06612_),
    .Y(_06613_));
 sky130_fd_sc_hd__or2_1 _14130_ (.A(_06579_),
    .B(_06587_),
    .X(_06614_));
 sky130_fd_sc_hd__a31o_1 _14131_ (.A1(_06451_),
    .A2(_06600_),
    .A3(_06567_),
    .B1(_06565_),
    .X(_06615_));
 sky130_fd_sc_hd__nand2_1 _14132_ (.A(_06495_),
    .B(_06615_),
    .Y(_06616_));
 sky130_fd_sc_hd__or2_1 _14133_ (.A(_06495_),
    .B(_06615_),
    .X(_06617_));
 sky130_fd_sc_hd__nand2_1 _14134_ (.A(_06616_),
    .B(_06617_),
    .Y(_06618_));
 sky130_fd_sc_hd__or2_1 _14135_ (.A(_06493_),
    .B(_06618_),
    .X(_06619_));
 sky130_fd_sc_hd__nand2_1 _14136_ (.A(_06493_),
    .B(_06618_),
    .Y(_06620_));
 sky130_fd_sc_hd__nand2_2 _14137_ (.A(_06619_),
    .B(_06620_),
    .Y(_06621_));
 sky130_fd_sc_hd__or3_1 _14138_ (.A(_06571_),
    .B(_06572_),
    .C(_06574_),
    .X(_06622_));
 sky130_fd_sc_hd__nand2_1 _14139_ (.A(_06568_),
    .B(_06575_),
    .Y(_06623_));
 sky130_fd_sc_hd__nand2_1 _14140_ (.A(_06509_),
    .B(_06525_),
    .Y(_06624_));
 sky130_fd_sc_hd__and4_1 _14141_ (.A(_06406_),
    .B(_06505_),
    .C(_06472_),
    .D(_06473_),
    .X(_06625_));
 sky130_fd_sc_hd__a22o_1 _14142_ (.A1(_06505_),
    .A2(_06472_),
    .B1(_06473_),
    .B2(_06406_),
    .X(_06626_));
 sky130_fd_sc_hd__and2b_1 _14143_ (.A_N(_06625_),
    .B(_06626_),
    .X(_06627_));
 sky130_fd_sc_hd__xnor2_1 _14144_ (.A(_06624_),
    .B(_06627_),
    .Y(_06628_));
 sky130_fd_sc_hd__nor2_1 _14145_ (.A(_06569_),
    .B(_06571_),
    .Y(_06629_));
 sky130_fd_sc_hd__xnor2_1 _14146_ (.A(_06628_),
    .B(_06629_),
    .Y(_06630_));
 sky130_fd_sc_hd__nand2_1 _14147_ (.A(_06568_),
    .B(_06630_),
    .Y(_06631_));
 sky130_fd_sc_hd__or2_1 _14148_ (.A(_06568_),
    .B(_06630_),
    .X(_06632_));
 sky130_fd_sc_hd__nand2_1 _14149_ (.A(_06631_),
    .B(_06632_),
    .Y(_06633_));
 sky130_fd_sc_hd__a21o_1 _14150_ (.A1(_06622_),
    .A2(_06623_),
    .B1(_06633_),
    .X(_06634_));
 sky130_fd_sc_hd__nand3_1 _14151_ (.A(_06633_),
    .B(_06622_),
    .C(_06623_),
    .Y(_06635_));
 sky130_fd_sc_hd__nand2_1 _14152_ (.A(_06634_),
    .B(_06635_),
    .Y(_06636_));
 sky130_fd_sc_hd__xnor2_1 _14153_ (.A(_06621_),
    .B(_06636_),
    .Y(_06637_));
 sky130_fd_sc_hd__a21oi_1 _14154_ (.A1(_06577_),
    .A2(_06614_),
    .B1(_06637_),
    .Y(_06638_));
 sky130_fd_sc_hd__and3_1 _14155_ (.A(_06637_),
    .B(_06577_),
    .C(_06614_),
    .X(_06639_));
 sky130_fd_sc_hd__a21oi_1 _14156_ (.A1(_06582_),
    .A2(_06585_),
    .B1(_06557_),
    .Y(_06640_));
 sky130_fd_sc_hd__and3_1 _14157_ (.A(_06557_),
    .B(_06582_),
    .C(_06585_),
    .X(_06641_));
 sky130_fd_sc_hd__nor2_1 _14158_ (.A(_06640_),
    .B(_06641_),
    .Y(_06642_));
 sky130_fd_sc_hd__xnor2_1 _14159_ (.A(_06556_),
    .B(_06642_),
    .Y(_06643_));
 sky130_fd_sc_hd__or3_1 _14160_ (.A(_06638_),
    .B(_06639_),
    .C(_06643_),
    .X(_06644_));
 sky130_fd_sc_hd__o21ai_1 _14161_ (.A1(_06638_),
    .A2(_06639_),
    .B1(_06643_),
    .Y(_06645_));
 sky130_fd_sc_hd__o211a_1 _14162_ (.A1(_06589_),
    .A2(_06594_),
    .B1(_06644_),
    .C1(_06645_),
    .X(_06646_));
 sky130_fd_sc_hd__a211oi_1 _14163_ (.A1(_06644_),
    .A2(_06645_),
    .B1(_06589_),
    .C1(_06594_),
    .Y(_06647_));
 sky130_fd_sc_hd__xnor2_4 _14164_ (.A(_06541_),
    .B(_06542_),
    .Y(_06648_));
 sky130_fd_sc_hd__xnor2_4 _14165_ (.A(_06648_),
    .B(_06554_),
    .Y(_06649_));
 sky130_fd_sc_hd__and2_1 _14166_ (.A(_06649_),
    .B(_06591_),
    .X(_06650_));
 sky130_fd_sc_hd__a21oi_1 _14167_ (.A1(_06556_),
    .A2(_06592_),
    .B1(_06650_),
    .Y(_06651_));
 sky130_fd_sc_hd__or2_1 _14168_ (.A(_06607_),
    .B(_06651_),
    .X(_06652_));
 sky130_fd_sc_hd__buf_4 _14169_ (.A(_06607_),
    .X(_06653_));
 sky130_fd_sc_hd__nand2_1 _14170_ (.A(_06653_),
    .B(_06651_),
    .Y(_06654_));
 sky130_fd_sc_hd__nand2_1 _14171_ (.A(_06652_),
    .B(_06654_),
    .Y(_06655_));
 sky130_fd_sc_hd__xnor2_1 _14172_ (.A(_06603_),
    .B(_06655_),
    .Y(_06656_));
 sky130_fd_sc_hd__or3_1 _14173_ (.A(_06646_),
    .B(_06647_),
    .C(_06656_),
    .X(_06657_));
 sky130_fd_sc_hd__o21ai_1 _14174_ (.A1(_06646_),
    .A2(_06647_),
    .B1(_06656_),
    .Y(_06658_));
 sky130_fd_sc_hd__o211a_1 _14175_ (.A1(_06597_),
    .A2(_06613_),
    .B1(_06657_),
    .C1(_06658_),
    .X(_06659_));
 sky130_fd_sc_hd__o21a_1 _14176_ (.A1(_06603_),
    .A2(_06611_),
    .B1(_06609_),
    .X(_06660_));
 sky130_fd_sc_hd__a211oi_1 _14177_ (.A1(_06657_),
    .A2(_06658_),
    .B1(_06597_),
    .C1(_06613_),
    .Y(_06661_));
 sky130_fd_sc_hd__nor2_1 _14178_ (.A(_06659_),
    .B(_06661_),
    .Y(_06662_));
 sky130_fd_sc_hd__and2b_1 _14179_ (.A_N(_06660_),
    .B(_06662_),
    .X(_06663_));
 sky130_fd_sc_hd__and2b_1 _14180_ (.A_N(_06646_),
    .B(_06657_),
    .X(_06664_));
 sky130_fd_sc_hd__a21o_1 _14181_ (.A1(_06577_),
    .A2(_06614_),
    .B1(_06637_),
    .X(_06665_));
 sky130_fd_sc_hd__a21oi_1 _14182_ (.A1(_06616_),
    .A2(_06619_),
    .B1(_06557_),
    .Y(_06666_));
 sky130_fd_sc_hd__and3_1 _14183_ (.A(_06557_),
    .B(_06616_),
    .C(_06619_),
    .X(_06667_));
 sky130_fd_sc_hd__nor2_1 _14184_ (.A(_06666_),
    .B(_06667_),
    .Y(_06668_));
 sky130_fd_sc_hd__xnor2_2 _14185_ (.A(_06556_),
    .B(_06668_),
    .Y(_06669_));
 sky130_fd_sc_hd__or2b_1 _14186_ (.A(_06629_),
    .B_N(_06628_),
    .X(_06670_));
 sky130_fd_sc_hd__a31o_1 _14187_ (.A1(_06509_),
    .A2(_06600_),
    .A3(_06626_),
    .B1(_06625_),
    .X(_06671_));
 sky130_fd_sc_hd__buf_6 _14188_ (.A(_06454_),
    .X(_06672_));
 sky130_fd_sc_hd__nand2_1 _14189_ (.A(_06406_),
    .B(_06672_),
    .Y(_06673_));
 sky130_fd_sc_hd__nand2_2 _14190_ (.A(_06412_),
    .B(\wfg_stim_sine_top.gain_val_q[13] ),
    .Y(_06674_));
 sky130_fd_sc_hd__or2_1 _14191_ (.A(_06505_),
    .B(_06509_),
    .X(_06675_));
 sky130_fd_sc_hd__and3_1 _14192_ (.A(_06525_),
    .B(_06674_),
    .C(_06675_),
    .X(_06676_));
 sky130_fd_sc_hd__xnor2_1 _14193_ (.A(_06673_),
    .B(_06676_),
    .Y(_06677_));
 sky130_fd_sc_hd__and2_1 _14194_ (.A(_06671_),
    .B(_06677_),
    .X(_06678_));
 sky130_fd_sc_hd__nor2_1 _14195_ (.A(_06671_),
    .B(_06677_),
    .Y(_06679_));
 sky130_fd_sc_hd__nor2_1 _14196_ (.A(_06678_),
    .B(_06679_),
    .Y(_06680_));
 sky130_fd_sc_hd__xnor2_1 _14197_ (.A(_06568_),
    .B(_06680_),
    .Y(_06681_));
 sky130_fd_sc_hd__a21o_1 _14198_ (.A1(_06670_),
    .A2(_06631_),
    .B1(_06681_),
    .X(_06682_));
 sky130_fd_sc_hd__nand3_1 _14199_ (.A(_06681_),
    .B(_06670_),
    .C(_06631_),
    .Y(_06683_));
 sky130_fd_sc_hd__nand2_1 _14200_ (.A(_06682_),
    .B(_06683_),
    .Y(_06684_));
 sky130_fd_sc_hd__xnor2_1 _14201_ (.A(_06621_),
    .B(_06684_),
    .Y(_06685_));
 sky130_fd_sc_hd__o21a_1 _14202_ (.A1(_06621_),
    .A2(_06636_),
    .B1(_06634_),
    .X(_06686_));
 sky130_fd_sc_hd__or2_1 _14203_ (.A(_06685_),
    .B(_06686_),
    .X(_06687_));
 sky130_fd_sc_hd__nand2_1 _14204_ (.A(_06685_),
    .B(_06686_),
    .Y(_06688_));
 sky130_fd_sc_hd__nand2_1 _14205_ (.A(_06687_),
    .B(_06688_),
    .Y(_06689_));
 sky130_fd_sc_hd__xnor2_1 _14206_ (.A(_06669_),
    .B(_06689_),
    .Y(_06690_));
 sky130_fd_sc_hd__a21o_1 _14207_ (.A1(_06665_),
    .A2(_06644_),
    .B1(_06690_),
    .X(_06691_));
 sky130_fd_sc_hd__nand3_1 _14208_ (.A(_06690_),
    .B(_06665_),
    .C(_06644_),
    .Y(_06692_));
 sky130_fd_sc_hd__nand2_1 _14209_ (.A(_06691_),
    .B(_06692_),
    .Y(_06693_));
 sky130_fd_sc_hd__a21oi_1 _14210_ (.A1(_06556_),
    .A2(_06642_),
    .B1(_06640_),
    .Y(_06694_));
 sky130_fd_sc_hd__or2_1 _14211_ (.A(_06653_),
    .B(_06694_),
    .X(_06695_));
 sky130_fd_sc_hd__nand2_1 _14212_ (.A(_06653_),
    .B(_06694_),
    .Y(_06696_));
 sky130_fd_sc_hd__nand2_1 _14213_ (.A(_06695_),
    .B(_06696_),
    .Y(_06697_));
 sky130_fd_sc_hd__xor2_1 _14214_ (.A(_06603_),
    .B(_06697_),
    .X(_06698_));
 sky130_fd_sc_hd__xnor2_1 _14215_ (.A(_06693_),
    .B(_06698_),
    .Y(_06699_));
 sky130_fd_sc_hd__and2b_1 _14216_ (.A_N(_06664_),
    .B(_06699_),
    .X(_06700_));
 sky130_fd_sc_hd__and2b_1 _14217_ (.A_N(_06699_),
    .B(_06664_),
    .X(_06701_));
 sky130_fd_sc_hd__nor2_1 _14218_ (.A(_06700_),
    .B(_06701_),
    .Y(_06702_));
 sky130_fd_sc_hd__o21ai_1 _14219_ (.A1(_06603_),
    .A2(_06655_),
    .B1(_06652_),
    .Y(_06703_));
 sky130_fd_sc_hd__xor2_1 _14220_ (.A(_06702_),
    .B(_06703_),
    .X(_06704_));
 sky130_fd_sc_hd__o21a_1 _14221_ (.A1(_06659_),
    .A2(_06663_),
    .B1(_06704_),
    .X(_06705_));
 sky130_fd_sc_hd__a22o_1 _14222_ (.A1(_06549_),
    .A2(_06409_),
    .B1(_06452_),
    .B2(_06547_),
    .X(_06706_));
 sky130_fd_sc_hd__nand2_1 _14223_ (.A(_06472_),
    .B(_06552_),
    .Y(_06707_));
 sky130_fd_sc_hd__mux2_1 _14224_ (.A0(_06706_),
    .A1(_06707_),
    .S(_06545_),
    .X(_06708_));
 sky130_fd_sc_hd__or2_1 _14225_ (.A(_06552_),
    .B(_06550_),
    .X(_06709_));
 sky130_fd_sc_hd__xnor2_1 _14226_ (.A(_06708_),
    .B(_06709_),
    .Y(_06710_));
 sky130_fd_sc_hd__o21bai_2 _14227_ (.A1(_06543_),
    .A2(_06710_),
    .B1_N(_06553_),
    .Y(_06711_));
 sky130_fd_sc_hd__and4_1 _14228_ (.A(_06487_),
    .B(_06490_),
    .C(_06440_),
    .D(_06443_),
    .X(_06712_));
 sky130_fd_sc_hd__buf_2 _14229_ (.A(\wfg_stim_sine_top.gain_val_q[9] ),
    .X(_06713_));
 sky130_fd_sc_hd__buf_4 _14230_ (.A(_06713_),
    .X(_06714_));
 sky130_fd_sc_hd__a22o_1 _14231_ (.A1(_06490_),
    .A2(_06441_),
    .B1(_06443_),
    .B2(_06714_),
    .X(_06715_));
 sky130_fd_sc_hd__or2b_1 _14232_ (.A(_06712_),
    .B_N(_06715_),
    .X(_06716_));
 sky130_fd_sc_hd__nand2_1 _14233_ (.A(_06486_),
    .B(_06472_),
    .Y(_06717_));
 sky130_fd_sc_hd__xnor2_1 _14234_ (.A(_06716_),
    .B(_06717_),
    .Y(_06718_));
 sky130_fd_sc_hd__a22oi_1 _14235_ (.A1(_06439_),
    .A2(_06416_),
    .B1(_06430_),
    .B2(_06444_),
    .Y(_06719_));
 sky130_fd_sc_hd__and4_1 _14236_ (.A(_06444_),
    .B(_06439_),
    .C(_06416_),
    .D(_06428_),
    .X(_06720_));
 sky130_fd_sc_hd__nor2_1 _14237_ (.A(_06719_),
    .B(_06720_),
    .Y(_06721_));
 sky130_fd_sc_hd__a31o_1 _14238_ (.A1(_06451_),
    .A2(_06432_),
    .A3(_06721_),
    .B1(_06720_),
    .X(_06722_));
 sky130_fd_sc_hd__and2b_1 _14239_ (.A_N(_06718_),
    .B(_06722_),
    .X(_06723_));
 sky130_fd_sc_hd__and4_1 _14240_ (.A(_06487_),
    .B(_06490_),
    .C(_06442_),
    .D(_06421_),
    .X(_06724_));
 sky130_fd_sc_hd__buf_6 _14241_ (.A(_06490_),
    .X(_06725_));
 sky130_fd_sc_hd__a22oi_1 _14242_ (.A1(_06725_),
    .A2(_06443_),
    .B1(_06422_),
    .B2(_06714_),
    .Y(_06726_));
 sky130_fd_sc_hd__and4bb_1 _14243_ (.A_N(_06724_),
    .B_N(_06726_),
    .C(_06485_),
    .D(_06441_),
    .X(_06727_));
 sky130_fd_sc_hd__xnor2_1 _14244_ (.A(_06722_),
    .B(_06718_),
    .Y(_06728_));
 sky130_fd_sc_hd__o21a_1 _14245_ (.A1(_06724_),
    .A2(_06727_),
    .B1(_06728_),
    .X(_06729_));
 sky130_fd_sc_hd__or3_1 _14246_ (.A(_06649_),
    .B(_06723_),
    .C(_06729_),
    .X(_06730_));
 sky130_fd_sc_hd__o21a_1 _14247_ (.A1(_06723_),
    .A2(_06729_),
    .B1(_06649_),
    .X(_06731_));
 sky130_fd_sc_hd__a21oi_1 _14248_ (.A1(_06711_),
    .A2(_06730_),
    .B1(_06731_),
    .Y(_06732_));
 sky130_fd_sc_hd__or2_1 _14249_ (.A(_06653_),
    .B(_06732_),
    .X(_06733_));
 sky130_fd_sc_hd__xnor2_1 _14250_ (.A(_06607_),
    .B(_06732_),
    .Y(_06734_));
 sky130_fd_sc_hd__or2_1 _14251_ (.A(_06602_),
    .B(_06734_),
    .X(_06735_));
 sky130_fd_sc_hd__buf_8 _14252_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[7] ),
    .X(_06736_));
 sky130_fd_sc_hd__buf_4 _14253_ (.A(_06736_),
    .X(_06737_));
 sky130_fd_sc_hd__clkbuf_4 _14254_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[6] ),
    .X(_06738_));
 sky130_fd_sc_hd__clkbuf_4 _14255_ (.A(_06738_),
    .X(_06739_));
 sky130_fd_sc_hd__and4_1 _14256_ (.A(\wfg_stim_sine_top.gain_val_q[15] ),
    .B(\wfg_stim_sine_top.gain_val_q[14] ),
    .C(_06737_),
    .D(_06739_),
    .X(_06740_));
 sky130_fd_sc_hd__buf_4 _14257_ (.A(_06736_),
    .X(_06741_));
 sky130_fd_sc_hd__clkbuf_8 _14258_ (.A(_06738_),
    .X(_06742_));
 sky130_fd_sc_hd__a22oi_1 _14259_ (.A1(_06459_),
    .A2(_06741_),
    .B1(_06742_),
    .B2(_06458_),
    .Y(_06743_));
 sky130_fd_sc_hd__buf_8 _14260_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[8] ),
    .X(_06744_));
 sky130_fd_sc_hd__buf_4 _14261_ (.A(_06744_),
    .X(_06745_));
 sky130_fd_sc_hd__and4bb_1 _14262_ (.A_N(_06740_),
    .B_N(_06743_),
    .C(\wfg_stim_sine_top.gain_val_q[13] ),
    .D(_06745_),
    .X(_06746_));
 sky130_fd_sc_hd__buf_4 _14263_ (.A(_06744_),
    .X(_06747_));
 sky130_fd_sc_hd__buf_6 _14264_ (.A(_06747_),
    .X(_06748_));
 sky130_fd_sc_hd__o2bb2a_1 _14265_ (.A1_N(_06419_),
    .A2_N(_06748_),
    .B1(_06740_),
    .B2(_06743_),
    .X(_06749_));
 sky130_fd_sc_hd__buf_6 _14266_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[5] ),
    .X(_06750_));
 sky130_fd_sc_hd__and4_1 _14267_ (.A(\wfg_stim_sine_top.gain_val_q[15] ),
    .B(\wfg_stim_sine_top.gain_val_q[14] ),
    .C(_06739_),
    .D(_06750_),
    .X(_06751_));
 sky130_fd_sc_hd__buf_6 _14268_ (.A(_06750_),
    .X(_06752_));
 sky130_fd_sc_hd__a22oi_1 _14269_ (.A1(_06459_),
    .A2(_06739_),
    .B1(_06752_),
    .B2(_06458_),
    .Y(_06753_));
 sky130_fd_sc_hd__buf_6 _14270_ (.A(_06741_),
    .X(_06754_));
 sky130_fd_sc_hd__and4bb_1 _14271_ (.A_N(_06751_),
    .B_N(_06753_),
    .C(_06419_),
    .D(_06754_),
    .X(_06755_));
 sky130_fd_sc_hd__nor2_1 _14272_ (.A(_06751_),
    .B(_06755_),
    .Y(_06756_));
 sky130_fd_sc_hd__or3_1 _14273_ (.A(_06746_),
    .B(_06749_),
    .C(_06756_),
    .X(_06757_));
 sky130_fd_sc_hd__nor2_1 _14274_ (.A(_06746_),
    .B(_06749_),
    .Y(_06758_));
 sky130_fd_sc_hd__xnor2_1 _14275_ (.A(_06758_),
    .B(_06756_),
    .Y(_06759_));
 sky130_fd_sc_hd__nand2_1 _14276_ (.A(_06468_),
    .B(_06432_),
    .Y(_06760_));
 sky130_fd_sc_hd__xnor2_1 _14277_ (.A(_06721_),
    .B(_06760_),
    .Y(_06761_));
 sky130_fd_sc_hd__nand2_1 _14278_ (.A(_06759_),
    .B(_06761_),
    .Y(_06762_));
 sky130_fd_sc_hd__and4_1 _14279_ (.A(_06458_),
    .B(_06459_),
    .C(_06745_),
    .D(_06741_),
    .X(_06763_));
 sky130_fd_sc_hd__a22oi_1 _14280_ (.A1(_06412_),
    .A2(_06745_),
    .B1(_06754_),
    .B2(_06405_),
    .Y(_06764_));
 sky130_fd_sc_hd__and4bb_1 _14281_ (.A_N(_06763_),
    .B_N(_06764_),
    .C(_06419_),
    .D(_06430_),
    .X(_06765_));
 sky130_fd_sc_hd__o2bb2a_1 _14282_ (.A1_N(_06420_),
    .A2_N(_06430_),
    .B1(_06763_),
    .B2(_06764_),
    .X(_06766_));
 sky130_fd_sc_hd__nor2_1 _14283_ (.A(_06765_),
    .B(_06766_),
    .Y(_06767_));
 sky130_fd_sc_hd__nor2_1 _14284_ (.A(_06740_),
    .B(_06746_),
    .Y(_06768_));
 sky130_fd_sc_hd__xnor2_1 _14285_ (.A(_06767_),
    .B(_06768_),
    .Y(_06769_));
 sky130_fd_sc_hd__buf_6 _14286_ (.A(_06416_),
    .X(_06770_));
 sky130_fd_sc_hd__a22oi_1 _14287_ (.A1(_06471_),
    .A2(_06432_),
    .B1(_06770_),
    .B2(_06474_),
    .Y(_06771_));
 sky130_fd_sc_hd__and4_1 _14288_ (.A(_06474_),
    .B(_06471_),
    .C(_06432_),
    .D(_06770_),
    .X(_06772_));
 sky130_fd_sc_hd__nor2_1 _14289_ (.A(_06771_),
    .B(_06772_),
    .Y(_06773_));
 sky130_fd_sc_hd__nand2_1 _14290_ (.A(_06451_),
    .B(_06423_),
    .Y(_06774_));
 sky130_fd_sc_hd__xnor2_1 _14291_ (.A(_06773_),
    .B(_06774_),
    .Y(_06775_));
 sky130_fd_sc_hd__xnor2_1 _14292_ (.A(_06769_),
    .B(_06775_),
    .Y(_06776_));
 sky130_fd_sc_hd__a21o_1 _14293_ (.A1(_06757_),
    .A2(_06762_),
    .B1(_06776_),
    .X(_06777_));
 sky130_fd_sc_hd__nand3_1 _14294_ (.A(_06776_),
    .B(_06757_),
    .C(_06762_),
    .Y(_06778_));
 sky130_fd_sc_hd__nor3_1 _14295_ (.A(_06724_),
    .B(_06727_),
    .C(_06728_),
    .Y(_06779_));
 sky130_fd_sc_hd__nor2_1 _14296_ (.A(_06729_),
    .B(_06779_),
    .Y(_06780_));
 sky130_fd_sc_hd__nand3_1 _14297_ (.A(_06777_),
    .B(_06778_),
    .C(_06780_),
    .Y(_06781_));
 sky130_fd_sc_hd__or3_1 _14298_ (.A(_06765_),
    .B(_06766_),
    .C(_06768_),
    .X(_06782_));
 sky130_fd_sc_hd__nand2_1 _14299_ (.A(_06769_),
    .B(_06775_),
    .Y(_06783_));
 sky130_fd_sc_hd__and4_1 _14300_ (.A(_06458_),
    .B(_06459_),
    .C(_06428_),
    .D(_06745_),
    .X(_06784_));
 sky130_fd_sc_hd__a22oi_1 _14301_ (.A1(_06412_),
    .A2(_06428_),
    .B1(_06748_),
    .B2(_06405_),
    .Y(_06785_));
 sky130_fd_sc_hd__and4bb_1 _14302_ (.A_N(_06784_),
    .B_N(_06785_),
    .C(_06419_),
    .D(_06770_),
    .X(_06786_));
 sky130_fd_sc_hd__o2bb2a_1 _14303_ (.A1_N(_06420_),
    .A2_N(_06770_),
    .B1(_06784_),
    .B2(_06785_),
    .X(_06787_));
 sky130_fd_sc_hd__nor2_1 _14304_ (.A(_06786_),
    .B(_06787_),
    .Y(_06788_));
 sky130_fd_sc_hd__nor2_1 _14305_ (.A(_06763_),
    .B(_06765_),
    .Y(_06789_));
 sky130_fd_sc_hd__xnor2_1 _14306_ (.A(_06788_),
    .B(_06789_),
    .Y(_06790_));
 sky130_fd_sc_hd__a22oi_1 _14307_ (.A1(_06439_),
    .A2(_06422_),
    .B1(_06414_),
    .B2(_06444_),
    .Y(_06791_));
 sky130_fd_sc_hd__and4_1 _14308_ (.A(_06446_),
    .B(_06447_),
    .C(_06421_),
    .D(_06413_),
    .X(_06792_));
 sky130_fd_sc_hd__or2_1 _14309_ (.A(_06791_),
    .B(_06792_),
    .X(_06793_));
 sky130_fd_sc_hd__nand2_1 _14310_ (.A(_06468_),
    .B(_06463_),
    .Y(_06794_));
 sky130_fd_sc_hd__xnor2_1 _14311_ (.A(_06793_),
    .B(_06794_),
    .Y(_06795_));
 sky130_fd_sc_hd__inv_2 _14312_ (.A(_06795_),
    .Y(_06796_));
 sky130_fd_sc_hd__xnor2_1 _14313_ (.A(_06790_),
    .B(_06796_),
    .Y(_06797_));
 sky130_fd_sc_hd__a21oi_2 _14314_ (.A1(_06782_),
    .A2(_06783_),
    .B1(_06797_),
    .Y(_06798_));
 sky130_fd_sc_hd__and3_1 _14315_ (.A(_06797_),
    .B(_06782_),
    .C(_06783_),
    .X(_06799_));
 sky130_fd_sc_hd__a31o_1 _14316_ (.A1(_06486_),
    .A2(_06672_),
    .A3(_06715_),
    .B1(_06712_),
    .X(_06800_));
 sky130_fd_sc_hd__o21ba_1 _14317_ (.A1(_06771_),
    .A2(_06774_),
    .B1_N(_06772_),
    .X(_06801_));
 sky130_fd_sc_hd__and4_1 _14318_ (.A(_06714_),
    .B(_06725_),
    .C(_06452_),
    .D(_06441_),
    .X(_06802_));
 sky130_fd_sc_hd__a22o_1 _14319_ (.A1(_06725_),
    .A2(_06453_),
    .B1(_06441_),
    .B2(_06714_),
    .X(_06803_));
 sky130_fd_sc_hd__and2b_1 _14320_ (.A_N(_06802_),
    .B(_06803_),
    .X(_06804_));
 sky130_fd_sc_hd__xnor2_1 _14321_ (.A(_06494_),
    .B(_06804_),
    .Y(_06805_));
 sky130_fd_sc_hd__xnor2_1 _14322_ (.A(_06801_),
    .B(_06805_),
    .Y(_06806_));
 sky130_fd_sc_hd__xnor2_1 _14323_ (.A(_06800_),
    .B(_06806_),
    .Y(_06807_));
 sky130_fd_sc_hd__nor3_2 _14324_ (.A(_06798_),
    .B(_06799_),
    .C(_06807_),
    .Y(_06808_));
 sky130_fd_sc_hd__o21a_1 _14325_ (.A1(_06798_),
    .A2(_06799_),
    .B1(_06807_),
    .X(_06809_));
 sky130_fd_sc_hd__a211oi_2 _14326_ (.A1(_06777_),
    .A2(_06781_),
    .B1(_06808_),
    .C1(_06809_),
    .Y(_06810_));
 sky130_fd_sc_hd__o211a_1 _14327_ (.A1(_06808_),
    .A2(_06809_),
    .B1(_06777_),
    .C1(_06781_),
    .X(_06811_));
 sky130_fd_sc_hd__and2b_1 _14328_ (.A_N(_06731_),
    .B(_06730_),
    .X(_06812_));
 sky130_fd_sc_hd__xnor2_1 _14329_ (.A(_06711_),
    .B(_06812_),
    .Y(_06813_));
 sky130_fd_sc_hd__nor3_2 _14330_ (.A(_06810_),
    .B(_06811_),
    .C(_06813_),
    .Y(_06814_));
 sky130_fd_sc_hd__or3_1 _14331_ (.A(_06786_),
    .B(_06787_),
    .C(_06789_),
    .X(_06815_));
 sky130_fd_sc_hd__nand2_1 _14332_ (.A(_06790_),
    .B(_06796_),
    .Y(_06816_));
 sky130_fd_sc_hd__o2bb2a_1 _14333_ (.A1_N(_06420_),
    .A2_N(_06432_),
    .B1(_06429_),
    .B2(_06431_),
    .X(_06817_));
 sky130_fd_sc_hd__nor2_1 _14334_ (.A(_06433_),
    .B(_06817_),
    .Y(_06818_));
 sky130_fd_sc_hd__nor2_1 _14335_ (.A(_06784_),
    .B(_06786_),
    .Y(_06819_));
 sky130_fd_sc_hd__xnor2_1 _14336_ (.A(_06818_),
    .B(_06819_),
    .Y(_06820_));
 sky130_fd_sc_hd__a22o_1 _14337_ (.A1(_06439_),
    .A2(_06463_),
    .B1(_06423_),
    .B2(_06444_),
    .X(_06821_));
 sky130_fd_sc_hd__and4_1 _14338_ (.A(_06444_),
    .B(_06439_),
    .C(_06443_),
    .D(_06422_),
    .X(_06822_));
 sky130_fd_sc_hd__inv_2 _14339_ (.A(_06822_),
    .Y(_06823_));
 sky130_fd_sc_hd__a22oi_1 _14340_ (.A1(_06451_),
    .A2(_06510_),
    .B1(_06821_),
    .B2(_06823_),
    .Y(_06824_));
 sky130_fd_sc_hd__and4_1 _14341_ (.A(_06451_),
    .B(_06510_),
    .C(_06821_),
    .D(_06823_),
    .X(_06825_));
 sky130_fd_sc_hd__nor2_1 _14342_ (.A(_06824_),
    .B(_06825_),
    .Y(_06826_));
 sky130_fd_sc_hd__xnor2_1 _14343_ (.A(_06820_),
    .B(_06826_),
    .Y(_06827_));
 sky130_fd_sc_hd__a21o_1 _14344_ (.A1(_06815_),
    .A2(_06816_),
    .B1(_06827_),
    .X(_06828_));
 sky130_fd_sc_hd__nand3_1 _14345_ (.A(_06827_),
    .B(_06815_),
    .C(_06816_),
    .Y(_06829_));
 sky130_fd_sc_hd__a31o_1 _14346_ (.A1(_06486_),
    .A2(_06525_),
    .A3(_06803_),
    .B1(_06802_),
    .X(_06830_));
 sky130_fd_sc_hd__o21ba_1 _14347_ (.A1(_06791_),
    .A2(_06794_),
    .B1_N(_06792_),
    .X(_06831_));
 sky130_fd_sc_hd__nand2_1 _14348_ (.A(_06472_),
    .B(_06489_),
    .Y(_06832_));
 sky130_fd_sc_hd__a22o_1 _14349_ (.A1(_06725_),
    .A2(_06469_),
    .B1(_06453_),
    .B2(_06714_),
    .X(_06833_));
 sky130_fd_sc_hd__and3b_1 _14350_ (.A_N(_06494_),
    .B(_06832_),
    .C(_06833_),
    .X(_06834_));
 sky130_fd_sc_hd__a21boi_1 _14351_ (.A1(_06832_),
    .A2(_06833_),
    .B1_N(_06494_),
    .Y(_06835_));
 sky130_fd_sc_hd__nor2_1 _14352_ (.A(_06834_),
    .B(_06835_),
    .Y(_06836_));
 sky130_fd_sc_hd__xnor2_1 _14353_ (.A(_06831_),
    .B(_06836_),
    .Y(_06837_));
 sky130_fd_sc_hd__xor2_1 _14354_ (.A(_06830_),
    .B(_06837_),
    .X(_06838_));
 sky130_fd_sc_hd__nand3_2 _14355_ (.A(_06828_),
    .B(_06829_),
    .C(_06838_),
    .Y(_06839_));
 sky130_fd_sc_hd__a21o_1 _14356_ (.A1(_06828_),
    .A2(_06829_),
    .B1(_06838_),
    .X(_06840_));
 sky130_fd_sc_hd__o211a_1 _14357_ (.A1(_06798_),
    .A2(_06808_),
    .B1(_06839_),
    .C1(_06840_),
    .X(_06841_));
 sky130_fd_sc_hd__a211oi_2 _14358_ (.A1(_06839_),
    .A2(_06840_),
    .B1(_06798_),
    .C1(_06808_),
    .Y(_06842_));
 sky130_fd_sc_hd__or2b_1 _14359_ (.A(_06801_),
    .B_N(_06805_),
    .X(_06843_));
 sky130_fd_sc_hd__a21bo_1 _14360_ (.A1(_06800_),
    .A2(_06806_),
    .B1_N(_06843_),
    .X(_06844_));
 sky130_fd_sc_hd__xnor2_1 _14361_ (.A(_06557_),
    .B(_06844_),
    .Y(_06845_));
 sky130_fd_sc_hd__xnor2_1 _14362_ (.A(_06555_),
    .B(_06845_),
    .Y(_06846_));
 sky130_fd_sc_hd__or3_1 _14363_ (.A(_06841_),
    .B(_06842_),
    .C(_06846_),
    .X(_06847_));
 sky130_fd_sc_hd__o21ai_1 _14364_ (.A1(_06841_),
    .A2(_06842_),
    .B1(_06846_),
    .Y(_06848_));
 sky130_fd_sc_hd__o211a_1 _14365_ (.A1(_06810_),
    .A2(_06814_),
    .B1(_06847_),
    .C1(_06848_),
    .X(_06849_));
 sky130_fd_sc_hd__a211oi_1 _14366_ (.A1(_06847_),
    .A2(_06848_),
    .B1(_06810_),
    .C1(_06814_),
    .Y(_06850_));
 sky130_fd_sc_hd__or2_1 _14367_ (.A(_06849_),
    .B(_06850_),
    .X(_06851_));
 sky130_fd_sc_hd__nand2_1 _14368_ (.A(_06602_),
    .B(_06734_),
    .Y(_06852_));
 sky130_fd_sc_hd__nand2_1 _14369_ (.A(_06735_),
    .B(_06852_),
    .Y(_06853_));
 sky130_fd_sc_hd__nor2_1 _14370_ (.A(_06851_),
    .B(_06853_),
    .Y(_06854_));
 sky130_fd_sc_hd__nor3_1 _14371_ (.A(_06841_),
    .B(_06842_),
    .C(_06846_),
    .Y(_06855_));
 sky130_fd_sc_hd__or3_1 _14372_ (.A(_06433_),
    .B(_06817_),
    .C(_06819_),
    .X(_06856_));
 sky130_fd_sc_hd__nand2_1 _14373_ (.A(_06820_),
    .B(_06826_),
    .Y(_06857_));
 sky130_fd_sc_hd__or2_1 _14374_ (.A(_06437_),
    .B(_06456_),
    .X(_06858_));
 sky130_fd_sc_hd__nand2_1 _14375_ (.A(_06457_),
    .B(_06858_),
    .Y(_06859_));
 sky130_fd_sc_hd__a21o_2 _14376_ (.A1(_06856_),
    .A2(_06857_),
    .B1(_06859_),
    .X(_06860_));
 sky130_fd_sc_hd__nand3_1 _14377_ (.A(_06859_),
    .B(_06856_),
    .C(_06857_),
    .Y(_06861_));
 sky130_fd_sc_hd__a21o_1 _14378_ (.A1(_06672_),
    .A2(_06489_),
    .B1(_06834_),
    .X(_06862_));
 sky130_fd_sc_hd__nor2_1 _14379_ (.A(_06822_),
    .B(_06825_),
    .Y(_06863_));
 sky130_fd_sc_hd__xnor2_1 _14380_ (.A(_06495_),
    .B(_06863_),
    .Y(_06864_));
 sky130_fd_sc_hd__xor2_2 _14381_ (.A(_06862_),
    .B(_06864_),
    .X(_06865_));
 sky130_fd_sc_hd__and3_1 _14382_ (.A(_06860_),
    .B(_06861_),
    .C(_06865_),
    .X(_06866_));
 sky130_fd_sc_hd__a21oi_2 _14383_ (.A1(_06860_),
    .A2(_06861_),
    .B1(_06865_),
    .Y(_06867_));
 sky130_fd_sc_hd__a211oi_4 _14384_ (.A1(_06828_),
    .A2(_06839_),
    .B1(_06866_),
    .C1(_06867_),
    .Y(_06868_));
 sky130_fd_sc_hd__o211a_1 _14385_ (.A1(_06866_),
    .A2(_06867_),
    .B1(_06828_),
    .C1(_06839_),
    .X(_06869_));
 sky130_fd_sc_hd__or2b_1 _14386_ (.A(_06831_),
    .B_N(_06836_),
    .X(_06870_));
 sky130_fd_sc_hd__a21bo_1 _14387_ (.A1(_06830_),
    .A2(_06837_),
    .B1_N(_06870_),
    .X(_06871_));
 sky130_fd_sc_hd__xnor2_1 _14388_ (.A(_06557_),
    .B(_06871_),
    .Y(_06872_));
 sky130_fd_sc_hd__xnor2_1 _14389_ (.A(_06556_),
    .B(_06872_),
    .Y(_06873_));
 sky130_fd_sc_hd__or3_1 _14390_ (.A(_06868_),
    .B(_06869_),
    .C(_06873_),
    .X(_06874_));
 sky130_fd_sc_hd__o21ai_1 _14391_ (.A1(_06868_),
    .A2(_06869_),
    .B1(_06873_),
    .Y(_06875_));
 sky130_fd_sc_hd__o211a_2 _14392_ (.A1(_06841_),
    .A2(_06855_),
    .B1(_06874_),
    .C1(_06875_),
    .X(_06876_));
 sky130_fd_sc_hd__a211oi_2 _14393_ (.A1(_06874_),
    .A2(_06875_),
    .B1(_06841_),
    .C1(_06855_),
    .Y(_06877_));
 sky130_fd_sc_hd__and2_1 _14394_ (.A(_06649_),
    .B(_06844_),
    .X(_06878_));
 sky130_fd_sc_hd__a21oi_1 _14395_ (.A1(_06555_),
    .A2(_06845_),
    .B1(_06878_),
    .Y(_06879_));
 sky130_fd_sc_hd__nor2_1 _14396_ (.A(_06606_),
    .B(_06879_),
    .Y(_06880_));
 sky130_fd_sc_hd__and2_1 _14397_ (.A(_06606_),
    .B(_06879_),
    .X(_06881_));
 sky130_fd_sc_hd__or2_1 _14398_ (.A(_06880_),
    .B(_06881_),
    .X(_06882_));
 sky130_fd_sc_hd__nor2_1 _14399_ (.A(_06602_),
    .B(_06882_),
    .Y(_06883_));
 sky130_fd_sc_hd__and2_1 _14400_ (.A(_06602_),
    .B(_06882_),
    .X(_06884_));
 sky130_fd_sc_hd__or2_1 _14401_ (.A(_06883_),
    .B(_06884_),
    .X(_06885_));
 sky130_fd_sc_hd__or3_1 _14402_ (.A(_06876_),
    .B(_06877_),
    .C(_06885_),
    .X(_06886_));
 sky130_fd_sc_hd__o21ai_1 _14403_ (.A1(_06876_),
    .A2(_06877_),
    .B1(_06885_),
    .Y(_06887_));
 sky130_fd_sc_hd__o211a_1 _14404_ (.A1(_06849_),
    .A2(_06854_),
    .B1(_06886_),
    .C1(_06887_),
    .X(_06888_));
 sky130_fd_sc_hd__a211oi_1 _14405_ (.A1(_06886_),
    .A2(_06887_),
    .B1(_06849_),
    .C1(_06854_),
    .Y(_06889_));
 sky130_fd_sc_hd__a211oi_2 _14406_ (.A1(_06733_),
    .A2(_06735_),
    .B1(_06888_),
    .C1(_06889_),
    .Y(_06890_));
 sky130_fd_sc_hd__o211a_1 _14407_ (.A1(_06888_),
    .A2(_06889_),
    .B1(_06733_),
    .C1(_06735_),
    .X(_06891_));
 sky130_fd_sc_hd__xnor2_1 _14408_ (.A(_06851_),
    .B(_06853_),
    .Y(_06892_));
 sky130_fd_sc_hd__o2bb2a_1 _14409_ (.A1_N(_06419_),
    .A2_N(_06754_),
    .B1(_06751_),
    .B2(_06753_),
    .X(_06893_));
 sky130_fd_sc_hd__buf_4 _14410_ (.A(_06750_),
    .X(_06894_));
 sky130_fd_sc_hd__buf_6 _14411_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[4] ),
    .X(_06895_));
 sky130_fd_sc_hd__buf_4 _14412_ (.A(_06895_),
    .X(_06896_));
 sky130_fd_sc_hd__nand4_1 _14413_ (.A(_06458_),
    .B(_06459_),
    .C(_06894_),
    .D(_06896_),
    .Y(_06897_));
 sky130_fd_sc_hd__a22o_1 _14414_ (.A1(_06459_),
    .A2(_06894_),
    .B1(_06896_),
    .B2(_06458_),
    .X(_06898_));
 sky130_fd_sc_hd__nand4_1 _14415_ (.A(_06419_),
    .B(_06742_),
    .C(_06897_),
    .D(_06898_),
    .Y(_06899_));
 sky130_fd_sc_hd__and2_1 _14416_ (.A(_06897_),
    .B(_06899_),
    .X(_06900_));
 sky130_fd_sc_hd__or3_1 _14417_ (.A(_06755_),
    .B(_06893_),
    .C(_06900_),
    .X(_06901_));
 sky130_fd_sc_hd__nor2_1 _14418_ (.A(_06755_),
    .B(_06893_),
    .Y(_06902_));
 sky130_fd_sc_hd__xnor2_1 _14419_ (.A(_06902_),
    .B(_06900_),
    .Y(_06903_));
 sky130_fd_sc_hd__a22o_1 _14420_ (.A1(_06439_),
    .A2(_06430_),
    .B1(_06748_),
    .B2(_06444_),
    .X(_06904_));
 sky130_fd_sc_hd__and4_1 _14421_ (.A(_06446_),
    .B(_06447_),
    .C(_06427_),
    .D(_06747_),
    .X(_06905_));
 sky130_fd_sc_hd__inv_2 _14422_ (.A(_06905_),
    .Y(_06906_));
 sky130_fd_sc_hd__nand2_1 _14423_ (.A(_06904_),
    .B(_06906_),
    .Y(_06907_));
 sky130_fd_sc_hd__nand2_1 _14424_ (.A(_06468_),
    .B(_06770_),
    .Y(_06908_));
 sky130_fd_sc_hd__xor2_1 _14425_ (.A(_06907_),
    .B(_06908_),
    .X(_06909_));
 sky130_fd_sc_hd__nand2_1 _14426_ (.A(_06903_),
    .B(_06909_),
    .Y(_06910_));
 sky130_fd_sc_hd__xnor2_1 _14427_ (.A(_06759_),
    .B(_06761_),
    .Y(_06911_));
 sky130_fd_sc_hd__a21o_1 _14428_ (.A1(_06901_),
    .A2(_06910_),
    .B1(_06911_),
    .X(_06912_));
 sky130_fd_sc_hd__nand3_1 _14429_ (.A(_06911_),
    .B(_06901_),
    .C(_06910_),
    .Y(_06913_));
 sky130_fd_sc_hd__and4_1 _14430_ (.A(_06714_),
    .B(_06490_),
    .C(_06422_),
    .D(_06414_),
    .X(_06914_));
 sky130_fd_sc_hd__a22oi_1 _14431_ (.A1(_06725_),
    .A2(_06422_),
    .B1(_06414_),
    .B2(_06714_),
    .Y(_06915_));
 sky130_fd_sc_hd__nand2_1 _14432_ (.A(_06485_),
    .B(_06463_),
    .Y(_06916_));
 sky130_fd_sc_hd__or3_1 _14433_ (.A(_06914_),
    .B(_06915_),
    .C(_06916_),
    .X(_06917_));
 sky130_fd_sc_hd__or2b_1 _14434_ (.A(_06914_),
    .B_N(_06917_),
    .X(_06918_));
 sky130_fd_sc_hd__a31oi_2 _14435_ (.A1(_06468_),
    .A2(_06770_),
    .A3(_06904_),
    .B1(_06905_),
    .Y(_06919_));
 sky130_fd_sc_hd__o2bb2a_1 _14436_ (.A1_N(_06486_),
    .A2_N(_06473_),
    .B1(_06724_),
    .B2(_06726_),
    .X(_06920_));
 sky130_fd_sc_hd__nor2_1 _14437_ (.A(_06727_),
    .B(_06920_),
    .Y(_06921_));
 sky130_fd_sc_hd__xnor2_1 _14438_ (.A(_06919_),
    .B(_06921_),
    .Y(_06922_));
 sky130_fd_sc_hd__xor2_1 _14439_ (.A(_06918_),
    .B(_06922_),
    .X(_06923_));
 sky130_fd_sc_hd__nand3_1 _14440_ (.A(_06912_),
    .B(_06913_),
    .C(_06923_),
    .Y(_06924_));
 sky130_fd_sc_hd__and3_1 _14441_ (.A(_06777_),
    .B(_06778_),
    .C(_06780_),
    .X(_06925_));
 sky130_fd_sc_hd__a21oi_1 _14442_ (.A1(_06777_),
    .A2(_06778_),
    .B1(_06780_),
    .Y(_06926_));
 sky130_fd_sc_hd__a211o_1 _14443_ (.A1(_06912_),
    .A2(_06924_),
    .B1(_06925_),
    .C1(_06926_),
    .X(_06927_));
 sky130_fd_sc_hd__o211ai_2 _14444_ (.A1(_06925_),
    .A2(_06926_),
    .B1(_06912_),
    .C1(_06924_),
    .Y(_06928_));
 sky130_fd_sc_hd__clkbuf_4 _14445_ (.A(\wfg_stim_sine_top.gain_val_q[6] ),
    .X(_06929_));
 sky130_fd_sc_hd__clkbuf_4 _14446_ (.A(\wfg_stim_sine_top.gain_val_q[5] ),
    .X(_06930_));
 sky130_fd_sc_hd__and4_1 _14447_ (.A(_06929_),
    .B(_06930_),
    .C(_06452_),
    .D(\wfg_stim_sine_top.wfg_stim_sine.sin_17[14] ),
    .X(_06931_));
 sky130_fd_sc_hd__a22oi_1 _14448_ (.A1(_06930_),
    .A2(_06452_),
    .B1(_06440_),
    .B2(_06547_),
    .Y(_06932_));
 sky130_fd_sc_hd__nor2_1 _14449_ (.A(_06931_),
    .B(_06932_),
    .Y(_06933_));
 sky130_fd_sc_hd__a31o_1 _14450_ (.A1(_06551_),
    .A2(_06469_),
    .A3(_06933_),
    .B1(_06931_),
    .X(_06934_));
 sky130_fd_sc_hd__a21bo_1 _14451_ (.A1(_06453_),
    .A2(_06552_),
    .B1_N(_06706_),
    .X(_06935_));
 sky130_fd_sc_hd__xor2_1 _14452_ (.A(_06545_),
    .B(_06935_),
    .X(_06936_));
 sky130_fd_sc_hd__xnor2_1 _14453_ (.A(_06934_),
    .B(_06936_),
    .Y(_06937_));
 sky130_fd_sc_hd__nand2_1 _14454_ (.A(_06934_),
    .B(_06936_),
    .Y(_06938_));
 sky130_fd_sc_hd__o21a_1 _14455_ (.A1(_06543_),
    .A2(_06937_),
    .B1(_06938_),
    .X(_06939_));
 sky130_fd_sc_hd__and2b_1 _14456_ (.A_N(_06919_),
    .B(_06921_),
    .X(_06940_));
 sky130_fd_sc_hd__a21oi_1 _14457_ (.A1(_06918_),
    .A2(_06922_),
    .B1(_06940_),
    .Y(_06941_));
 sky130_fd_sc_hd__xnor2_1 _14458_ (.A(_06648_),
    .B(_06710_),
    .Y(_06942_));
 sky130_fd_sc_hd__xnor2_1 _14459_ (.A(_06941_),
    .B(_06942_),
    .Y(_06943_));
 sky130_fd_sc_hd__xnor2_1 _14460_ (.A(_06939_),
    .B(_06943_),
    .Y(_06944_));
 sky130_fd_sc_hd__nand3_1 _14461_ (.A(_06927_),
    .B(_06928_),
    .C(_06944_),
    .Y(_06945_));
 sky130_fd_sc_hd__o21a_1 _14462_ (.A1(_06810_),
    .A2(_06811_),
    .B1(_06813_),
    .X(_06946_));
 sky130_fd_sc_hd__a211oi_2 _14463_ (.A1(_06927_),
    .A2(_06945_),
    .B1(_06814_),
    .C1(_06946_),
    .Y(_06947_));
 sky130_fd_sc_hd__o211a_1 _14464_ (.A1(_06814_),
    .A2(_06946_),
    .B1(_06927_),
    .C1(_06945_),
    .X(_06948_));
 sky130_fd_sc_hd__or2b_1 _14465_ (.A(_06941_),
    .B_N(_06942_),
    .X(_06949_));
 sky130_fd_sc_hd__or2b_1 _14466_ (.A(_06939_),
    .B_N(_06943_),
    .X(_06950_));
 sky130_fd_sc_hd__and2_1 _14467_ (.A(_06949_),
    .B(_06950_),
    .X(_06951_));
 sky130_fd_sc_hd__xnor2_1 _14468_ (.A(_06607_),
    .B(_06951_),
    .Y(_06952_));
 sky130_fd_sc_hd__xor2_1 _14469_ (.A(_06601_),
    .B(_06952_),
    .X(_06953_));
 sky130_fd_sc_hd__nor3b_2 _14470_ (.A(_06947_),
    .B(_06948_),
    .C_N(_06953_),
    .Y(_06954_));
 sky130_fd_sc_hd__nor2_1 _14471_ (.A(_06947_),
    .B(_06954_),
    .Y(_06955_));
 sky130_fd_sc_hd__or2_1 _14472_ (.A(_06892_),
    .B(_06955_),
    .X(_06956_));
 sky130_fd_sc_hd__nand2_1 _14473_ (.A(_06892_),
    .B(_06955_),
    .Y(_06957_));
 sky130_fd_sc_hd__nand2_1 _14474_ (.A(_06956_),
    .B(_06957_),
    .Y(_06958_));
 sky130_fd_sc_hd__or2_1 _14475_ (.A(_06653_),
    .B(_06951_),
    .X(_06959_));
 sky130_fd_sc_hd__o21a_1 _14476_ (.A1(_06603_),
    .A2(_06952_),
    .B1(_06959_),
    .X(_06960_));
 sky130_fd_sc_hd__or2_1 _14477_ (.A(_06958_),
    .B(_06960_),
    .X(_06961_));
 sky130_fd_sc_hd__o211a_1 _14478_ (.A1(_06890_),
    .A2(_06891_),
    .B1(_06956_),
    .C1(_06961_),
    .X(_06962_));
 sky130_fd_sc_hd__a211o_1 _14479_ (.A1(_06956_),
    .A2(_06961_),
    .B1(_06890_),
    .C1(_06891_),
    .X(_06963_));
 sky130_fd_sc_hd__or2b_1 _14480_ (.A(_06962_),
    .B_N(_06963_),
    .X(_06964_));
 sky130_fd_sc_hd__buf_4 _14481_ (.A(_06895_),
    .X(_06965_));
 sky130_fd_sc_hd__and4_1 _14482_ (.A(_06713_),
    .B(_06488_),
    .C(_06750_),
    .D(_06965_),
    .X(_06966_));
 sky130_fd_sc_hd__nand2_1 _14483_ (.A(_06484_),
    .B(_06742_),
    .Y(_06967_));
 sky130_fd_sc_hd__a22oi_1 _14484_ (.A1(_06488_),
    .A2(_06894_),
    .B1(_06896_),
    .B2(_06487_),
    .Y(_06968_));
 sky130_fd_sc_hd__or3_1 _14485_ (.A(_06966_),
    .B(_06967_),
    .C(_06968_),
    .X(_06969_));
 sky130_fd_sc_hd__buf_8 _14486_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[2] ),
    .X(_06970_));
 sky130_fd_sc_hd__clkbuf_4 _14487_ (.A(_06970_),
    .X(_06971_));
 sky130_fd_sc_hd__clkbuf_8 _14488_ (.A(_06971_),
    .X(_06972_));
 sky130_fd_sc_hd__buf_4 _14489_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[1] ),
    .X(_06973_));
 sky130_fd_sc_hd__buf_4 _14490_ (.A(_06973_),
    .X(_06974_));
 sky130_fd_sc_hd__buf_4 _14491_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[0] ),
    .X(_06975_));
 sky130_fd_sc_hd__a22o_1 _14492_ (.A1(_06447_),
    .A2(_06974_),
    .B1(_06975_),
    .B2(_06446_),
    .X(_06976_));
 sky130_fd_sc_hd__and4_1 _14493_ (.A(_06446_),
    .B(_06438_),
    .C(_06974_),
    .D(_06975_),
    .X(_06977_));
 sky130_fd_sc_hd__a31o_1 _14494_ (.A1(_06450_),
    .A2(_06972_),
    .A3(_06976_),
    .B1(_06977_),
    .X(_06978_));
 sky130_fd_sc_hd__o21ai_1 _14495_ (.A1(_06966_),
    .A2(_06968_),
    .B1(_06967_),
    .Y(_06979_));
 sky130_fd_sc_hd__nand3_1 _14496_ (.A(_06969_),
    .B(_06978_),
    .C(_06979_),
    .Y(_06980_));
 sky130_fd_sc_hd__a21o_1 _14497_ (.A1(_06969_),
    .A2(_06979_),
    .B1(_06978_),
    .X(_06981_));
 sky130_fd_sc_hd__clkbuf_4 _14498_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[3] ),
    .X(_06982_));
 sky130_fd_sc_hd__nand4_2 _14499_ (.A(_06487_),
    .B(_06488_),
    .C(_06896_),
    .D(_06982_),
    .Y(_06983_));
 sky130_fd_sc_hd__a22o_1 _14500_ (.A1(_06488_),
    .A2(_06965_),
    .B1(_06982_),
    .B2(_06713_),
    .X(_06984_));
 sky130_fd_sc_hd__nand4_2 _14501_ (.A(_06485_),
    .B(_06752_),
    .C(_06983_),
    .D(_06984_),
    .Y(_06985_));
 sky130_fd_sc_hd__nand2_1 _14502_ (.A(_06983_),
    .B(_06985_),
    .Y(_06986_));
 sky130_fd_sc_hd__nand3_1 _14503_ (.A(_06980_),
    .B(_06981_),
    .C(_06986_),
    .Y(_06987_));
 sky130_fd_sc_hd__a21o_1 _14504_ (.A1(_06980_),
    .A2(_06981_),
    .B1(_06986_),
    .X(_06988_));
 sky130_fd_sc_hd__clkbuf_4 _14505_ (.A(_06975_),
    .X(_06989_));
 sky130_fd_sc_hd__nand2_1 _14506_ (.A(_06420_),
    .B(_06989_),
    .Y(_06990_));
 sky130_fd_sc_hd__buf_4 _14507_ (.A(_06970_),
    .X(_06991_));
 sky130_fd_sc_hd__and3_1 _14508_ (.A(\wfg_stim_sine_top.gain_val_q[12] ),
    .B(\wfg_stim_sine_top.gain_val_q[11] ),
    .C(_06991_),
    .X(_06992_));
 sky130_fd_sc_hd__a22o_1 _14509_ (.A1(_06438_),
    .A2(_06991_),
    .B1(_06973_),
    .B2(\wfg_stim_sine_top.gain_val_q[12] ),
    .X(_06993_));
 sky130_fd_sc_hd__a21bo_1 _14510_ (.A1(_06974_),
    .A2(_06992_),
    .B1_N(_06993_),
    .X(_06994_));
 sky130_fd_sc_hd__clkbuf_8 _14511_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[3] ),
    .X(_06995_));
 sky130_fd_sc_hd__buf_6 _14512_ (.A(_06995_),
    .X(_06996_));
 sky130_fd_sc_hd__nand2_1 _14513_ (.A(\wfg_stim_sine_top.gain_val_q[10] ),
    .B(_06996_),
    .Y(_06997_));
 sky130_fd_sc_hd__xor2_1 _14514_ (.A(_06994_),
    .B(_06997_),
    .X(_06998_));
 sky130_fd_sc_hd__xnor2_1 _14515_ (.A(_06990_),
    .B(_06998_),
    .Y(_06999_));
 sky130_fd_sc_hd__nand3_2 _14516_ (.A(_06987_),
    .B(_06988_),
    .C(_06999_),
    .Y(_07000_));
 sky130_fd_sc_hd__nand2_4 _14517_ (.A(_06973_),
    .B(_06975_),
    .Y(_07001_));
 sky130_fd_sc_hd__a22o_1 _14518_ (.A1(\wfg_stim_sine_top.gain_val_q[13] ),
    .A2(_06974_),
    .B1(_06975_),
    .B2(_06412_),
    .X(_07002_));
 sky130_fd_sc_hd__o21ai_2 _14519_ (.A1(_06674_),
    .A2(_07001_),
    .B1(_07002_),
    .Y(_07003_));
 sky130_fd_sc_hd__a22oi_1 _14520_ (.A1(_06438_),
    .A2(_06995_),
    .B1(_06971_),
    .B2(\wfg_stim_sine_top.gain_val_q[12] ),
    .Y(_07004_));
 sky130_fd_sc_hd__and4_1 _14521_ (.A(\wfg_stim_sine_top.gain_val_q[12] ),
    .B(_06438_),
    .C(_06995_),
    .D(_06991_),
    .X(_07005_));
 sky130_fd_sc_hd__nor2_1 _14522_ (.A(_07004_),
    .B(_07005_),
    .Y(_07006_));
 sky130_fd_sc_hd__buf_6 _14523_ (.A(_06965_),
    .X(_07007_));
 sky130_fd_sc_hd__nand2_1 _14524_ (.A(\wfg_stim_sine_top.gain_val_q[10] ),
    .B(_07007_),
    .Y(_07008_));
 sky130_fd_sc_hd__xnor2_1 _14525_ (.A(_07006_),
    .B(_07008_),
    .Y(_07009_));
 sky130_fd_sc_hd__xnor2_2 _14526_ (.A(_07003_),
    .B(_07009_),
    .Y(_07010_));
 sky130_fd_sc_hd__or2b_1 _14527_ (.A(_06990_),
    .B_N(_06998_),
    .X(_07011_));
 sky130_fd_sc_hd__xor2_1 _14528_ (.A(_07010_),
    .B(_07011_),
    .X(_07012_));
 sky130_fd_sc_hd__or2b_1 _14529_ (.A(_06966_),
    .B_N(_06969_),
    .X(_07013_));
 sky130_fd_sc_hd__and4_1 _14530_ (.A(\wfg_stim_sine_top.gain_val_q[9] ),
    .B(\wfg_stim_sine_top.gain_val_q[8] ),
    .C(\wfg_stim_sine_top.wfg_stim_sine.sin_17[6] ),
    .D(\wfg_stim_sine_top.wfg_stim_sine.sin_17[5] ),
    .X(_07014_));
 sky130_fd_sc_hd__a22oi_1 _14531_ (.A1(\wfg_stim_sine_top.gain_val_q[8] ),
    .A2(_06738_),
    .B1(_06750_),
    .B2(\wfg_stim_sine_top.gain_val_q[9] ),
    .Y(_07015_));
 sky130_fd_sc_hd__nand2_1 _14532_ (.A(\wfg_stim_sine_top.gain_val_q[7] ),
    .B(_06737_),
    .Y(_07016_));
 sky130_fd_sc_hd__or3_1 _14533_ (.A(_07014_),
    .B(_07015_),
    .C(_07016_),
    .X(_07017_));
 sky130_fd_sc_hd__a32o_1 _14534_ (.A1(\wfg_stim_sine_top.gain_val_q[10] ),
    .A2(_06982_),
    .A3(_06993_),
    .B1(_06992_),
    .B2(_06974_),
    .X(_07018_));
 sky130_fd_sc_hd__o21ai_1 _14535_ (.A1(_07014_),
    .A2(_07015_),
    .B1(_07016_),
    .Y(_07019_));
 sky130_fd_sc_hd__and3_1 _14536_ (.A(_07017_),
    .B(_07018_),
    .C(_07019_),
    .X(_07020_));
 sky130_fd_sc_hd__a21o_1 _14537_ (.A1(_07017_),
    .A2(_07019_),
    .B1(_07018_),
    .X(_07021_));
 sky130_fd_sc_hd__and2b_1 _14538_ (.A_N(_07020_),
    .B(_07021_),
    .X(_07022_));
 sky130_fd_sc_hd__xnor2_1 _14539_ (.A(_07013_),
    .B(_07022_),
    .Y(_07023_));
 sky130_fd_sc_hd__nand2_1 _14540_ (.A(_07012_),
    .B(_07023_),
    .Y(_07024_));
 sky130_fd_sc_hd__or2_2 _14541_ (.A(_07012_),
    .B(_07023_),
    .X(_07025_));
 sky130_fd_sc_hd__and3b_1 _14542_ (.A_N(_07000_),
    .B(_07024_),
    .C(_07025_),
    .X(_07026_));
 sky130_fd_sc_hd__inv_2 _14543_ (.A(_07026_),
    .Y(_07027_));
 sky130_fd_sc_hd__a21boi_1 _14544_ (.A1(_07025_),
    .A2(_07024_),
    .B1_N(_07000_),
    .Y(_07028_));
 sky130_fd_sc_hd__and4_1 _14545_ (.A(_06546_),
    .B(_06548_),
    .C(_06744_),
    .D(_06736_),
    .X(_07029_));
 sky130_fd_sc_hd__nand2_1 _14546_ (.A(\wfg_stim_sine_top.gain_val_q[4] ),
    .B(_06427_),
    .Y(_07030_));
 sky130_fd_sc_hd__a22oi_2 _14547_ (.A1(_06548_),
    .A2(_06747_),
    .B1(_06737_),
    .B2(_06929_),
    .Y(_07031_));
 sky130_fd_sc_hd__or3_1 _14548_ (.A(_07029_),
    .B(_07030_),
    .C(_07031_),
    .X(_07032_));
 sky130_fd_sc_hd__o21ai_1 _14549_ (.A1(_07029_),
    .A2(_07031_),
    .B1(_07030_),
    .Y(_07033_));
 sky130_fd_sc_hd__and2_1 _14550_ (.A(_06544_),
    .B(_06747_),
    .X(_07034_));
 sky130_fd_sc_hd__a22o_1 _14551_ (.A1(_06930_),
    .A2(_06741_),
    .B1(_06739_),
    .B2(_06929_),
    .X(_07035_));
 sky130_fd_sc_hd__nand4_1 _14552_ (.A(_06547_),
    .B(_06930_),
    .C(_06741_),
    .D(_06739_),
    .Y(_07036_));
 sky130_fd_sc_hd__a21bo_1 _14553_ (.A1(_07034_),
    .A2(_07035_),
    .B1_N(_07036_),
    .X(_07037_));
 sky130_fd_sc_hd__nand3_2 _14554_ (.A(_07032_),
    .B(_07033_),
    .C(_07037_),
    .Y(_07038_));
 sky130_fd_sc_hd__a21o_1 _14555_ (.A1(_07032_),
    .A2(_07033_),
    .B1(_07037_),
    .X(_07039_));
 sky130_fd_sc_hd__nand2_1 _14556_ (.A(\wfg_stim_sine_top.gain_val_q[2] ),
    .B(_06414_),
    .Y(_07040_));
 sky130_fd_sc_hd__nand2_4 _14557_ (.A(\wfg_stim_sine_top.gain_val_q[1] ),
    .B(\wfg_stim_sine_top.gain_val_q[0] ),
    .Y(_07041_));
 sky130_fd_sc_hd__nand2_2 _14558_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[13] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.sin_17[12] ),
    .Y(_07042_));
 sky130_fd_sc_hd__buf_4 _14559_ (.A(\wfg_stim_sine_top.gain_val_q[0] ),
    .X(_07043_));
 sky130_fd_sc_hd__buf_4 _14560_ (.A(\wfg_stim_sine_top.gain_val_q[1] ),
    .X(_07044_));
 sky130_fd_sc_hd__a22o_1 _14561_ (.A1(_07043_),
    .A2(_06442_),
    .B1(_06421_),
    .B2(_07044_),
    .X(_07045_));
 sky130_fd_sc_hd__o21ai_1 _14562_ (.A1(_07041_),
    .A2(_07042_),
    .B1(_07045_),
    .Y(_07046_));
 sky130_fd_sc_hd__xor2_1 _14563_ (.A(_07040_),
    .B(_07046_),
    .X(_07047_));
 sky130_fd_sc_hd__nand3_2 _14564_ (.A(_07038_),
    .B(_07039_),
    .C(_07047_),
    .Y(_07048_));
 sky130_fd_sc_hd__nand4_1 _14565_ (.A(_06547_),
    .B(_06549_),
    .C(_06428_),
    .D(_06745_),
    .Y(_07049_));
 sky130_fd_sc_hd__a22o_1 _14566_ (.A1(_06930_),
    .A2(_06427_),
    .B1(_06745_),
    .B2(_06929_),
    .X(_07050_));
 sky130_fd_sc_hd__and2_1 _14567_ (.A(_06544_),
    .B(_06415_),
    .X(_07051_));
 sky130_fd_sc_hd__nand3_1 _14568_ (.A(_07049_),
    .B(_07050_),
    .C(_07051_),
    .Y(_07052_));
 sky130_fd_sc_hd__a21o_1 _14569_ (.A1(_07049_),
    .A2(_07050_),
    .B1(_07051_),
    .X(_07053_));
 sky130_fd_sc_hd__o21bai_1 _14570_ (.A1(_07030_),
    .A2(_07031_),
    .B1_N(_07029_),
    .Y(_07054_));
 sky130_fd_sc_hd__nand3_2 _14571_ (.A(_07052_),
    .B(_07053_),
    .C(_07054_),
    .Y(_07055_));
 sky130_fd_sc_hd__and3_1 _14572_ (.A(_06538_),
    .B(_06539_),
    .C(_06440_),
    .X(_07056_));
 sky130_fd_sc_hd__a22o_1 _14573_ (.A1(_06539_),
    .A2(_06440_),
    .B1(_06442_),
    .B2(_06538_),
    .X(_07057_));
 sky130_fd_sc_hd__a21bo_1 _14574_ (.A1(_06443_),
    .A2(_07056_),
    .B1_N(_07057_),
    .X(_07058_));
 sky130_fd_sc_hd__nand2_1 _14575_ (.A(_06604_),
    .B(_06423_),
    .Y(_07059_));
 sky130_fd_sc_hd__xor2_1 _14576_ (.A(_07058_),
    .B(_07059_),
    .X(_07060_));
 sky130_fd_sc_hd__a21o_1 _14577_ (.A1(_07052_),
    .A2(_07053_),
    .B1(_07054_),
    .X(_07061_));
 sky130_fd_sc_hd__nand3_2 _14578_ (.A(_07055_),
    .B(_07060_),
    .C(_07061_),
    .Y(_07062_));
 sky130_fd_sc_hd__a21bo_1 _14579_ (.A1(_06981_),
    .A2(_06986_),
    .B1_N(_06980_),
    .X(_07063_));
 sky130_fd_sc_hd__a21o_1 _14580_ (.A1(_07055_),
    .A2(_07061_),
    .B1(_07060_),
    .X(_07064_));
 sky130_fd_sc_hd__and3_1 _14581_ (.A(_07062_),
    .B(_07063_),
    .C(_07064_),
    .X(_07065_));
 sky130_fd_sc_hd__a21oi_1 _14582_ (.A1(_07062_),
    .A2(_07064_),
    .B1(_07063_),
    .Y(_07066_));
 sky130_fd_sc_hd__a211oi_2 _14583_ (.A1(_07038_),
    .A2(_07048_),
    .B1(_07065_),
    .C1(_07066_),
    .Y(_07067_));
 sky130_fd_sc_hd__o211a_1 _14584_ (.A1(_07065_),
    .A2(_07066_),
    .B1(_07038_),
    .C1(_07048_),
    .X(_07068_));
 sky130_fd_sc_hd__or4_4 _14585_ (.A(_07026_),
    .B(_07028_),
    .C(_07067_),
    .D(_07068_),
    .X(_07069_));
 sky130_fd_sc_hd__inv_2 _14586_ (.A(_07011_),
    .Y(_07070_));
 sky130_fd_sc_hd__nand2_1 _14587_ (.A(_07010_),
    .B(_07070_),
    .Y(_07071_));
 sky130_fd_sc_hd__nand4_1 _14588_ (.A(_06405_),
    .B(_06459_),
    .C(_06974_),
    .D(_06975_),
    .Y(_07072_));
 sky130_fd_sc_hd__a22o_1 _14589_ (.A1(\wfg_stim_sine_top.gain_val_q[14] ),
    .A2(_06973_),
    .B1(_06975_),
    .B2(_06458_),
    .X(_07073_));
 sky130_fd_sc_hd__and2_1 _14590_ (.A(\wfg_stim_sine_top.gain_val_q[13] ),
    .B(_06971_),
    .X(_07074_));
 sky130_fd_sc_hd__nand3_1 _14591_ (.A(_07072_),
    .B(_07073_),
    .C(_07074_),
    .Y(_07075_));
 sky130_fd_sc_hd__a22o_1 _14592_ (.A1(_06419_),
    .A2(_06971_),
    .B1(_07072_),
    .B2(_07073_),
    .X(_07076_));
 sky130_fd_sc_hd__nor2_1 _14593_ (.A(_06674_),
    .B(_07001_),
    .Y(_07077_));
 sky130_fd_sc_hd__nand3_1 _14594_ (.A(_07075_),
    .B(_07076_),
    .C(_07077_),
    .Y(_07078_));
 sky130_fd_sc_hd__a21o_1 _14595_ (.A1(_07075_),
    .A2(_07076_),
    .B1(_07077_),
    .X(_07079_));
 sky130_fd_sc_hd__and3_1 _14596_ (.A(\wfg_stim_sine_top.gain_val_q[12] ),
    .B(_06438_),
    .C(_06982_),
    .X(_07080_));
 sky130_fd_sc_hd__a22o_1 _14597_ (.A1(_06438_),
    .A2(_06896_),
    .B1(_06982_),
    .B2(\wfg_stim_sine_top.gain_val_q[12] ),
    .X(_07081_));
 sky130_fd_sc_hd__a21bo_1 _14598_ (.A1(_07007_),
    .A2(_07080_),
    .B1_N(_07081_),
    .X(_07082_));
 sky130_fd_sc_hd__nand2_1 _14599_ (.A(_06450_),
    .B(_06752_),
    .Y(_07083_));
 sky130_fd_sc_hd__xor2_1 _14600_ (.A(_07082_),
    .B(_07083_),
    .X(_07084_));
 sky130_fd_sc_hd__nand3_1 _14601_ (.A(_07078_),
    .B(_07079_),
    .C(_07084_),
    .Y(_07085_));
 sky130_fd_sc_hd__a21o_1 _14602_ (.A1(_07078_),
    .A2(_07079_),
    .B1(_07084_),
    .X(_07086_));
 sky130_fd_sc_hd__and2b_1 _14603_ (.A_N(_07003_),
    .B(_07009_),
    .X(_07087_));
 sky130_fd_sc_hd__nand3_4 _14604_ (.A(_07085_),
    .B(_07086_),
    .C(_07087_),
    .Y(_07088_));
 sky130_fd_sc_hd__a21o_1 _14605_ (.A1(_07085_),
    .A2(_07086_),
    .B1(_07087_),
    .X(_07089_));
 sky130_fd_sc_hd__or2b_1 _14606_ (.A(_07014_),
    .B_N(_07017_),
    .X(_07090_));
 sky130_fd_sc_hd__and4_1 _14607_ (.A(_06713_),
    .B(\wfg_stim_sine_top.gain_val_q[8] ),
    .C(_06737_),
    .D(_06738_),
    .X(_07091_));
 sky130_fd_sc_hd__a22oi_1 _14608_ (.A1(_06488_),
    .A2(_06737_),
    .B1(_06739_),
    .B2(_06713_),
    .Y(_07092_));
 sky130_fd_sc_hd__nand2_1 _14609_ (.A(_06484_),
    .B(_06745_),
    .Y(_07093_));
 sky130_fd_sc_hd__or3_1 _14610_ (.A(_07091_),
    .B(_07092_),
    .C(_07093_),
    .X(_07094_));
 sky130_fd_sc_hd__o21bai_1 _14611_ (.A1(_07004_),
    .A2(_07008_),
    .B1_N(_07005_),
    .Y(_07095_));
 sky130_fd_sc_hd__o21ai_1 _14612_ (.A1(_07091_),
    .A2(_07092_),
    .B1(_07093_),
    .Y(_07096_));
 sky130_fd_sc_hd__nand3_1 _14613_ (.A(_07094_),
    .B(_07095_),
    .C(_07096_),
    .Y(_07097_));
 sky130_fd_sc_hd__a21o_1 _14614_ (.A1(_07094_),
    .A2(_07096_),
    .B1(_07095_),
    .X(_07098_));
 sky130_fd_sc_hd__and3_1 _14615_ (.A(_07090_),
    .B(_07097_),
    .C(_07098_),
    .X(_07099_));
 sky130_fd_sc_hd__a21oi_1 _14616_ (.A1(_07097_),
    .A2(_07098_),
    .B1(_07090_),
    .Y(_07100_));
 sky130_fd_sc_hd__nor2_1 _14617_ (.A(_07099_),
    .B(_07100_),
    .Y(_07101_));
 sky130_fd_sc_hd__and3_1 _14618_ (.A(_07088_),
    .B(_07089_),
    .C(_07101_),
    .X(_07102_));
 sky130_fd_sc_hd__a21oi_2 _14619_ (.A1(_07088_),
    .A2(_07089_),
    .B1(_07101_),
    .Y(_07103_));
 sky130_fd_sc_hd__a211oi_4 _14620_ (.A1(_07071_),
    .A2(_07025_),
    .B1(_07102_),
    .C1(_07103_),
    .Y(_07104_));
 sky130_fd_sc_hd__o211a_1 _14621_ (.A1(_07102_),
    .A2(_07103_),
    .B1(_07071_),
    .C1(_07025_),
    .X(_07105_));
 sky130_fd_sc_hd__and4_1 _14622_ (.A(_06929_),
    .B(_06930_),
    .C(_06415_),
    .D(_06427_),
    .X(_07106_));
 sky130_fd_sc_hd__a22oi_2 _14623_ (.A1(_06930_),
    .A2(_06415_),
    .B1(_06428_),
    .B2(_06929_),
    .Y(_07107_));
 sky130_fd_sc_hd__nand2_1 _14624_ (.A(_06544_),
    .B(_06413_),
    .Y(_07108_));
 sky130_fd_sc_hd__or3_1 _14625_ (.A(_07106_),
    .B(_07107_),
    .C(_07108_),
    .X(_07109_));
 sky130_fd_sc_hd__o21ai_1 _14626_ (.A1(_07106_),
    .A2(_07107_),
    .B1(_07108_),
    .Y(_07110_));
 sky130_fd_sc_hd__a21bo_1 _14627_ (.A1(_07050_),
    .A2(_07051_),
    .B1_N(_07049_),
    .X(_07111_));
 sky130_fd_sc_hd__nand3_2 _14628_ (.A(_07109_),
    .B(_07110_),
    .C(_07111_),
    .Y(_07112_));
 sky130_fd_sc_hd__a22o_1 _14629_ (.A1(_07043_),
    .A2(_06452_),
    .B1(_06440_),
    .B2(_07044_),
    .X(_07113_));
 sky130_fd_sc_hd__a21bo_1 _14630_ (.A1(_06452_),
    .A2(_07056_),
    .B1_N(_07113_),
    .X(_07114_));
 sky130_fd_sc_hd__nand2_1 _14631_ (.A(_06604_),
    .B(_06463_),
    .Y(_07115_));
 sky130_fd_sc_hd__xor2_1 _14632_ (.A(_07114_),
    .B(_07115_),
    .X(_07116_));
 sky130_fd_sc_hd__a21o_1 _14633_ (.A1(_07109_),
    .A2(_07110_),
    .B1(_07111_),
    .X(_07117_));
 sky130_fd_sc_hd__nand3_2 _14634_ (.A(_07112_),
    .B(_07116_),
    .C(_07117_),
    .Y(_07118_));
 sky130_fd_sc_hd__a21o_1 _14635_ (.A1(_07013_),
    .A2(_07021_),
    .B1(_07020_),
    .X(_07119_));
 sky130_fd_sc_hd__a21o_1 _14636_ (.A1(_07112_),
    .A2(_07117_),
    .B1(_07116_),
    .X(_07120_));
 sky130_fd_sc_hd__and3_2 _14637_ (.A(_07118_),
    .B(_07119_),
    .C(_07120_),
    .X(_07121_));
 sky130_fd_sc_hd__a21oi_2 _14638_ (.A1(_07118_),
    .A2(_07120_),
    .B1(_07119_),
    .Y(_07122_));
 sky130_fd_sc_hd__a211oi_4 _14639_ (.A1(_07055_),
    .A2(_07062_),
    .B1(_07121_),
    .C1(_07122_),
    .Y(_07123_));
 sky130_fd_sc_hd__o211a_1 _14640_ (.A1(_07121_),
    .A2(_07122_),
    .B1(_07055_),
    .C1(_07062_),
    .X(_07124_));
 sky130_fd_sc_hd__nor4_4 _14641_ (.A(_07104_),
    .B(_07105_),
    .C(_07123_),
    .D(_07124_),
    .Y(_07125_));
 sky130_fd_sc_hd__o22a_1 _14642_ (.A1(_07104_),
    .A2(_07105_),
    .B1(_07123_),
    .B2(_07124_),
    .X(_07126_));
 sky130_fd_sc_hd__a211oi_4 _14643_ (.A1(_07027_),
    .A2(_07069_),
    .B1(_07125_),
    .C1(_07126_),
    .Y(_07127_));
 sky130_fd_sc_hd__o211a_1 _14644_ (.A1(_07125_),
    .A2(_07126_),
    .B1(_07027_),
    .C1(_07069_),
    .X(_07128_));
 sky130_fd_sc_hd__o2bb2a_1 _14645_ (.A1_N(_06513_),
    .A2_N(_07056_),
    .B1(_07058_),
    .B2(_07059_),
    .X(_07129_));
 sky130_fd_sc_hd__o21ba_1 _14646_ (.A1(_07065_),
    .A2(_07067_),
    .B1_N(_07129_),
    .X(_07130_));
 sky130_fd_sc_hd__or3b_1 _14647_ (.A(_07065_),
    .B(_07067_),
    .C_N(_07129_),
    .X(_07131_));
 sky130_fd_sc_hd__and2b_1 _14648_ (.A_N(_07130_),
    .B(_07131_),
    .X(_07132_));
 sky130_fd_sc_hd__nand2_1 _14649_ (.A(_06599_),
    .B(_06423_),
    .Y(_07133_));
 sky130_fd_sc_hd__xor2_1 _14650_ (.A(_07132_),
    .B(_07133_),
    .X(_07134_));
 sky130_fd_sc_hd__nor3_1 _14651_ (.A(_07127_),
    .B(_07128_),
    .C(_07134_),
    .Y(_07135_));
 sky130_fd_sc_hd__nand3_2 _14652_ (.A(_07088_),
    .B(_07089_),
    .C(_07101_),
    .Y(_07136_));
 sky130_fd_sc_hd__and4_1 _14653_ (.A(\wfg_stim_sine_top.gain_val_q[15] ),
    .B(\wfg_stim_sine_top.gain_val_q[14] ),
    .C(_06971_),
    .D(_06973_),
    .X(_07137_));
 sky130_fd_sc_hd__a22oi_2 _14654_ (.A1(_06459_),
    .A2(_06971_),
    .B1(_06974_),
    .B2(_06458_),
    .Y(_07138_));
 sky130_fd_sc_hd__nand2_1 _14655_ (.A(\wfg_stim_sine_top.gain_val_q[13] ),
    .B(_06996_),
    .Y(_07139_));
 sky130_fd_sc_hd__or3_1 _14656_ (.A(_07137_),
    .B(_07138_),
    .C(_07139_),
    .X(_07140_));
 sky130_fd_sc_hd__o21ai_1 _14657_ (.A1(_07137_),
    .A2(_07138_),
    .B1(_07139_),
    .Y(_07141_));
 sky130_fd_sc_hd__a21bo_1 _14658_ (.A1(_07073_),
    .A2(_07074_),
    .B1_N(_07072_),
    .X(_07142_));
 sky130_fd_sc_hd__nand3_1 _14659_ (.A(_07140_),
    .B(_07141_),
    .C(_07142_),
    .Y(_07143_));
 sky130_fd_sc_hd__a21o_1 _14660_ (.A1(_07140_),
    .A2(_07141_),
    .B1(_07142_),
    .X(_07144_));
 sky130_fd_sc_hd__a22oi_1 _14661_ (.A1(_06447_),
    .A2(_06752_),
    .B1(_07007_),
    .B2(_06444_),
    .Y(_07145_));
 sky130_fd_sc_hd__and4_1 _14662_ (.A(\wfg_stim_sine_top.gain_val_q[12] ),
    .B(_06438_),
    .C(_06894_),
    .D(_06896_),
    .X(_07146_));
 sky130_fd_sc_hd__nor2_1 _14663_ (.A(_07145_),
    .B(_07146_),
    .Y(_07147_));
 sky130_fd_sc_hd__nand2_1 _14664_ (.A(_06450_),
    .B(_06742_),
    .Y(_07148_));
 sky130_fd_sc_hd__xnor2_1 _14665_ (.A(_07147_),
    .B(_07148_),
    .Y(_07149_));
 sky130_fd_sc_hd__nand3_1 _14666_ (.A(_07143_),
    .B(_07144_),
    .C(_07149_),
    .Y(_07150_));
 sky130_fd_sc_hd__a21o_1 _14667_ (.A1(_07143_),
    .A2(_07144_),
    .B1(_07149_),
    .X(_07151_));
 sky130_fd_sc_hd__a21bo_1 _14668_ (.A1(_07079_),
    .A2(_07084_),
    .B1_N(_07078_),
    .X(_07152_));
 sky130_fd_sc_hd__nand3_4 _14669_ (.A(_07150_),
    .B(_07151_),
    .C(_07152_),
    .Y(_07153_));
 sky130_fd_sc_hd__a21o_1 _14670_ (.A1(_07150_),
    .A2(_07151_),
    .B1(_07152_),
    .X(_07154_));
 sky130_fd_sc_hd__or2b_1 _14671_ (.A(_07091_),
    .B_N(_07094_),
    .X(_07155_));
 sky130_fd_sc_hd__and4_1 _14672_ (.A(_06713_),
    .B(_06488_),
    .C(_06747_),
    .D(_06737_),
    .X(_07156_));
 sky130_fd_sc_hd__a22oi_1 _14673_ (.A1(_06488_),
    .A2(_06747_),
    .B1(_06741_),
    .B2(_06713_),
    .Y(_07157_));
 sky130_fd_sc_hd__nand2_1 _14674_ (.A(_06484_),
    .B(_06428_),
    .Y(_07158_));
 sky130_fd_sc_hd__or3_1 _14675_ (.A(_07156_),
    .B(_07157_),
    .C(_07158_),
    .X(_07159_));
 sky130_fd_sc_hd__a32o_1 _14676_ (.A1(_06450_),
    .A2(_06752_),
    .A3(_07081_),
    .B1(_07080_),
    .B2(_07007_),
    .X(_07160_));
 sky130_fd_sc_hd__o21ai_1 _14677_ (.A1(_07156_),
    .A2(_07157_),
    .B1(_07158_),
    .Y(_07161_));
 sky130_fd_sc_hd__and3_1 _14678_ (.A(_07159_),
    .B(_07160_),
    .C(_07161_),
    .X(_07162_));
 sky130_fd_sc_hd__a21o_1 _14679_ (.A1(_07159_),
    .A2(_07161_),
    .B1(_07160_),
    .X(_07163_));
 sky130_fd_sc_hd__and2b_1 _14680_ (.A_N(_07162_),
    .B(_07163_),
    .X(_07164_));
 sky130_fd_sc_hd__xor2_2 _14681_ (.A(_07155_),
    .B(_07164_),
    .X(_07165_));
 sky130_fd_sc_hd__and3_1 _14682_ (.A(_07153_),
    .B(_07154_),
    .C(_07165_),
    .X(_07166_));
 sky130_fd_sc_hd__a21oi_2 _14683_ (.A1(_07153_),
    .A2(_07154_),
    .B1(_07165_),
    .Y(_07167_));
 sky130_fd_sc_hd__a211oi_4 _14684_ (.A1(_07088_),
    .A2(_07136_),
    .B1(_07166_),
    .C1(_07167_),
    .Y(_07168_));
 sky130_fd_sc_hd__and4_1 _14685_ (.A(_06546_),
    .B(_06548_),
    .C(\wfg_stim_sine_top.wfg_stim_sine.sin_17[11] ),
    .D(\wfg_stim_sine_top.wfg_stim_sine.sin_17[10] ),
    .X(_07169_));
 sky130_fd_sc_hd__a22oi_2 _14686_ (.A1(_06930_),
    .A2(_06413_),
    .B1(_06415_),
    .B2(_06929_),
    .Y(_07170_));
 sky130_fd_sc_hd__nand2_1 _14687_ (.A(_06544_),
    .B(_06421_),
    .Y(_07171_));
 sky130_fd_sc_hd__or3_1 _14688_ (.A(_07169_),
    .B(_07170_),
    .C(_07171_),
    .X(_07172_));
 sky130_fd_sc_hd__o21ai_1 _14689_ (.A1(_07169_),
    .A2(_07170_),
    .B1(_07171_),
    .Y(_07173_));
 sky130_fd_sc_hd__o21bai_1 _14690_ (.A1(_07107_),
    .A2(_07108_),
    .B1_N(_07106_),
    .Y(_07174_));
 sky130_fd_sc_hd__nand3_1 _14691_ (.A(_07172_),
    .B(_07173_),
    .C(_07174_),
    .Y(_07175_));
 sky130_fd_sc_hd__a22oi_1 _14692_ (.A1(_07043_),
    .A2(_06409_),
    .B1(_06452_),
    .B2(_07044_),
    .Y(_07176_));
 sky130_fd_sc_hd__and4_1 _14693_ (.A(_06538_),
    .B(_06539_),
    .C(_06409_),
    .D(_06452_),
    .X(_07177_));
 sky130_fd_sc_hd__nor2_1 _14694_ (.A(_07176_),
    .B(_07177_),
    .Y(_07178_));
 sky130_fd_sc_hd__nand2_1 _14695_ (.A(_06604_),
    .B(_06441_),
    .Y(_07179_));
 sky130_fd_sc_hd__xnor2_1 _14696_ (.A(_07178_),
    .B(_07179_),
    .Y(_07180_));
 sky130_fd_sc_hd__a21o_1 _14697_ (.A1(_07172_),
    .A2(_07173_),
    .B1(_07174_),
    .X(_07181_));
 sky130_fd_sc_hd__nand3_1 _14698_ (.A(_07175_),
    .B(_07180_),
    .C(_07181_),
    .Y(_07182_));
 sky130_fd_sc_hd__a21bo_1 _14699_ (.A1(_07090_),
    .A2(_07098_),
    .B1_N(_07097_),
    .X(_07183_));
 sky130_fd_sc_hd__a21o_1 _14700_ (.A1(_07175_),
    .A2(_07181_),
    .B1(_07180_),
    .X(_07184_));
 sky130_fd_sc_hd__and3_1 _14701_ (.A(_07182_),
    .B(_07183_),
    .C(_07184_),
    .X(_07185_));
 sky130_fd_sc_hd__a21oi_1 _14702_ (.A1(_07182_),
    .A2(_07184_),
    .B1(_07183_),
    .Y(_07186_));
 sky130_fd_sc_hd__a211oi_1 _14703_ (.A1(_07112_),
    .A2(_07118_),
    .B1(_07185_),
    .C1(_07186_),
    .Y(_07187_));
 sky130_fd_sc_hd__o211a_1 _14704_ (.A1(_07185_),
    .A2(_07186_),
    .B1(_07112_),
    .C1(_07118_),
    .X(_07188_));
 sky130_fd_sc_hd__or2_1 _14705_ (.A(_07187_),
    .B(_07188_),
    .X(_07189_));
 sky130_fd_sc_hd__o211ai_1 _14706_ (.A1(_07166_),
    .A2(_07167_),
    .B1(_07088_),
    .C1(_07136_),
    .Y(_07190_));
 sky130_fd_sc_hd__or3b_2 _14707_ (.A(_07168_),
    .B(_07189_),
    .C_N(_07190_),
    .X(_07191_));
 sky130_fd_sc_hd__a211o_1 _14708_ (.A1(_07088_),
    .A2(_07136_),
    .B1(_07166_),
    .C1(_07167_),
    .X(_07192_));
 sky130_fd_sc_hd__a21bo_1 _14709_ (.A1(_07192_),
    .A2(_07190_),
    .B1_N(_07189_),
    .X(_07193_));
 sky130_fd_sc_hd__o211ai_4 _14710_ (.A1(_07104_),
    .A2(_07125_),
    .B1(_07191_),
    .C1(_07193_),
    .Y(_07194_));
 sky130_fd_sc_hd__a211o_1 _14711_ (.A1(_07191_),
    .A2(_07193_),
    .B1(_07104_),
    .C1(_07125_),
    .X(_07195_));
 sky130_fd_sc_hd__a32oi_1 _14712_ (.A1(_06605_),
    .A2(_06513_),
    .A3(_07113_),
    .B1(_07056_),
    .B2(_06672_),
    .Y(_07196_));
 sky130_fd_sc_hd__o21bai_1 _14713_ (.A1(_07121_),
    .A2(_07123_),
    .B1_N(_07196_),
    .Y(_07197_));
 sky130_fd_sc_hd__or3b_1 _14714_ (.A(_07121_),
    .B(_07123_),
    .C_N(_07196_),
    .X(_07198_));
 sky130_fd_sc_hd__and2_1 _14715_ (.A(_07197_),
    .B(_07198_),
    .X(_07199_));
 sky130_fd_sc_hd__buf_4 _14716_ (.A(_06599_),
    .X(_07200_));
 sky130_fd_sc_hd__nand2_1 _14717_ (.A(_07200_),
    .B(_06513_),
    .Y(_07201_));
 sky130_fd_sc_hd__xnor2_1 _14718_ (.A(_07199_),
    .B(_07201_),
    .Y(_07202_));
 sky130_fd_sc_hd__nand3_2 _14719_ (.A(_07194_),
    .B(_07195_),
    .C(_07202_),
    .Y(_07203_));
 sky130_fd_sc_hd__a21o_1 _14720_ (.A1(_07194_),
    .A2(_07195_),
    .B1(_07202_),
    .X(_07204_));
 sky130_fd_sc_hd__o211ai_2 _14721_ (.A1(_07127_),
    .A2(_07135_),
    .B1(_07203_),
    .C1(_07204_),
    .Y(_07205_));
 sky130_fd_sc_hd__buf_6 _14722_ (.A(_07200_),
    .X(_07206_));
 sky130_fd_sc_hd__and3_1 _14723_ (.A(_07206_),
    .B(_06423_),
    .C(_07132_),
    .X(_07207_));
 sky130_fd_sc_hd__a211o_1 _14724_ (.A1(_07203_),
    .A2(_07204_),
    .B1(_07127_),
    .C1(_07135_),
    .X(_07208_));
 sky130_fd_sc_hd__o211ai_2 _14725_ (.A1(_07130_),
    .A2(_07207_),
    .B1(_07205_),
    .C1(_07208_),
    .Y(_07209_));
 sky130_fd_sc_hd__nand3_1 _14726_ (.A(_07206_),
    .B(_06513_),
    .C(_07199_),
    .Y(_07210_));
 sky130_fd_sc_hd__and3b_1 _14727_ (.A_N(_07189_),
    .B(_07190_),
    .C(_07192_),
    .X(_07211_));
 sky130_fd_sc_hd__and4_1 _14728_ (.A(\wfg_stim_sine_top.gain_val_q[6] ),
    .B(\wfg_stim_sine_top.gain_val_q[5] ),
    .C(\wfg_stim_sine_top.wfg_stim_sine.sin_17[12] ),
    .D(\wfg_stim_sine_top.wfg_stim_sine.sin_17[11] ),
    .X(_07212_));
 sky130_fd_sc_hd__a22oi_1 _14729_ (.A1(_06548_),
    .A2(\wfg_stim_sine_top.wfg_stim_sine.sin_17[12] ),
    .B1(\wfg_stim_sine_top.wfg_stim_sine.sin_17[11] ),
    .B2(_06546_),
    .Y(_07213_));
 sky130_fd_sc_hd__nand2_1 _14730_ (.A(\wfg_stim_sine_top.gain_val_q[4] ),
    .B(_06442_),
    .Y(_07214_));
 sky130_fd_sc_hd__or3_1 _14731_ (.A(_07212_),
    .B(_07213_),
    .C(_07214_),
    .X(_07215_));
 sky130_fd_sc_hd__o21ai_1 _14732_ (.A1(_07212_),
    .A2(_07213_),
    .B1(_07214_),
    .Y(_07216_));
 sky130_fd_sc_hd__o21bai_1 _14733_ (.A1(_07170_),
    .A2(_07171_),
    .B1_N(_07169_),
    .Y(_07217_));
 sky130_fd_sc_hd__nand3_1 _14734_ (.A(_07215_),
    .B(_07216_),
    .C(_07217_),
    .Y(_07218_));
 sky130_fd_sc_hd__nand2_1 _14735_ (.A(_06604_),
    .B(_06453_),
    .Y(_07219_));
 sky130_fd_sc_hd__xnor2_1 _14736_ (.A(_06541_),
    .B(_07219_),
    .Y(_07220_));
 sky130_fd_sc_hd__a21o_1 _14737_ (.A1(_07215_),
    .A2(_07216_),
    .B1(_07217_),
    .X(_07221_));
 sky130_fd_sc_hd__nand3_1 _14738_ (.A(_07218_),
    .B(_07220_),
    .C(_07221_),
    .Y(_07222_));
 sky130_fd_sc_hd__a21o_1 _14739_ (.A1(_07155_),
    .A2(_07163_),
    .B1(_07162_),
    .X(_07223_));
 sky130_fd_sc_hd__a21o_1 _14740_ (.A1(_07218_),
    .A2(_07221_),
    .B1(_07220_),
    .X(_07224_));
 sky130_fd_sc_hd__and3_1 _14741_ (.A(_07222_),
    .B(_07223_),
    .C(_07224_),
    .X(_07225_));
 sky130_fd_sc_hd__a21oi_1 _14742_ (.A1(_07222_),
    .A2(_07224_),
    .B1(_07223_),
    .Y(_07226_));
 sky130_fd_sc_hd__a211oi_1 _14743_ (.A1(_07175_),
    .A2(_07182_),
    .B1(_07225_),
    .C1(_07226_),
    .Y(_07227_));
 sky130_fd_sc_hd__o211a_1 _14744_ (.A1(_07225_),
    .A2(_07226_),
    .B1(_07175_),
    .C1(_07182_),
    .X(_07228_));
 sky130_fd_sc_hd__or2_1 _14745_ (.A(_07227_),
    .B(_07228_),
    .X(_07229_));
 sky130_fd_sc_hd__nand4_1 _14746_ (.A(_06458_),
    .B(_06459_),
    .C(_06996_),
    .D(_06971_),
    .Y(_07230_));
 sky130_fd_sc_hd__a22o_1 _14747_ (.A1(\wfg_stim_sine_top.gain_val_q[14] ),
    .A2(_06982_),
    .B1(_06971_),
    .B2(\wfg_stim_sine_top.gain_val_q[15] ),
    .X(_07231_));
 sky130_fd_sc_hd__and2_1 _14748_ (.A(\wfg_stim_sine_top.gain_val_q[13] ),
    .B(_06896_),
    .X(_07232_));
 sky130_fd_sc_hd__nand3_1 _14749_ (.A(_07230_),
    .B(_07231_),
    .C(_07232_),
    .Y(_07233_));
 sky130_fd_sc_hd__a22o_1 _14750_ (.A1(_06419_),
    .A2(_07007_),
    .B1(_07230_),
    .B2(_07231_),
    .X(_07234_));
 sky130_fd_sc_hd__o21bai_1 _14751_ (.A1(_07138_),
    .A2(_07139_),
    .B1_N(_07137_),
    .Y(_07235_));
 sky130_fd_sc_hd__nand3_1 _14752_ (.A(_07233_),
    .B(_07234_),
    .C(_07235_),
    .Y(_07236_));
 sky130_fd_sc_hd__a21o_1 _14753_ (.A1(_07233_),
    .A2(_07234_),
    .B1(_07235_),
    .X(_07237_));
 sky130_fd_sc_hd__a22oi_1 _14754_ (.A1(_06447_),
    .A2(_06739_),
    .B1(_06894_),
    .B2(_06446_),
    .Y(_07238_));
 sky130_fd_sc_hd__and4_1 _14755_ (.A(\wfg_stim_sine_top.gain_val_q[12] ),
    .B(_06438_),
    .C(_06739_),
    .D(_06894_),
    .X(_07239_));
 sky130_fd_sc_hd__nor2_1 _14756_ (.A(_07238_),
    .B(_07239_),
    .Y(_07240_));
 sky130_fd_sc_hd__nand2_1 _14757_ (.A(_06450_),
    .B(_06754_),
    .Y(_07241_));
 sky130_fd_sc_hd__xnor2_1 _14758_ (.A(_07240_),
    .B(_07241_),
    .Y(_07242_));
 sky130_fd_sc_hd__nand3_1 _14759_ (.A(_07236_),
    .B(_07237_),
    .C(_07242_),
    .Y(_07243_));
 sky130_fd_sc_hd__a21o_1 _14760_ (.A1(_07236_),
    .A2(_07237_),
    .B1(_07242_),
    .X(_07244_));
 sky130_fd_sc_hd__a21bo_1 _14761_ (.A1(_07144_),
    .A2(_07149_),
    .B1_N(_07143_),
    .X(_07245_));
 sky130_fd_sc_hd__nand3_2 _14762_ (.A(_07243_),
    .B(_07244_),
    .C(_07245_),
    .Y(_07246_));
 sky130_fd_sc_hd__a21o_1 _14763_ (.A1(_07243_),
    .A2(_07244_),
    .B1(_07245_),
    .X(_07247_));
 sky130_fd_sc_hd__or2b_1 _14764_ (.A(_07156_),
    .B_N(_07159_),
    .X(_07248_));
 sky130_fd_sc_hd__and4_1 _14765_ (.A(_06713_),
    .B(_06488_),
    .C(_06427_),
    .D(_06747_),
    .X(_07249_));
 sky130_fd_sc_hd__a22oi_1 _14766_ (.A1(_06490_),
    .A2(_06427_),
    .B1(_06745_),
    .B2(_06487_),
    .Y(_07250_));
 sky130_fd_sc_hd__nand2_1 _14767_ (.A(_06484_),
    .B(_06415_),
    .Y(_07251_));
 sky130_fd_sc_hd__or3_1 _14768_ (.A(_07249_),
    .B(_07250_),
    .C(_07251_),
    .X(_07252_));
 sky130_fd_sc_hd__o21bai_1 _14769_ (.A1(_07145_),
    .A2(_07148_),
    .B1_N(_07146_),
    .Y(_07253_));
 sky130_fd_sc_hd__o21ai_1 _14770_ (.A1(_07249_),
    .A2(_07250_),
    .B1(_07251_),
    .Y(_07254_));
 sky130_fd_sc_hd__and3_1 _14771_ (.A(_07252_),
    .B(_07253_),
    .C(_07254_),
    .X(_07255_));
 sky130_fd_sc_hd__a21o_1 _14772_ (.A1(_07252_),
    .A2(_07254_),
    .B1(_07253_),
    .X(_07256_));
 sky130_fd_sc_hd__or2b_1 _14773_ (.A(_07255_),
    .B_N(_07256_),
    .X(_07257_));
 sky130_fd_sc_hd__xnor2_1 _14774_ (.A(_07248_),
    .B(_07257_),
    .Y(_07258_));
 sky130_fd_sc_hd__and3_1 _14775_ (.A(_07246_),
    .B(_07247_),
    .C(_07258_),
    .X(_07259_));
 sky130_fd_sc_hd__a21oi_2 _14776_ (.A1(_07246_),
    .A2(_07247_),
    .B1(_07258_),
    .Y(_07260_));
 sky130_fd_sc_hd__nand3_2 _14777_ (.A(_07153_),
    .B(_07154_),
    .C(_07165_),
    .Y(_07261_));
 sky130_fd_sc_hd__o211ai_4 _14778_ (.A1(_07259_),
    .A2(_07260_),
    .B1(_07153_),
    .C1(_07261_),
    .Y(_07262_));
 sky130_fd_sc_hd__a211o_2 _14779_ (.A1(_07153_),
    .A2(_07261_),
    .B1(_07259_),
    .C1(_07260_),
    .X(_07263_));
 sky130_fd_sc_hd__nand3b_4 _14780_ (.A_N(_07229_),
    .B(_07262_),
    .C(_07263_),
    .Y(_07264_));
 sky130_fd_sc_hd__a21bo_1 _14781_ (.A1(_07263_),
    .A2(_07262_),
    .B1_N(_07229_),
    .X(_07265_));
 sky130_fd_sc_hd__o211ai_4 _14782_ (.A1(_07168_),
    .A2(_07211_),
    .B1(_07264_),
    .C1(_07265_),
    .Y(_07266_));
 sky130_fd_sc_hd__a211o_1 _14783_ (.A1(_07264_),
    .A2(_07265_),
    .B1(_07168_),
    .C1(_07211_),
    .X(_07267_));
 sky130_fd_sc_hd__or2_1 _14784_ (.A(_07185_),
    .B(_07187_),
    .X(_07268_));
 sky130_fd_sc_hd__and3_1 _14785_ (.A(_06605_),
    .B(_06510_),
    .C(_07178_),
    .X(_07269_));
 sky130_fd_sc_hd__nor2_1 _14786_ (.A(_07177_),
    .B(_07269_),
    .Y(_07270_));
 sky130_fd_sc_hd__xnor2_1 _14787_ (.A(_07268_),
    .B(_07270_),
    .Y(_07271_));
 sky130_fd_sc_hd__nand2_1 _14788_ (.A(_07200_),
    .B(_06510_),
    .Y(_07272_));
 sky130_fd_sc_hd__xnor2_1 _14789_ (.A(_07271_),
    .B(_07272_),
    .Y(_07273_));
 sky130_fd_sc_hd__and3_1 _14790_ (.A(_07266_),
    .B(_07267_),
    .C(_07273_),
    .X(_07274_));
 sky130_fd_sc_hd__a21oi_1 _14791_ (.A1(_07266_),
    .A2(_07267_),
    .B1(_07273_),
    .Y(_07275_));
 sky130_fd_sc_hd__a211oi_2 _14792_ (.A1(_07194_),
    .A2(_07203_),
    .B1(_07274_),
    .C1(_07275_),
    .Y(_07276_));
 sky130_fd_sc_hd__o211a_1 _14793_ (.A1(_07274_),
    .A2(_07275_),
    .B1(_07194_),
    .C1(_07203_),
    .X(_07277_));
 sky130_fd_sc_hd__a211oi_2 _14794_ (.A1(_07197_),
    .A2(_07210_),
    .B1(_07276_),
    .C1(_07277_),
    .Y(_07278_));
 sky130_fd_sc_hd__o211a_1 _14795_ (.A1(_07276_),
    .A2(_07277_),
    .B1(_07197_),
    .C1(_07210_),
    .X(_07279_));
 sky130_fd_sc_hd__a211oi_1 _14796_ (.A1(_07205_),
    .A2(_07209_),
    .B1(_07278_),
    .C1(_07279_),
    .Y(_07280_));
 sky130_fd_sc_hd__inv_2 _14797_ (.A(_07280_),
    .Y(_07281_));
 sky130_fd_sc_hd__a21o_1 _14798_ (.A1(_06987_),
    .A2(_06988_),
    .B1(_06999_),
    .X(_07282_));
 sky130_fd_sc_hd__a22o_1 _14799_ (.A1(_06485_),
    .A2(_06752_),
    .B1(_06983_),
    .B2(_06984_),
    .X(_07283_));
 sky130_fd_sc_hd__and4_1 _14800_ (.A(_06439_),
    .B(\wfg_stim_sine_top.gain_val_q[10] ),
    .C(_06974_),
    .D(_06989_),
    .X(_07284_));
 sky130_fd_sc_hd__nand3_2 _14801_ (.A(_06985_),
    .B(_07283_),
    .C(_07284_),
    .Y(_07285_));
 sky130_fd_sc_hd__a21o_1 _14802_ (.A1(_06985_),
    .A2(_07283_),
    .B1(_07284_),
    .X(_07286_));
 sky130_fd_sc_hd__and4_1 _14803_ (.A(\wfg_stim_sine_top.gain_val_q[9] ),
    .B(\wfg_stim_sine_top.gain_val_q[8] ),
    .C(\wfg_stim_sine_top.wfg_stim_sine.sin_17[3] ),
    .D(_06970_),
    .X(_07287_));
 sky130_fd_sc_hd__a22oi_1 _14804_ (.A1(\wfg_stim_sine_top.gain_val_q[8] ),
    .A2(_06995_),
    .B1(_06991_),
    .B2(_06713_),
    .Y(_07288_));
 sky130_fd_sc_hd__nor2_1 _14805_ (.A(_07287_),
    .B(_07288_),
    .Y(_07289_));
 sky130_fd_sc_hd__a31o_1 _14806_ (.A1(_06486_),
    .A2(_07007_),
    .A3(_07289_),
    .B1(_07287_),
    .X(_07290_));
 sky130_fd_sc_hd__nand3_1 _14807_ (.A(_07285_),
    .B(_07286_),
    .C(_07290_),
    .Y(_07291_));
 sky130_fd_sc_hd__a21o_1 _14808_ (.A1(_07285_),
    .A2(_07286_),
    .B1(_07290_),
    .X(_07292_));
 sky130_fd_sc_hd__nand2_1 _14809_ (.A(_06468_),
    .B(_06972_),
    .Y(_07293_));
 sky130_fd_sc_hd__and2b_1 _14810_ (.A_N(_06977_),
    .B(_06976_),
    .X(_07294_));
 sky130_fd_sc_hd__xnor2_2 _14811_ (.A(_07293_),
    .B(_07294_),
    .Y(_07295_));
 sky130_fd_sc_hd__and3_1 _14812_ (.A(_07291_),
    .B(_07292_),
    .C(_07295_),
    .X(_07296_));
 sky130_fd_sc_hd__and3_2 _14813_ (.A(_07000_),
    .B(_07282_),
    .C(_07296_),
    .X(_07297_));
 sky130_fd_sc_hd__nand3_1 _14814_ (.A(_07036_),
    .B(_07034_),
    .C(_07035_),
    .Y(_07298_));
 sky130_fd_sc_hd__a22o_1 _14815_ (.A1(_06544_),
    .A2(_06748_),
    .B1(_07036_),
    .B2(_07035_),
    .X(_07299_));
 sky130_fd_sc_hd__nand2_1 _14816_ (.A(\wfg_stim_sine_top.gain_val_q[4] ),
    .B(_06737_),
    .Y(_07300_));
 sky130_fd_sc_hd__a22oi_2 _14817_ (.A1(\wfg_stim_sine_top.gain_val_q[5] ),
    .A2(_06738_),
    .B1(_06750_),
    .B2(\wfg_stim_sine_top.gain_val_q[6] ),
    .Y(_07301_));
 sky130_fd_sc_hd__and4_1 _14818_ (.A(\wfg_stim_sine_top.gain_val_q[6] ),
    .B(\wfg_stim_sine_top.gain_val_q[5] ),
    .C(_06738_),
    .D(\wfg_stim_sine_top.wfg_stim_sine.sin_17[5] ),
    .X(_07302_));
 sky130_fd_sc_hd__o21bai_1 _14819_ (.A1(_07300_),
    .A2(_07301_),
    .B1_N(_07302_),
    .Y(_07303_));
 sky130_fd_sc_hd__nand3_2 _14820_ (.A(_07298_),
    .B(_07299_),
    .C(_07303_),
    .Y(_07304_));
 sky130_fd_sc_hd__a21o_1 _14821_ (.A1(_07298_),
    .A2(_07299_),
    .B1(_07303_),
    .X(_07305_));
 sky130_fd_sc_hd__nand2_1 _14822_ (.A(_06604_),
    .B(_06770_),
    .Y(_07306_));
 sky130_fd_sc_hd__nand2_2 _14823_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[12] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.sin_17[11] ),
    .Y(_07307_));
 sky130_fd_sc_hd__a22o_1 _14824_ (.A1(_07043_),
    .A2(_06421_),
    .B1(_06414_),
    .B2(_07044_),
    .X(_07308_));
 sky130_fd_sc_hd__o21ai_1 _14825_ (.A1(_07041_),
    .A2(_07307_),
    .B1(_07308_),
    .Y(_07309_));
 sky130_fd_sc_hd__xor2_1 _14826_ (.A(_07306_),
    .B(_07309_),
    .X(_07310_));
 sky130_fd_sc_hd__nand3_2 _14827_ (.A(_07304_),
    .B(_07305_),
    .C(_07310_),
    .Y(_07311_));
 sky130_fd_sc_hd__a21bo_1 _14828_ (.A1(_07286_),
    .A2(_07290_),
    .B1_N(_07285_),
    .X(_07312_));
 sky130_fd_sc_hd__a21o_1 _14829_ (.A1(_07038_),
    .A2(_07039_),
    .B1(_07047_),
    .X(_07313_));
 sky130_fd_sc_hd__and3_1 _14830_ (.A(_07048_),
    .B(_07312_),
    .C(_07313_),
    .X(_07314_));
 sky130_fd_sc_hd__a21oi_2 _14831_ (.A1(_07048_),
    .A2(_07313_),
    .B1(_07312_),
    .Y(_07315_));
 sky130_fd_sc_hd__a211oi_4 _14832_ (.A1(_07304_),
    .A2(_07311_),
    .B1(_07314_),
    .C1(_07315_),
    .Y(_07316_));
 sky130_fd_sc_hd__o211a_1 _14833_ (.A1(_07314_),
    .A2(_07315_),
    .B1(_07304_),
    .C1(_07311_),
    .X(_07317_));
 sky130_fd_sc_hd__a21oi_2 _14834_ (.A1(_07000_),
    .A2(_07282_),
    .B1(_07296_),
    .Y(_07318_));
 sky130_fd_sc_hd__nor4_4 _14835_ (.A(_07297_),
    .B(_07316_),
    .C(_07317_),
    .D(_07318_),
    .Y(_07319_));
 sky130_fd_sc_hd__o22ai_2 _14836_ (.A1(_07026_),
    .A2(_07028_),
    .B1(_07067_),
    .B2(_07068_),
    .Y(_07320_));
 sky130_fd_sc_hd__o211a_1 _14837_ (.A1(_07297_),
    .A2(_07319_),
    .B1(_07069_),
    .C1(_07320_),
    .X(_07321_));
 sky130_fd_sc_hd__a211oi_2 _14838_ (.A1(_07069_),
    .A2(_07320_),
    .B1(_07297_),
    .C1(_07319_),
    .Y(_07322_));
 sky130_fd_sc_hd__or2_1 _14839_ (.A(_07314_),
    .B(_07316_),
    .X(_07323_));
 sky130_fd_sc_hd__buf_4 _14840_ (.A(_07041_),
    .X(_07324_));
 sky130_fd_sc_hd__o22a_1 _14841_ (.A1(_07324_),
    .A2(_07042_),
    .B1(_07046_),
    .B2(_07040_),
    .X(_07325_));
 sky130_fd_sc_hd__xnor2_1 _14842_ (.A(_07323_),
    .B(_07325_),
    .Y(_07326_));
 sky130_fd_sc_hd__nand2_1 _14843_ (.A(_06599_),
    .B(_06432_),
    .Y(_07327_));
 sky130_fd_sc_hd__xor2_1 _14844_ (.A(_07326_),
    .B(_07327_),
    .X(_07328_));
 sky130_fd_sc_hd__nor3_1 _14845_ (.A(_07321_),
    .B(_07322_),
    .C(_07328_),
    .Y(_07329_));
 sky130_fd_sc_hd__or3_1 _14846_ (.A(_07127_),
    .B(_07128_),
    .C(_07134_),
    .X(_07330_));
 sky130_fd_sc_hd__o21ai_1 _14847_ (.A1(_07127_),
    .A2(_07128_),
    .B1(_07134_),
    .Y(_07331_));
 sky130_fd_sc_hd__o211a_1 _14848_ (.A1(_07321_),
    .A2(_07329_),
    .B1(_07330_),
    .C1(_07331_),
    .X(_07332_));
 sky130_fd_sc_hd__a211o_1 _14849_ (.A1(_07330_),
    .A2(_07331_),
    .B1(_07321_),
    .C1(_07329_),
    .X(_07333_));
 sky130_fd_sc_hd__o21ba_1 _14850_ (.A1(_07314_),
    .A2(_07316_),
    .B1_N(_07325_),
    .X(_07334_));
 sky130_fd_sc_hd__a31o_1 _14851_ (.A1(_07206_),
    .A2(_06432_),
    .A3(_07326_),
    .B1(_07334_),
    .X(_07335_));
 sky130_fd_sc_hd__and3b_1 _14852_ (.A_N(_07332_),
    .B(_07333_),
    .C(_07335_),
    .X(_07336_));
 sky130_fd_sc_hd__nor2_1 _14853_ (.A(_07332_),
    .B(_07336_),
    .Y(_07337_));
 sky130_fd_sc_hd__a211o_1 _14854_ (.A1(_07205_),
    .A2(_07208_),
    .B1(_07130_),
    .C1(_07207_),
    .X(_07338_));
 sky130_fd_sc_hd__and2_1 _14855_ (.A(_07209_),
    .B(_07338_),
    .X(_07339_));
 sky130_fd_sc_hd__or2b_1 _14856_ (.A(_07337_),
    .B_N(_07339_),
    .X(_07340_));
 sky130_fd_sc_hd__o211a_1 _14857_ (.A1(_07278_),
    .A2(_07279_),
    .B1(_07205_),
    .C1(_07209_),
    .X(_07341_));
 sky130_fd_sc_hd__a21o_1 _14858_ (.A1(_07281_),
    .A2(_07340_),
    .B1(_07341_),
    .X(_07342_));
 sky130_fd_sc_hd__nand3_1 _14859_ (.A(_07266_),
    .B(_07267_),
    .C(_07273_),
    .Y(_07343_));
 sky130_fd_sc_hd__nand3_1 _14860_ (.A(_07246_),
    .B(_07247_),
    .C(_07258_),
    .Y(_07344_));
 sky130_fd_sc_hd__and4_1 _14861_ (.A(\wfg_stim_sine_top.gain_val_q[15] ),
    .B(\wfg_stim_sine_top.gain_val_q[14] ),
    .C(_06965_),
    .D(_06995_),
    .X(_07345_));
 sky130_fd_sc_hd__a22oi_2 _14862_ (.A1(\wfg_stim_sine_top.gain_val_q[14] ),
    .A2(_06965_),
    .B1(_06982_),
    .B2(\wfg_stim_sine_top.gain_val_q[15] ),
    .Y(_07346_));
 sky130_fd_sc_hd__nand2_1 _14863_ (.A(\wfg_stim_sine_top.gain_val_q[13] ),
    .B(_06894_),
    .Y(_07347_));
 sky130_fd_sc_hd__or3_1 _14864_ (.A(_07345_),
    .B(_07346_),
    .C(_07347_),
    .X(_07348_));
 sky130_fd_sc_hd__o21ai_1 _14865_ (.A1(_07345_),
    .A2(_07346_),
    .B1(_07347_),
    .Y(_07349_));
 sky130_fd_sc_hd__a21bo_1 _14866_ (.A1(_07231_),
    .A2(_07232_),
    .B1_N(_07230_),
    .X(_07350_));
 sky130_fd_sc_hd__nand3_1 _14867_ (.A(_07348_),
    .B(_07349_),
    .C(_07350_),
    .Y(_07351_));
 sky130_fd_sc_hd__a21o_1 _14868_ (.A1(_07348_),
    .A2(_07349_),
    .B1(_07350_),
    .X(_07352_));
 sky130_fd_sc_hd__a22oi_1 _14869_ (.A1(_06447_),
    .A2(_06741_),
    .B1(_06742_),
    .B2(_06446_),
    .Y(_07353_));
 sky130_fd_sc_hd__and4_1 _14870_ (.A(_06446_),
    .B(_06447_),
    .C(_06741_),
    .D(_06739_),
    .X(_07354_));
 sky130_fd_sc_hd__nor2_1 _14871_ (.A(_07353_),
    .B(_07354_),
    .Y(_07355_));
 sky130_fd_sc_hd__nand2_1 _14872_ (.A(_06450_),
    .B(_06748_),
    .Y(_07356_));
 sky130_fd_sc_hd__xnor2_1 _14873_ (.A(_07355_),
    .B(_07356_),
    .Y(_07357_));
 sky130_fd_sc_hd__nand3_1 _14874_ (.A(_07351_),
    .B(_07352_),
    .C(_07357_),
    .Y(_07358_));
 sky130_fd_sc_hd__a21o_1 _14875_ (.A1(_07351_),
    .A2(_07352_),
    .B1(_07357_),
    .X(_07359_));
 sky130_fd_sc_hd__a21bo_1 _14876_ (.A1(_07237_),
    .A2(_07242_),
    .B1_N(_07236_),
    .X(_07360_));
 sky130_fd_sc_hd__nand3_2 _14877_ (.A(_07358_),
    .B(_07359_),
    .C(_07360_),
    .Y(_07361_));
 sky130_fd_sc_hd__a21o_1 _14878_ (.A1(_07358_),
    .A2(_07359_),
    .B1(_07360_),
    .X(_07362_));
 sky130_fd_sc_hd__or2b_1 _14879_ (.A(_07249_),
    .B_N(_07252_),
    .X(_07363_));
 sky130_fd_sc_hd__a31o_1 _14880_ (.A1(_06450_),
    .A2(_06754_),
    .A3(_07240_),
    .B1(_07239_),
    .X(_07364_));
 sky130_fd_sc_hd__nand4_1 _14881_ (.A(_06487_),
    .B(_06490_),
    .C(_06416_),
    .D(_06428_),
    .Y(_07365_));
 sky130_fd_sc_hd__a22o_1 _14882_ (.A1(_06490_),
    .A2(_06415_),
    .B1(_06427_),
    .B2(_06487_),
    .X(_07366_));
 sky130_fd_sc_hd__nand4_1 _14883_ (.A(_06485_),
    .B(_06432_),
    .C(_07365_),
    .D(_07366_),
    .Y(_07367_));
 sky130_fd_sc_hd__a22o_1 _14884_ (.A1(_06485_),
    .A2(_06414_),
    .B1(_07365_),
    .B2(_07366_),
    .X(_07368_));
 sky130_fd_sc_hd__nand2_1 _14885_ (.A(_07367_),
    .B(_07368_),
    .Y(_07369_));
 sky130_fd_sc_hd__xnor2_1 _14886_ (.A(_07364_),
    .B(_07369_),
    .Y(_07370_));
 sky130_fd_sc_hd__xor2_1 _14887_ (.A(_07363_),
    .B(_07370_),
    .X(_07371_));
 sky130_fd_sc_hd__and3_1 _14888_ (.A(_07361_),
    .B(_07362_),
    .C(_07371_),
    .X(_07372_));
 sky130_fd_sc_hd__a21oi_1 _14889_ (.A1(_07361_),
    .A2(_07362_),
    .B1(_07371_),
    .Y(_07373_));
 sky130_fd_sc_hd__a211oi_2 _14890_ (.A1(_07246_),
    .A2(_07344_),
    .B1(_07372_),
    .C1(_07373_),
    .Y(_07374_));
 sky130_fd_sc_hd__o211a_1 _14891_ (.A1(_07372_),
    .A2(_07373_),
    .B1(_07246_),
    .C1(_07344_),
    .X(_07375_));
 sky130_fd_sc_hd__nand2_1 _14892_ (.A(_07218_),
    .B(_07222_),
    .Y(_07376_));
 sky130_fd_sc_hd__nand4_1 _14893_ (.A(_06547_),
    .B(_06549_),
    .C(_06443_),
    .D(_06422_),
    .Y(_07377_));
 sky130_fd_sc_hd__a22o_1 _14894_ (.A1(_06549_),
    .A2(_06442_),
    .B1(_06421_),
    .B2(_06547_),
    .X(_07378_));
 sky130_fd_sc_hd__nand4_1 _14895_ (.A(_06551_),
    .B(_06441_),
    .C(_07377_),
    .D(_07378_),
    .Y(_07379_));
 sky130_fd_sc_hd__a22o_1 _14896_ (.A1(_06551_),
    .A2(_06441_),
    .B1(_07377_),
    .B2(_07378_),
    .X(_07380_));
 sky130_fd_sc_hd__or2b_1 _14897_ (.A(_07212_),
    .B_N(_07215_),
    .X(_07381_));
 sky130_fd_sc_hd__nand3_2 _14898_ (.A(_07379_),
    .B(_07380_),
    .C(_07381_),
    .Y(_07382_));
 sky130_fd_sc_hd__a21o_1 _14899_ (.A1(_07379_),
    .A2(_07380_),
    .B1(_07381_),
    .X(_07383_));
 sky130_fd_sc_hd__and3_1 _14900_ (.A(_06648_),
    .B(_07382_),
    .C(_07383_),
    .X(_07384_));
 sky130_fd_sc_hd__a21oi_1 _14901_ (.A1(_07248_),
    .A2(_07256_),
    .B1(_07255_),
    .Y(_07385_));
 sky130_fd_sc_hd__a21oi_1 _14902_ (.A1(_07382_),
    .A2(_07383_),
    .B1(_06648_),
    .Y(_07386_));
 sky130_fd_sc_hd__or3_1 _14903_ (.A(_07384_),
    .B(_07385_),
    .C(_07386_),
    .X(_07387_));
 sky130_fd_sc_hd__o21ai_1 _14904_ (.A1(_07384_),
    .A2(_07386_),
    .B1(_07385_),
    .Y(_07388_));
 sky130_fd_sc_hd__and3_1 _14905_ (.A(_07376_),
    .B(_07387_),
    .C(_07388_),
    .X(_07389_));
 sky130_fd_sc_hd__a21oi_1 _14906_ (.A1(_07387_),
    .A2(_07388_),
    .B1(_07376_),
    .Y(_07390_));
 sky130_fd_sc_hd__nor4_1 _14907_ (.A(_07374_),
    .B(_07375_),
    .C(_07389_),
    .D(_07390_),
    .Y(_07391_));
 sky130_fd_sc_hd__o22a_1 _14908_ (.A1(_07374_),
    .A2(_07375_),
    .B1(_07389_),
    .B2(_07390_),
    .X(_07392_));
 sky130_fd_sc_hd__a211o_1 _14909_ (.A1(_07263_),
    .A2(_07264_),
    .B1(_07391_),
    .C1(_07392_),
    .X(_07393_));
 sky130_fd_sc_hd__o211ai_2 _14910_ (.A1(_07391_),
    .A2(_07392_),
    .B1(_07263_),
    .C1(_07264_),
    .Y(_07394_));
 sky130_fd_sc_hd__or2_1 _14911_ (.A(_07225_),
    .B(_07227_),
    .X(_07395_));
 sky130_fd_sc_hd__and3_1 _14912_ (.A(_06605_),
    .B(_06672_),
    .C(_06541_),
    .X(_07396_));
 sky130_fd_sc_hd__nor2_1 _14913_ (.A(_06537_),
    .B(_07396_),
    .Y(_07397_));
 sky130_fd_sc_hd__xnor2_1 _14914_ (.A(_07395_),
    .B(_07397_),
    .Y(_07398_));
 sky130_fd_sc_hd__nand2_1 _14915_ (.A(_07200_),
    .B(_06672_),
    .Y(_07399_));
 sky130_fd_sc_hd__xnor2_1 _14916_ (.A(_07398_),
    .B(_07399_),
    .Y(_07400_));
 sky130_fd_sc_hd__and3_1 _14917_ (.A(_07393_),
    .B(_07394_),
    .C(_07400_),
    .X(_07401_));
 sky130_fd_sc_hd__a21oi_1 _14918_ (.A1(_07393_),
    .A2(_07394_),
    .B1(_07400_),
    .Y(_07402_));
 sky130_fd_sc_hd__a211o_1 _14919_ (.A1(_07266_),
    .A2(_07343_),
    .B1(_07401_),
    .C1(_07402_),
    .X(_07403_));
 sky130_fd_sc_hd__o211ai_1 _14920_ (.A1(_07401_),
    .A2(_07402_),
    .B1(_07266_),
    .C1(_07343_),
    .Y(_07404_));
 sky130_fd_sc_hd__nand2_1 _14921_ (.A(_07403_),
    .B(_07404_),
    .Y(_07405_));
 sky130_fd_sc_hd__o21a_1 _14922_ (.A1(_07177_),
    .A2(_07269_),
    .B1(_07268_),
    .X(_07406_));
 sky130_fd_sc_hd__and3_1 _14923_ (.A(_07206_),
    .B(_06510_),
    .C(_07271_),
    .X(_07407_));
 sky130_fd_sc_hd__nor2_1 _14924_ (.A(_07406_),
    .B(_07407_),
    .Y(_07408_));
 sky130_fd_sc_hd__xnor2_1 _14925_ (.A(_07405_),
    .B(_07408_),
    .Y(_07409_));
 sky130_fd_sc_hd__nor2_1 _14926_ (.A(_07276_),
    .B(_07278_),
    .Y(_07410_));
 sky130_fd_sc_hd__xor2_1 _14927_ (.A(_07409_),
    .B(_07410_),
    .X(_07411_));
 sky130_fd_sc_hd__o211ai_1 _14928_ (.A1(_07406_),
    .A2(_07407_),
    .B1(_07403_),
    .C1(_07404_),
    .Y(_07412_));
 sky130_fd_sc_hd__o21ai_1 _14929_ (.A1(_06537_),
    .A2(_07396_),
    .B1(_07395_),
    .Y(_07413_));
 sky130_fd_sc_hd__nand3_1 _14930_ (.A(_07206_),
    .B(_06672_),
    .C(_07398_),
    .Y(_07414_));
 sky130_fd_sc_hd__nand3_1 _14931_ (.A(_07393_),
    .B(_07394_),
    .C(_07400_),
    .Y(_07415_));
 sky130_fd_sc_hd__inv_2 _14932_ (.A(_07374_),
    .Y(_07416_));
 sky130_fd_sc_hd__or4_1 _14933_ (.A(_07374_),
    .B(_07375_),
    .C(_07389_),
    .D(_07390_),
    .X(_07417_));
 sky130_fd_sc_hd__nand3_2 _14934_ (.A(_07361_),
    .B(_07362_),
    .C(_07371_),
    .Y(_07418_));
 sky130_fd_sc_hd__a22o_1 _14935_ (.A1(_06419_),
    .A2(_06742_),
    .B1(_06897_),
    .B2(_06898_),
    .X(_07419_));
 sky130_fd_sc_hd__o21bai_1 _14936_ (.A1(_07346_),
    .A2(_07347_),
    .B1_N(_07345_),
    .Y(_07420_));
 sky130_fd_sc_hd__nand3_2 _14937_ (.A(_06899_),
    .B(_07419_),
    .C(_07420_),
    .Y(_07421_));
 sky130_fd_sc_hd__a21o_1 _14938_ (.A1(_06899_),
    .A2(_07419_),
    .B1(_07420_),
    .X(_07422_));
 sky130_fd_sc_hd__and3_1 _14939_ (.A(_06446_),
    .B(_06447_),
    .C(_06741_),
    .X(_07423_));
 sky130_fd_sc_hd__a22o_1 _14940_ (.A1(_06447_),
    .A2(_06745_),
    .B1(_06741_),
    .B2(_06446_),
    .X(_07424_));
 sky130_fd_sc_hd__a21bo_1 _14941_ (.A1(_06748_),
    .A2(_07423_),
    .B1_N(_07424_),
    .X(_07425_));
 sky130_fd_sc_hd__nand2_1 _14942_ (.A(_06468_),
    .B(_06430_),
    .Y(_07426_));
 sky130_fd_sc_hd__xor2_1 _14943_ (.A(_07425_),
    .B(_07426_),
    .X(_07427_));
 sky130_fd_sc_hd__nand3_2 _14944_ (.A(_07421_),
    .B(_07422_),
    .C(_07427_),
    .Y(_07428_));
 sky130_fd_sc_hd__a21o_1 _14945_ (.A1(_07421_),
    .A2(_07422_),
    .B1(_07427_),
    .X(_07429_));
 sky130_fd_sc_hd__a21bo_1 _14946_ (.A1(_07352_),
    .A2(_07357_),
    .B1_N(_07351_),
    .X(_07430_));
 sky130_fd_sc_hd__and3_2 _14947_ (.A(_07428_),
    .B(_07429_),
    .C(_07430_),
    .X(_07431_));
 sky130_fd_sc_hd__a21oi_2 _14948_ (.A1(_07428_),
    .A2(_07429_),
    .B1(_07430_),
    .Y(_07432_));
 sky130_fd_sc_hd__and2_1 _14949_ (.A(_07365_),
    .B(_07367_),
    .X(_07433_));
 sky130_fd_sc_hd__and4_1 _14950_ (.A(_06487_),
    .B(_06490_),
    .C(_06413_),
    .D(_06416_),
    .X(_07434_));
 sky130_fd_sc_hd__a22oi_1 _14951_ (.A1(_06725_),
    .A2(_06414_),
    .B1(_06416_),
    .B2(_06714_),
    .Y(_07435_));
 sky130_fd_sc_hd__nand2_1 _14952_ (.A(_06485_),
    .B(_06422_),
    .Y(_07436_));
 sky130_fd_sc_hd__or3_1 _14953_ (.A(_07434_),
    .B(_07435_),
    .C(_07436_),
    .X(_07437_));
 sky130_fd_sc_hd__o21bai_1 _14954_ (.A1(_07353_),
    .A2(_07356_),
    .B1_N(_07354_),
    .Y(_07438_));
 sky130_fd_sc_hd__o21ai_1 _14955_ (.A1(_07434_),
    .A2(_07435_),
    .B1(_07436_),
    .Y(_07439_));
 sky130_fd_sc_hd__and3_1 _14956_ (.A(_07437_),
    .B(_07438_),
    .C(_07439_),
    .X(_07440_));
 sky130_fd_sc_hd__a21oi_1 _14957_ (.A1(_07437_),
    .A2(_07439_),
    .B1(_07438_),
    .Y(_07441_));
 sky130_fd_sc_hd__nor2_1 _14958_ (.A(_07440_),
    .B(_07441_),
    .Y(_07442_));
 sky130_fd_sc_hd__xor2_2 _14959_ (.A(_07433_),
    .B(_07442_),
    .X(_07443_));
 sky130_fd_sc_hd__nor3_4 _14960_ (.A(_07431_),
    .B(_07432_),
    .C(_07443_),
    .Y(_07444_));
 sky130_fd_sc_hd__o21a_1 _14961_ (.A1(_07431_),
    .A2(_07432_),
    .B1(_07443_),
    .X(_07445_));
 sky130_fd_sc_hd__a211oi_4 _14962_ (.A1(_07361_),
    .A2(_07418_),
    .B1(_07444_),
    .C1(_07445_),
    .Y(_07446_));
 sky130_fd_sc_hd__o211a_1 _14963_ (.A1(_07444_),
    .A2(_07445_),
    .B1(_07361_),
    .C1(_07418_),
    .X(_07447_));
 sky130_fd_sc_hd__nand3_1 _14964_ (.A(_06648_),
    .B(_07382_),
    .C(_07383_),
    .Y(_07448_));
 sky130_fd_sc_hd__a32o_1 _14965_ (.A1(_07367_),
    .A2(_07364_),
    .A3(_07368_),
    .B1(_07370_),
    .B2(_07363_),
    .X(_07449_));
 sky130_fd_sc_hd__and4_1 _14966_ (.A(_06929_),
    .B(_06930_),
    .C(_06440_),
    .D(_06442_),
    .X(_07450_));
 sky130_fd_sc_hd__a22o_1 _14967_ (.A1(_06930_),
    .A2(_06440_),
    .B1(_06442_),
    .B2(_06929_),
    .X(_07451_));
 sky130_fd_sc_hd__and2b_1 _14968_ (.A_N(_07450_),
    .B(_07451_),
    .X(_07452_));
 sky130_fd_sc_hd__nand2_1 _14969_ (.A(_06551_),
    .B(_06453_),
    .Y(_07453_));
 sky130_fd_sc_hd__xnor2_1 _14970_ (.A(_07452_),
    .B(_07453_),
    .Y(_07454_));
 sky130_fd_sc_hd__nand2_1 _14971_ (.A(_07377_),
    .B(_07379_),
    .Y(_07455_));
 sky130_fd_sc_hd__xor2_1 _14972_ (.A(_07454_),
    .B(_07455_),
    .X(_07456_));
 sky130_fd_sc_hd__xnor2_1 _14973_ (.A(_06543_),
    .B(_07456_),
    .Y(_07457_));
 sky130_fd_sc_hd__xnor2_1 _14974_ (.A(_07449_),
    .B(_07457_),
    .Y(_07458_));
 sky130_fd_sc_hd__a21oi_2 _14975_ (.A1(_07382_),
    .A2(_07448_),
    .B1(_07458_),
    .Y(_07459_));
 sky130_fd_sc_hd__and3_1 _14976_ (.A(_07382_),
    .B(_07448_),
    .C(_07458_),
    .X(_07460_));
 sky130_fd_sc_hd__nor4_4 _14977_ (.A(_07446_),
    .B(_07447_),
    .C(_07459_),
    .D(_07460_),
    .Y(_07461_));
 sky130_fd_sc_hd__o22a_1 _14978_ (.A1(_07446_),
    .A2(_07447_),
    .B1(_07459_),
    .B2(_07460_),
    .X(_07462_));
 sky130_fd_sc_hd__a211o_1 _14979_ (.A1(_07416_),
    .A2(_07417_),
    .B1(_07461_),
    .C1(_07462_),
    .X(_07463_));
 sky130_fd_sc_hd__o211ai_2 _14980_ (.A1(_07461_),
    .A2(_07462_),
    .B1(_07416_),
    .C1(_07417_),
    .Y(_07464_));
 sky130_fd_sc_hd__a21boi_2 _14981_ (.A1(_07376_),
    .A2(_07388_),
    .B1_N(_07387_),
    .Y(_07465_));
 sky130_fd_sc_hd__xnor2_1 _14982_ (.A(_06606_),
    .B(_07465_),
    .Y(_07466_));
 sky130_fd_sc_hd__xor2_1 _14983_ (.A(_06601_),
    .B(_07466_),
    .X(_07467_));
 sky130_fd_sc_hd__and3_1 _14984_ (.A(_07463_),
    .B(_07464_),
    .C(_07467_),
    .X(_07468_));
 sky130_fd_sc_hd__a21oi_1 _14985_ (.A1(_07463_),
    .A2(_07464_),
    .B1(_07467_),
    .Y(_07469_));
 sky130_fd_sc_hd__a211oi_2 _14986_ (.A1(_07393_),
    .A2(_07415_),
    .B1(_07468_),
    .C1(_07469_),
    .Y(_07470_));
 sky130_fd_sc_hd__o211a_1 _14987_ (.A1(_07468_),
    .A2(_07469_),
    .B1(_07393_),
    .C1(_07415_),
    .X(_07471_));
 sky130_fd_sc_hd__a211oi_2 _14988_ (.A1(_07413_),
    .A2(_07414_),
    .B1(_07470_),
    .C1(_07471_),
    .Y(_07472_));
 sky130_fd_sc_hd__o211a_1 _14989_ (.A1(_07470_),
    .A2(_07471_),
    .B1(_07413_),
    .C1(_07414_),
    .X(_07473_));
 sky130_fd_sc_hd__a211oi_1 _14990_ (.A1(_07403_),
    .A2(_07412_),
    .B1(_07472_),
    .C1(_07473_),
    .Y(_07474_));
 sky130_fd_sc_hd__o211ai_1 _14991_ (.A1(_07472_),
    .A2(_07473_),
    .B1(_07403_),
    .C1(_07412_),
    .Y(_07475_));
 sky130_fd_sc_hd__and2b_1 _14992_ (.A_N(_07474_),
    .B(_07475_),
    .X(_07476_));
 sky130_fd_sc_hd__nand2_1 _14993_ (.A(_07411_),
    .B(_07476_),
    .Y(_07477_));
 sky130_fd_sc_hd__nor2_1 _14994_ (.A(_07409_),
    .B(_07410_),
    .Y(_07478_));
 sky130_fd_sc_hd__nand2_1 _14995_ (.A(_07475_),
    .B(_07478_),
    .Y(_07479_));
 sky130_fd_sc_hd__inv_2 _14996_ (.A(_07474_),
    .Y(_07480_));
 sky130_fd_sc_hd__o211a_1 _14997_ (.A1(_07342_),
    .A2(_07477_),
    .B1(_07479_),
    .C1(_07480_),
    .X(_07481_));
 sky130_fd_sc_hd__and2b_1 _14998_ (.A_N(_07332_),
    .B(_07333_),
    .X(_07482_));
 sky130_fd_sc_hd__nor2_1 _14999_ (.A(_07482_),
    .B(_07335_),
    .Y(_07483_));
 sky130_fd_sc_hd__nand3_1 _15000_ (.A(_07291_),
    .B(_07292_),
    .C(_07295_),
    .Y(_07484_));
 sky130_fd_sc_hd__a21o_1 _15001_ (.A1(_07291_),
    .A2(_07292_),
    .B1(_07295_),
    .X(_07485_));
 sky130_fd_sc_hd__nand2_1 _15002_ (.A(_06484_),
    .B(_06896_),
    .Y(_07486_));
 sky130_fd_sc_hd__xnor2_1 _15003_ (.A(_07486_),
    .B(_07289_),
    .Y(_07487_));
 sky130_fd_sc_hd__and4_1 _15004_ (.A(\wfg_stim_sine_top.gain_val_q[9] ),
    .B(\wfg_stim_sine_top.gain_val_q[8] ),
    .C(_06970_),
    .D(\wfg_stim_sine_top.wfg_stim_sine.sin_17[1] ),
    .X(_07488_));
 sky130_fd_sc_hd__a22oi_1 _15005_ (.A1(\wfg_stim_sine_top.gain_val_q[8] ),
    .A2(_06991_),
    .B1(_06973_),
    .B2(\wfg_stim_sine_top.gain_val_q[9] ),
    .Y(_07489_));
 sky130_fd_sc_hd__and4bb_1 _15006_ (.A_N(_07488_),
    .B_N(_07489_),
    .C(_06484_),
    .D(_06982_),
    .X(_07490_));
 sky130_fd_sc_hd__nor2_1 _15007_ (.A(_07488_),
    .B(_07490_),
    .Y(_07491_));
 sky130_fd_sc_hd__xnor2_1 _15008_ (.A(_07487_),
    .B(_07491_),
    .Y(_07492_));
 sky130_fd_sc_hd__buf_6 _15009_ (.A(_06974_),
    .X(_07493_));
 sky130_fd_sc_hd__a22oi_1 _15010_ (.A1(_06450_),
    .A2(_07493_),
    .B1(_06989_),
    .B2(_06439_),
    .Y(_07494_));
 sky130_fd_sc_hd__nor2_1 _15011_ (.A(_07284_),
    .B(_07494_),
    .Y(_07495_));
 sky130_fd_sc_hd__and2_1 _15012_ (.A(_07492_),
    .B(_07495_),
    .X(_07496_));
 sky130_fd_sc_hd__nand3_4 _15013_ (.A(_07484_),
    .B(_07485_),
    .C(_07496_),
    .Y(_07497_));
 sky130_fd_sc_hd__and2b_1 _15014_ (.A_N(_07491_),
    .B(_07487_),
    .X(_07498_));
 sky130_fd_sc_hd__a21o_1 _15015_ (.A1(_07304_),
    .A2(_07305_),
    .B1(_07310_),
    .X(_07499_));
 sky130_fd_sc_hd__nand3_1 _15016_ (.A(_07311_),
    .B(_07498_),
    .C(_07499_),
    .Y(_07500_));
 sky130_fd_sc_hd__a21o_1 _15017_ (.A1(_07311_),
    .A2(_07499_),
    .B1(_07498_),
    .X(_07501_));
 sky130_fd_sc_hd__or3_1 _15018_ (.A(_07302_),
    .B(_07300_),
    .C(_07301_),
    .X(_07502_));
 sky130_fd_sc_hd__o21ai_1 _15019_ (.A1(_07302_),
    .A2(_07301_),
    .B1(_07300_),
    .Y(_07503_));
 sky130_fd_sc_hd__nand2_1 _15020_ (.A(\wfg_stim_sine_top.gain_val_q[4] ),
    .B(_06738_),
    .Y(_07504_));
 sky130_fd_sc_hd__a22oi_2 _15021_ (.A1(\wfg_stim_sine_top.gain_val_q[5] ),
    .A2(_06750_),
    .B1(_06965_),
    .B2(\wfg_stim_sine_top.gain_val_q[6] ),
    .Y(_07505_));
 sky130_fd_sc_hd__and4_1 _15022_ (.A(\wfg_stim_sine_top.gain_val_q[6] ),
    .B(\wfg_stim_sine_top.gain_val_q[5] ),
    .C(_06750_),
    .D(_06895_),
    .X(_07506_));
 sky130_fd_sc_hd__o21bai_1 _15023_ (.A1(_07504_),
    .A2(_07505_),
    .B1_N(_07506_),
    .Y(_07507_));
 sky130_fd_sc_hd__nand3_1 _15024_ (.A(_07502_),
    .B(_07503_),
    .C(_07507_),
    .Y(_07508_));
 sky130_fd_sc_hd__a21o_1 _15025_ (.A1(_07502_),
    .A2(_07503_),
    .B1(_07507_),
    .X(_07509_));
 sky130_fd_sc_hd__nand2_1 _15026_ (.A(\wfg_stim_sine_top.gain_val_q[2] ),
    .B(_06428_),
    .Y(_07510_));
 sky130_fd_sc_hd__nand2_1 _15027_ (.A(_06413_),
    .B(_06415_),
    .Y(_07511_));
 sky130_fd_sc_hd__a22o_1 _15028_ (.A1(_06539_),
    .A2(\wfg_stim_sine_top.wfg_stim_sine.sin_17[11] ),
    .B1(_06415_),
    .B2(_06538_),
    .X(_07512_));
 sky130_fd_sc_hd__o21ai_1 _15029_ (.A1(_07041_),
    .A2(_07511_),
    .B1(_07512_),
    .Y(_07513_));
 sky130_fd_sc_hd__xor2_1 _15030_ (.A(_07510_),
    .B(_07513_),
    .X(_07514_));
 sky130_fd_sc_hd__nand3_1 _15031_ (.A(_07508_),
    .B(_07509_),
    .C(_07514_),
    .Y(_07515_));
 sky130_fd_sc_hd__nand2_1 _15032_ (.A(_07508_),
    .B(_07515_),
    .Y(_07516_));
 sky130_fd_sc_hd__nand3_2 _15033_ (.A(_07500_),
    .B(_07501_),
    .C(_07516_),
    .Y(_07517_));
 sky130_fd_sc_hd__a21o_1 _15034_ (.A1(_07500_),
    .A2(_07501_),
    .B1(_07516_),
    .X(_07518_));
 sky130_fd_sc_hd__a21o_1 _15035_ (.A1(_07484_),
    .A2(_07485_),
    .B1(_07496_),
    .X(_07519_));
 sky130_fd_sc_hd__nand4_4 _15036_ (.A(_07497_),
    .B(_07517_),
    .C(_07518_),
    .D(_07519_),
    .Y(_07520_));
 sky130_fd_sc_hd__o22a_1 _15037_ (.A1(_07316_),
    .A2(_07317_),
    .B1(_07318_),
    .B2(_07297_),
    .X(_07521_));
 sky130_fd_sc_hd__a211oi_4 _15038_ (.A1(_07497_),
    .A2(_07520_),
    .B1(_07319_),
    .C1(_07521_),
    .Y(_07522_));
 sky130_fd_sc_hd__a21bo_1 _15039_ (.A1(_07501_),
    .A2(_07516_),
    .B1_N(_07500_),
    .X(_07523_));
 sky130_fd_sc_hd__o22a_1 _15040_ (.A1(_07324_),
    .A2(_07307_),
    .B1(_07309_),
    .B2(_07306_),
    .X(_07524_));
 sky130_fd_sc_hd__xnor2_1 _15041_ (.A(_07523_),
    .B(_07524_),
    .Y(_07525_));
 sky130_fd_sc_hd__nand2_1 _15042_ (.A(_06599_),
    .B(_06770_),
    .Y(_07526_));
 sky130_fd_sc_hd__xor2_1 _15043_ (.A(_07525_),
    .B(_07526_),
    .X(_07527_));
 sky130_fd_sc_hd__o211a_1 _15044_ (.A1(_07319_),
    .A2(_07521_),
    .B1(_07497_),
    .C1(_07520_),
    .X(_07528_));
 sky130_fd_sc_hd__nor3_1 _15045_ (.A(_07522_),
    .B(_07527_),
    .C(_07528_),
    .Y(_07529_));
 sky130_fd_sc_hd__or3_1 _15046_ (.A(_07321_),
    .B(_07322_),
    .C(_07328_),
    .X(_07530_));
 sky130_fd_sc_hd__o21ai_1 _15047_ (.A1(_07321_),
    .A2(_07322_),
    .B1(_07328_),
    .Y(_07531_));
 sky130_fd_sc_hd__o211a_1 _15048_ (.A1(_07522_),
    .A2(_07529_),
    .B1(_07530_),
    .C1(_07531_),
    .X(_07532_));
 sky130_fd_sc_hd__a21o_1 _15049_ (.A1(_07500_),
    .A2(_07517_),
    .B1(_07524_),
    .X(_07533_));
 sky130_fd_sc_hd__nand3_1 _15050_ (.A(_07206_),
    .B(_06770_),
    .C(_07525_),
    .Y(_07534_));
 sky130_fd_sc_hd__a211oi_1 _15051_ (.A1(_07530_),
    .A2(_07531_),
    .B1(_07522_),
    .C1(_07529_),
    .Y(_07535_));
 sky130_fd_sc_hd__a211oi_2 _15052_ (.A1(_07533_),
    .A2(_07534_),
    .B1(_07532_),
    .C1(_07535_),
    .Y(_07536_));
 sky130_fd_sc_hd__nor2_1 _15053_ (.A(_07532_),
    .B(_07536_),
    .Y(_07537_));
 sky130_fd_sc_hd__nor3_1 _15054_ (.A(_07336_),
    .B(_07483_),
    .C(_07537_),
    .Y(_07538_));
 sky130_fd_sc_hd__inv_2 _15055_ (.A(_07538_),
    .Y(_07539_));
 sky130_fd_sc_hd__xnor2_1 _15056_ (.A(_07492_),
    .B(_07495_),
    .Y(_07540_));
 sky130_fd_sc_hd__nand2_1 _15057_ (.A(_06468_),
    .B(_06989_),
    .Y(_07541_));
 sky130_fd_sc_hd__o2bb2a_1 _15058_ (.A1_N(_06484_),
    .A2_N(_06996_),
    .B1(_07488_),
    .B2(_07489_),
    .X(_07542_));
 sky130_fd_sc_hd__nor2_1 _15059_ (.A(_07490_),
    .B(_07542_),
    .Y(_07543_));
 sky130_fd_sc_hd__and4_1 _15060_ (.A(\wfg_stim_sine_top.gain_val_q[9] ),
    .B(\wfg_stim_sine_top.gain_val_q[8] ),
    .C(\wfg_stim_sine_top.wfg_stim_sine.sin_17[1] ),
    .D(\wfg_stim_sine_top.wfg_stim_sine.sin_17[0] ),
    .X(_07544_));
 sky130_fd_sc_hd__a22oi_1 _15061_ (.A1(_06488_),
    .A2(_06973_),
    .B1(_06975_),
    .B2(_06713_),
    .Y(_07545_));
 sky130_fd_sc_hd__and4bb_1 _15062_ (.A_N(_07544_),
    .B_N(_07545_),
    .C(_06484_),
    .D(_06971_),
    .X(_07546_));
 sky130_fd_sc_hd__nor2_1 _15063_ (.A(_07544_),
    .B(_07546_),
    .Y(_07547_));
 sky130_fd_sc_hd__xnor2_1 _15064_ (.A(_07543_),
    .B(_07547_),
    .Y(_07548_));
 sky130_fd_sc_hd__or2b_1 _15065_ (.A(_07541_),
    .B_N(_07548_),
    .X(_07549_));
 sky130_fd_sc_hd__nor2_1 _15066_ (.A(_07540_),
    .B(_07549_),
    .Y(_07550_));
 sky130_fd_sc_hd__xor2_1 _15067_ (.A(_07540_),
    .B(_07549_),
    .X(_07551_));
 sky130_fd_sc_hd__and2b_1 _15068_ (.A_N(_07547_),
    .B(_07543_),
    .X(_07552_));
 sky130_fd_sc_hd__a21o_1 _15069_ (.A1(_07508_),
    .A2(_07509_),
    .B1(_07514_),
    .X(_07553_));
 sky130_fd_sc_hd__nand3_1 _15070_ (.A(_07515_),
    .B(_07552_),
    .C(_07553_),
    .Y(_07554_));
 sky130_fd_sc_hd__a21o_1 _15071_ (.A1(_07515_),
    .A2(_07553_),
    .B1(_07552_),
    .X(_07555_));
 sky130_fd_sc_hd__or3_1 _15072_ (.A(_07506_),
    .B(_07504_),
    .C(_07505_),
    .X(_07556_));
 sky130_fd_sc_hd__o21ai_1 _15073_ (.A1(_07506_),
    .A2(_07505_),
    .B1(_07504_),
    .Y(_07557_));
 sky130_fd_sc_hd__nand2_1 _15074_ (.A(\wfg_stim_sine_top.gain_val_q[4] ),
    .B(_06894_),
    .Y(_07558_));
 sky130_fd_sc_hd__a22oi_2 _15075_ (.A1(_06548_),
    .A2(_06965_),
    .B1(_06982_),
    .B2(_06546_),
    .Y(_07559_));
 sky130_fd_sc_hd__and4_1 _15076_ (.A(_06546_),
    .B(\wfg_stim_sine_top.gain_val_q[5] ),
    .C(_06965_),
    .D(_06995_),
    .X(_07560_));
 sky130_fd_sc_hd__o21bai_1 _15077_ (.A1(_07558_),
    .A2(_07559_),
    .B1_N(_07560_),
    .Y(_07561_));
 sky130_fd_sc_hd__nand3_1 _15078_ (.A(_07556_),
    .B(_07557_),
    .C(_07561_),
    .Y(_07562_));
 sky130_fd_sc_hd__a21o_1 _15079_ (.A1(_07556_),
    .A2(_07557_),
    .B1(_07561_),
    .X(_07563_));
 sky130_fd_sc_hd__nand2_1 _15080_ (.A(\wfg_stim_sine_top.gain_val_q[2] ),
    .B(_06745_),
    .Y(_07564_));
 sky130_fd_sc_hd__and2_2 _15081_ (.A(_06538_),
    .B(_06539_),
    .X(_07565_));
 sky130_fd_sc_hd__and2_2 _15082_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[10] ),
    .B(_06426_),
    .X(_07566_));
 sky130_fd_sc_hd__a22o_1 _15083_ (.A1(\wfg_stim_sine_top.gain_val_q[0] ),
    .A2(\wfg_stim_sine_top.wfg_stim_sine.sin_17[10] ),
    .B1(_06427_),
    .B2(\wfg_stim_sine_top.gain_val_q[1] ),
    .X(_07567_));
 sky130_fd_sc_hd__a21bo_1 _15084_ (.A1(_07565_),
    .A2(_07566_),
    .B1_N(_07567_),
    .X(_07568_));
 sky130_fd_sc_hd__xor2_1 _15085_ (.A(_07564_),
    .B(_07568_),
    .X(_07569_));
 sky130_fd_sc_hd__nand3_1 _15086_ (.A(_07562_),
    .B(_07563_),
    .C(_07569_),
    .Y(_07570_));
 sky130_fd_sc_hd__nand2_1 _15087_ (.A(_07562_),
    .B(_07570_),
    .Y(_07571_));
 sky130_fd_sc_hd__nand3_1 _15088_ (.A(_07554_),
    .B(_07555_),
    .C(_07571_),
    .Y(_07572_));
 sky130_fd_sc_hd__a21o_1 _15089_ (.A1(_07554_),
    .A2(_07555_),
    .B1(_07571_),
    .X(_07573_));
 sky130_fd_sc_hd__and3_1 _15090_ (.A(_07551_),
    .B(_07572_),
    .C(_07573_),
    .X(_07574_));
 sky130_fd_sc_hd__a22o_1 _15091_ (.A1(_07517_),
    .A2(_07518_),
    .B1(_07519_),
    .B2(_07497_),
    .X(_07575_));
 sky130_fd_sc_hd__o211a_2 _15092_ (.A1(_07550_),
    .A2(_07574_),
    .B1(_07520_),
    .C1(_07575_),
    .X(_07576_));
 sky130_fd_sc_hd__a21bo_1 _15093_ (.A1(_07555_),
    .A2(_07571_),
    .B1_N(_07554_),
    .X(_07577_));
 sky130_fd_sc_hd__o22a_1 _15094_ (.A1(_07324_),
    .A2(_07511_),
    .B1(_07513_),
    .B2(_07510_),
    .X(_07578_));
 sky130_fd_sc_hd__xnor2_1 _15095_ (.A(_07577_),
    .B(_07578_),
    .Y(_07579_));
 sky130_fd_sc_hd__nand2_1 _15096_ (.A(_06599_),
    .B(_06430_),
    .Y(_07580_));
 sky130_fd_sc_hd__xor2_1 _15097_ (.A(_07579_),
    .B(_07580_),
    .X(_07581_));
 sky130_fd_sc_hd__a211oi_2 _15098_ (.A1(_07520_),
    .A2(_07575_),
    .B1(_07550_),
    .C1(_07574_),
    .Y(_07582_));
 sky130_fd_sc_hd__nor3_2 _15099_ (.A(_07576_),
    .B(_07581_),
    .C(_07582_),
    .Y(_07583_));
 sky130_fd_sc_hd__or3_1 _15100_ (.A(_07522_),
    .B(_07527_),
    .C(_07528_),
    .X(_07584_));
 sky130_fd_sc_hd__o21ai_2 _15101_ (.A1(_07522_),
    .A2(_07528_),
    .B1(_07527_),
    .Y(_07585_));
 sky130_fd_sc_hd__o211ai_4 _15102_ (.A1(_07576_),
    .A2(_07583_),
    .B1(_07584_),
    .C1(_07585_),
    .Y(_07586_));
 sky130_fd_sc_hd__a21oi_1 _15103_ (.A1(_07554_),
    .A2(_07572_),
    .B1(_07578_),
    .Y(_07587_));
 sky130_fd_sc_hd__and3_1 _15104_ (.A(_07200_),
    .B(_06430_),
    .C(_07579_),
    .X(_07588_));
 sky130_fd_sc_hd__a211o_1 _15105_ (.A1(_07584_),
    .A2(_07585_),
    .B1(_07576_),
    .C1(_07583_),
    .X(_07589_));
 sky130_fd_sc_hd__o211ai_2 _15106_ (.A1(_07587_),
    .A2(_07588_),
    .B1(_07586_),
    .C1(_07589_),
    .Y(_07590_));
 sky130_fd_sc_hd__o211a_1 _15107_ (.A1(_07532_),
    .A2(_07535_),
    .B1(_07533_),
    .C1(_07534_),
    .X(_07591_));
 sky130_fd_sc_hd__a211oi_1 _15108_ (.A1(_07586_),
    .A2(_07590_),
    .B1(_07536_),
    .C1(_07591_),
    .Y(_07592_));
 sky130_fd_sc_hd__inv_2 _15109_ (.A(_07592_),
    .Y(_07593_));
 sky130_fd_sc_hd__or3_1 _15110_ (.A(_07560_),
    .B(_07558_),
    .C(_07559_),
    .X(_07594_));
 sky130_fd_sc_hd__o21ai_1 _15111_ (.A1(_07560_),
    .A2(_07559_),
    .B1(_07558_),
    .Y(_07595_));
 sky130_fd_sc_hd__and2_1 _15112_ (.A(\wfg_stim_sine_top.gain_val_q[4] ),
    .B(_06965_),
    .X(_07596_));
 sky130_fd_sc_hd__a22o_1 _15113_ (.A1(_06548_),
    .A2(_06995_),
    .B1(_06991_),
    .B2(_06546_),
    .X(_07597_));
 sky130_fd_sc_hd__nand4_1 _15114_ (.A(_06546_),
    .B(_06548_),
    .C(_06982_),
    .D(_06991_),
    .Y(_07598_));
 sky130_fd_sc_hd__a21bo_1 _15115_ (.A1(_07596_),
    .A2(_07597_),
    .B1_N(_07598_),
    .X(_07599_));
 sky130_fd_sc_hd__nand3_1 _15116_ (.A(_07594_),
    .B(_07595_),
    .C(_07599_),
    .Y(_07600_));
 sky130_fd_sc_hd__and2_2 _15117_ (.A(_06426_),
    .B(_06744_),
    .X(_07601_));
 sky130_fd_sc_hd__a22o_1 _15118_ (.A1(_06539_),
    .A2(_06427_),
    .B1(_06747_),
    .B2(_06538_),
    .X(_07602_));
 sky130_fd_sc_hd__a21bo_1 _15119_ (.A1(_07565_),
    .A2(_07601_),
    .B1_N(_07602_),
    .X(_07603_));
 sky130_fd_sc_hd__nand2_1 _15120_ (.A(\wfg_stim_sine_top.gain_val_q[2] ),
    .B(_06754_),
    .Y(_07604_));
 sky130_fd_sc_hd__xor2_1 _15121_ (.A(_07603_),
    .B(_07604_),
    .X(_07605_));
 sky130_fd_sc_hd__a21o_1 _15122_ (.A1(_07594_),
    .A2(_07595_),
    .B1(_07599_),
    .X(_07606_));
 sky130_fd_sc_hd__nand3_1 _15123_ (.A(_07600_),
    .B(_07605_),
    .C(_07606_),
    .Y(_07607_));
 sky130_fd_sc_hd__a21o_1 _15124_ (.A1(_07600_),
    .A2(_07606_),
    .B1(_07605_),
    .X(_07608_));
 sky130_fd_sc_hd__nand2_1 _15125_ (.A(_06744_),
    .B(_06736_),
    .Y(_07609_));
 sky130_fd_sc_hd__a22o_1 _15126_ (.A1(_06539_),
    .A2(_06747_),
    .B1(_06737_),
    .B2(_06538_),
    .X(_07610_));
 sky130_fd_sc_hd__o21ai_1 _15127_ (.A1(_07041_),
    .A2(_07609_),
    .B1(_07610_),
    .Y(_07611_));
 sky130_fd_sc_hd__nand2_1 _15128_ (.A(\wfg_stim_sine_top.gain_val_q[2] ),
    .B(_06742_),
    .Y(_07612_));
 sky130_fd_sc_hd__xor2_1 _15129_ (.A(_07611_),
    .B(_07612_),
    .X(_07613_));
 sky130_fd_sc_hd__nand3_1 _15130_ (.A(_07598_),
    .B(_07596_),
    .C(_07597_),
    .Y(_07614_));
 sky130_fd_sc_hd__a22o_1 _15131_ (.A1(_06544_),
    .A2(_06896_),
    .B1(_07598_),
    .B2(_07597_),
    .X(_07615_));
 sky130_fd_sc_hd__nand2_1 _15132_ (.A(\wfg_stim_sine_top.gain_val_q[4] ),
    .B(_06995_),
    .Y(_07616_));
 sky130_fd_sc_hd__a22oi_2 _15133_ (.A1(\wfg_stim_sine_top.gain_val_q[5] ),
    .A2(_06991_),
    .B1(_06973_),
    .B2(_06546_),
    .Y(_07617_));
 sky130_fd_sc_hd__and4_1 _15134_ (.A(\wfg_stim_sine_top.gain_val_q[6] ),
    .B(\wfg_stim_sine_top.gain_val_q[5] ),
    .C(_06970_),
    .D(\wfg_stim_sine_top.wfg_stim_sine.sin_17[1] ),
    .X(_07618_));
 sky130_fd_sc_hd__o21bai_1 _15135_ (.A1(_07616_),
    .A2(_07617_),
    .B1_N(_07618_),
    .Y(_07619_));
 sky130_fd_sc_hd__a21o_1 _15136_ (.A1(_07614_),
    .A2(_07615_),
    .B1(_07619_),
    .X(_07620_));
 sky130_fd_sc_hd__nand3_1 _15137_ (.A(_07614_),
    .B(_07615_),
    .C(_07619_),
    .Y(_07621_));
 sky130_fd_sc_hd__a21bo_1 _15138_ (.A1(_07613_),
    .A2(_07620_),
    .B1_N(_07621_),
    .X(_07622_));
 sky130_fd_sc_hd__and3_1 _15139_ (.A(_07607_),
    .B(_07608_),
    .C(_07622_),
    .X(_07623_));
 sky130_fd_sc_hd__a32o_1 _15140_ (.A1(_06605_),
    .A2(_06754_),
    .A3(_07602_),
    .B1(_07601_),
    .B2(_07565_),
    .X(_07624_));
 sky130_fd_sc_hd__and2_1 _15141_ (.A(_07623_),
    .B(_07624_),
    .X(_07625_));
 sky130_fd_sc_hd__nor2_1 _15142_ (.A(_07623_),
    .B(_07624_),
    .Y(_07626_));
 sky130_fd_sc_hd__nor2_1 _15143_ (.A(_07625_),
    .B(_07626_),
    .Y(_07627_));
 sky130_fd_sc_hd__a31o_1 _15144_ (.A1(_07206_),
    .A2(_06754_),
    .A3(_07627_),
    .B1(_07625_),
    .X(_07628_));
 sky130_fd_sc_hd__o2bb2a_1 _15145_ (.A1_N(_06484_),
    .A2_N(_06971_),
    .B1(_07544_),
    .B2(_07545_),
    .X(_07629_));
 sky130_fd_sc_hd__nor2_1 _15146_ (.A(_07546_),
    .B(_07629_),
    .Y(_07630_));
 sky130_fd_sc_hd__and4_1 _15147_ (.A(_06725_),
    .B(_06485_),
    .C(_07493_),
    .D(_06989_),
    .X(_07631_));
 sky130_fd_sc_hd__and2_1 _15148_ (.A(_07630_),
    .B(_07631_),
    .X(_07632_));
 sky130_fd_sc_hd__a21o_1 _15149_ (.A1(_07562_),
    .A2(_07563_),
    .B1(_07569_),
    .X(_07633_));
 sky130_fd_sc_hd__nand3_1 _15150_ (.A(_07570_),
    .B(_07632_),
    .C(_07633_),
    .Y(_07634_));
 sky130_fd_sc_hd__a21o_1 _15151_ (.A1(_07570_),
    .A2(_07633_),
    .B1(_07632_),
    .X(_07635_));
 sky130_fd_sc_hd__nand2_1 _15152_ (.A(_07600_),
    .B(_07607_),
    .Y(_07636_));
 sky130_fd_sc_hd__nand3_1 _15153_ (.A(_07634_),
    .B(_07635_),
    .C(_07636_),
    .Y(_07637_));
 sky130_fd_sc_hd__a21o_1 _15154_ (.A1(_07634_),
    .A2(_07635_),
    .B1(_07636_),
    .X(_07638_));
 sky130_fd_sc_hd__xnor2_1 _15155_ (.A(_07541_),
    .B(_07548_),
    .Y(_07639_));
 sky130_fd_sc_hd__and3_1 _15156_ (.A(_07637_),
    .B(_07638_),
    .C(_07639_),
    .X(_07640_));
 sky130_fd_sc_hd__a21oi_1 _15157_ (.A1(_07607_),
    .A2(_07608_),
    .B1(_07622_),
    .Y(_07641_));
 sky130_fd_sc_hd__nor2_1 _15158_ (.A(_07630_),
    .B(_07631_),
    .Y(_07642_));
 sky130_fd_sc_hd__or2_1 _15159_ (.A(_07632_),
    .B(_07642_),
    .X(_07643_));
 sky130_fd_sc_hd__or3_2 _15160_ (.A(_07623_),
    .B(_07641_),
    .C(_07643_),
    .X(_07644_));
 sky130_fd_sc_hd__a21oi_1 _15161_ (.A1(_07637_),
    .A2(_07638_),
    .B1(_07639_),
    .Y(_07645_));
 sky130_fd_sc_hd__or3_2 _15162_ (.A(_07640_),
    .B(_07644_),
    .C(_07645_),
    .X(_07646_));
 sky130_fd_sc_hd__nand2_1 _15163_ (.A(_06599_),
    .B(_06754_),
    .Y(_07647_));
 sky130_fd_sc_hd__xnor2_1 _15164_ (.A(_07627_),
    .B(_07647_),
    .Y(_07648_));
 sky130_fd_sc_hd__o21ai_1 _15165_ (.A1(_07640_),
    .A2(_07645_),
    .B1(_07644_),
    .Y(_07649_));
 sky130_fd_sc_hd__nand3_2 _15166_ (.A(_07646_),
    .B(_07648_),
    .C(_07649_),
    .Y(_07650_));
 sky130_fd_sc_hd__a21oi_1 _15167_ (.A1(_07572_),
    .A2(_07573_),
    .B1(_07551_),
    .Y(_07651_));
 sky130_fd_sc_hd__or3b_1 _15168_ (.A(_07574_),
    .B(_07651_),
    .C_N(_07640_),
    .X(_07652_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15169_ (.A(_07652_),
    .X(_07653_));
 sky130_fd_sc_hd__a21bo_1 _15170_ (.A1(_07635_),
    .A2(_07636_),
    .B1_N(_07634_),
    .X(_07654_));
 sky130_fd_sc_hd__o2bb2a_1 _15171_ (.A1_N(_07565_),
    .A2_N(_07566_),
    .B1(_07568_),
    .B2(_07564_),
    .X(_07655_));
 sky130_fd_sc_hd__xnor2_1 _15172_ (.A(_07654_),
    .B(_07655_),
    .Y(_07656_));
 sky130_fd_sc_hd__nand2_1 _15173_ (.A(_06599_),
    .B(_06748_),
    .Y(_07657_));
 sky130_fd_sc_hd__xnor2_1 _15174_ (.A(_07656_),
    .B(_07657_),
    .Y(_07658_));
 sky130_fd_sc_hd__o21bai_1 _15175_ (.A1(_07574_),
    .A2(_07651_),
    .B1_N(_07640_),
    .Y(_07659_));
 sky130_fd_sc_hd__and3_1 _15176_ (.A(_07653_),
    .B(_07658_),
    .C(_07659_),
    .X(_07660_));
 sky130_fd_sc_hd__a21oi_1 _15177_ (.A1(_07653_),
    .A2(_07659_),
    .B1(_07658_),
    .Y(_07661_));
 sky130_fd_sc_hd__a211oi_1 _15178_ (.A1(_07646_),
    .A2(_07650_),
    .B1(_07660_),
    .C1(_07661_),
    .Y(_07662_));
 sky130_fd_sc_hd__o211a_1 _15179_ (.A1(_07660_),
    .A2(_07661_),
    .B1(_07646_),
    .C1(_07650_),
    .X(_07663_));
 sky130_fd_sc_hd__nor2_1 _15180_ (.A(_07662_),
    .B(_07663_),
    .Y(_07664_));
 sky130_fd_sc_hd__xor2_1 _15181_ (.A(_07628_),
    .B(_07664_),
    .X(_07665_));
 sky130_fd_sc_hd__nand3_1 _15182_ (.A(_07621_),
    .B(_07613_),
    .C(_07620_),
    .Y(_07666_));
 sky130_fd_sc_hd__a21o_1 _15183_ (.A1(_07621_),
    .A2(_07620_),
    .B1(_07613_),
    .X(_07667_));
 sky130_fd_sc_hd__nand2_2 _15184_ (.A(_06736_),
    .B(\wfg_stim_sine_top.wfg_stim_sine.sin_17[6] ),
    .Y(_07668_));
 sky130_fd_sc_hd__a22o_1 _15185_ (.A1(_06539_),
    .A2(_06737_),
    .B1(_06738_),
    .B2(_06538_),
    .X(_07669_));
 sky130_fd_sc_hd__o21ai_1 _15186_ (.A1(_07041_),
    .A2(_07668_),
    .B1(_07669_),
    .Y(_07670_));
 sky130_fd_sc_hd__nand2_1 _15187_ (.A(\wfg_stim_sine_top.gain_val_q[2] ),
    .B(_06752_),
    .Y(_07671_));
 sky130_fd_sc_hd__xor2_1 _15188_ (.A(_07670_),
    .B(_07671_),
    .X(_07672_));
 sky130_fd_sc_hd__or3_1 _15189_ (.A(_07618_),
    .B(_07616_),
    .C(_07617_),
    .X(_07673_));
 sky130_fd_sc_hd__o21ai_1 _15190_ (.A1(_07618_),
    .A2(_07617_),
    .B1(_07616_),
    .Y(_07674_));
 sky130_fd_sc_hd__and2_1 _15191_ (.A(\wfg_stim_sine_top.gain_val_q[4] ),
    .B(_06991_),
    .X(_07675_));
 sky130_fd_sc_hd__a22o_1 _15192_ (.A1(_06548_),
    .A2(_06973_),
    .B1(_06975_),
    .B2(_06546_),
    .X(_07676_));
 sky130_fd_sc_hd__nand4_1 _15193_ (.A(_06929_),
    .B(_06548_),
    .C(_06973_),
    .D(_06975_),
    .Y(_07677_));
 sky130_fd_sc_hd__a21bo_1 _15194_ (.A1(_07675_),
    .A2(_07676_),
    .B1_N(_07677_),
    .X(_07678_));
 sky130_fd_sc_hd__a21o_1 _15195_ (.A1(_07673_),
    .A2(_07674_),
    .B1(_07678_),
    .X(_07679_));
 sky130_fd_sc_hd__nand3_1 _15196_ (.A(_07673_),
    .B(_07674_),
    .C(_07678_),
    .Y(_07680_));
 sky130_fd_sc_hd__a21bo_1 _15197_ (.A1(_07672_),
    .A2(_07679_),
    .B1_N(_07680_),
    .X(_07681_));
 sky130_fd_sc_hd__and3_1 _15198_ (.A(_07666_),
    .B(_07667_),
    .C(_07681_),
    .X(_07682_));
 sky130_fd_sc_hd__o22ai_1 _15199_ (.A1(_07324_),
    .A2(_07609_),
    .B1(_07611_),
    .B2(_07612_),
    .Y(_07683_));
 sky130_fd_sc_hd__xor2_1 _15200_ (.A(_07682_),
    .B(_07683_),
    .X(_07684_));
 sky130_fd_sc_hd__and2_1 _15201_ (.A(_07682_),
    .B(_07683_),
    .X(_07685_));
 sky130_fd_sc_hd__a31o_1 _15202_ (.A1(_07206_),
    .A2(_06742_),
    .A3(_07684_),
    .B1(_07685_),
    .X(_07686_));
 sky130_fd_sc_hd__a21o_1 _15203_ (.A1(_07646_),
    .A2(_07649_),
    .B1(_07648_),
    .X(_07687_));
 sky130_fd_sc_hd__a21oi_1 _15204_ (.A1(_07666_),
    .A2(_07667_),
    .B1(_07681_),
    .Y(_07688_));
 sky130_fd_sc_hd__buf_4 _15205_ (.A(_06989_),
    .X(_07689_));
 sky130_fd_sc_hd__a22o_1 _15206_ (.A1(_06486_),
    .A2(_07493_),
    .B1(_07689_),
    .B2(_06725_),
    .X(_07690_));
 sky130_fd_sc_hd__or4b_2 _15207_ (.A(_07631_),
    .B(_07682_),
    .C(_07688_),
    .D_N(_07690_),
    .X(_07691_));
 sky130_fd_sc_hd__o21ai_1 _15208_ (.A1(_07623_),
    .A2(_07641_),
    .B1(_07643_),
    .Y(_07692_));
 sky130_fd_sc_hd__nand3b_1 _15209_ (.A_N(_07691_),
    .B(_07692_),
    .C(_07644_),
    .Y(_07693_));
 sky130_fd_sc_hd__inv_2 _15210_ (.A(_07693_),
    .Y(_07694_));
 sky130_fd_sc_hd__nand2_1 _15211_ (.A(_06599_),
    .B(_06742_),
    .Y(_07695_));
 sky130_fd_sc_hd__xnor2_1 _15212_ (.A(_07684_),
    .B(_07695_),
    .Y(_07696_));
 sky130_fd_sc_hd__a21bo_1 _15213_ (.A1(_07644_),
    .A2(_07692_),
    .B1_N(_07691_),
    .X(_07697_));
 sky130_fd_sc_hd__and3_1 _15214_ (.A(_07693_),
    .B(_07696_),
    .C(_07697_),
    .X(_07698_));
 sky130_fd_sc_hd__a211o_1 _15215_ (.A1(_07650_),
    .A2(_07687_),
    .B1(_07694_),
    .C1(_07698_),
    .X(_07699_));
 sky130_fd_sc_hd__o211a_1 _15216_ (.A1(_07694_),
    .A2(_07698_),
    .B1(_07650_),
    .C1(_07687_),
    .X(_07700_));
 sky130_fd_sc_hd__a21o_1 _15217_ (.A1(_07686_),
    .A2(_07699_),
    .B1(_07700_),
    .X(_07701_));
 sky130_fd_sc_hd__or2b_1 _15218_ (.A(_07700_),
    .B_N(_07699_),
    .X(_07702_));
 sky130_fd_sc_hd__xnor2_2 _15219_ (.A(_07686_),
    .B(_07702_),
    .Y(_07703_));
 sky130_fd_sc_hd__nand3_1 _15220_ (.A(_07680_),
    .B(_07672_),
    .C(_07679_),
    .Y(_07704_));
 sky130_fd_sc_hd__a21o_1 _15221_ (.A1(_07680_),
    .A2(_07679_),
    .B1(_07672_),
    .X(_07705_));
 sky130_fd_sc_hd__nand3_1 _15222_ (.A(_07677_),
    .B(_07675_),
    .C(_07676_),
    .Y(_07706_));
 sky130_fd_sc_hd__a21o_1 _15223_ (.A1(_07677_),
    .A2(_07676_),
    .B1(_07675_),
    .X(_07707_));
 sky130_fd_sc_hd__and4_1 _15224_ (.A(_06549_),
    .B(_06544_),
    .C(_06974_),
    .D(_06989_),
    .X(_07708_));
 sky130_fd_sc_hd__a21o_1 _15225_ (.A1(_07706_),
    .A2(_07707_),
    .B1(_07708_),
    .X(_07709_));
 sky130_fd_sc_hd__and2_1 _15226_ (.A(\wfg_stim_sine_top.gain_val_q[2] ),
    .B(_07007_),
    .X(_07710_));
 sky130_fd_sc_hd__nand2_1 _15227_ (.A(_06738_),
    .B(\wfg_stim_sine_top.wfg_stim_sine.sin_17[5] ),
    .Y(_07711_));
 sky130_fd_sc_hd__a22o_1 _15228_ (.A1(_06539_),
    .A2(_06739_),
    .B1(_06894_),
    .B2(_06538_),
    .X(_07712_));
 sky130_fd_sc_hd__o21ai_1 _15229_ (.A1(_07041_),
    .A2(_07711_),
    .B1(_07712_),
    .Y(_07713_));
 sky130_fd_sc_hd__xnor2_1 _15230_ (.A(_07710_),
    .B(_07713_),
    .Y(_07714_));
 sky130_fd_sc_hd__nand3_1 _15231_ (.A(_07706_),
    .B(_07708_),
    .C(_07707_),
    .Y(_07715_));
 sky130_fd_sc_hd__a21bo_1 _15232_ (.A1(_07709_),
    .A2(_07714_),
    .B1_N(_07715_),
    .X(_07716_));
 sky130_fd_sc_hd__and3_1 _15233_ (.A(_07704_),
    .B(_07705_),
    .C(_07716_),
    .X(_07717_));
 sky130_fd_sc_hd__o22ai_2 _15234_ (.A1(_07324_),
    .A2(_07668_),
    .B1(_07670_),
    .B2(_07671_),
    .Y(_07718_));
 sky130_fd_sc_hd__xor2_1 _15235_ (.A(_07717_),
    .B(_07718_),
    .X(_07719_));
 sky130_fd_sc_hd__and2_1 _15236_ (.A(_07717_),
    .B(_07718_),
    .X(_07720_));
 sky130_fd_sc_hd__a31o_1 _15237_ (.A1(_07200_),
    .A2(_06752_),
    .A3(_07719_),
    .B1(_07720_),
    .X(_07721_));
 sky130_fd_sc_hd__a21oi_1 _15238_ (.A1(_07693_),
    .A2(_07697_),
    .B1(_07696_),
    .Y(_07722_));
 sky130_fd_sc_hd__or2_1 _15239_ (.A(_07698_),
    .B(_07722_),
    .X(_07723_));
 sky130_fd_sc_hd__clkinv_2 _15240_ (.A(_07631_),
    .Y(_07724_));
 sky130_fd_sc_hd__a2bb2o_1 _15241_ (.A1_N(_07682_),
    .A2_N(_07688_),
    .B1(_07690_),
    .B2(_07724_),
    .X(_07725_));
 sky130_fd_sc_hd__nand2_1 _15242_ (.A(_06486_),
    .B(_07689_),
    .Y(_07726_));
 sky130_fd_sc_hd__a21oi_1 _15243_ (.A1(_07704_),
    .A2(_07705_),
    .B1(_07716_),
    .Y(_07727_));
 sky130_fd_sc_hd__nor3_1 _15244_ (.A(_07726_),
    .B(_07717_),
    .C(_07727_),
    .Y(_07728_));
 sky130_fd_sc_hd__a21o_1 _15245_ (.A1(_07691_),
    .A2(_07725_),
    .B1(_07728_),
    .X(_07729_));
 sky130_fd_sc_hd__nand2_1 _15246_ (.A(\wfg_stim_sine_top.gain_val_q[3] ),
    .B(_06752_),
    .Y(_07730_));
 sky130_fd_sc_hd__xnor2_1 _15247_ (.A(_07730_),
    .B(_07719_),
    .Y(_07731_));
 sky130_fd_sc_hd__nand3_1 _15248_ (.A(_07691_),
    .B(_07728_),
    .C(_07725_),
    .Y(_07732_));
 sky130_fd_sc_hd__a21boi_1 _15249_ (.A1(_07729_),
    .A2(_07731_),
    .B1_N(_07732_),
    .Y(_07733_));
 sky130_fd_sc_hd__nand2_1 _15250_ (.A(_07723_),
    .B(_07733_),
    .Y(_07734_));
 sky130_fd_sc_hd__nor2_1 _15251_ (.A(_07723_),
    .B(_07733_),
    .Y(_07735_));
 sky130_fd_sc_hd__a21o_1 _15252_ (.A1(_07721_),
    .A2(_07734_),
    .B1(_07735_),
    .X(_07736_));
 sky130_fd_sc_hd__a22o_1 _15253_ (.A1(_07665_),
    .A2(_07701_),
    .B1(_07703_),
    .B2(_07736_),
    .X(_07737_));
 sky130_fd_sc_hd__and3_1 _15254_ (.A(_07732_),
    .B(_07729_),
    .C(_07731_),
    .X(_07738_));
 sky130_fd_sc_hd__nand3_1 _15255_ (.A(_07715_),
    .B(_07709_),
    .C(_07714_),
    .Y(_07739_));
 sky130_fd_sc_hd__nand2_2 _15256_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[5] ),
    .B(_06895_),
    .Y(_07740_));
 sky130_fd_sc_hd__a22o_1 _15257_ (.A1(_07043_),
    .A2(_06894_),
    .B1(_06896_),
    .B2(_07044_),
    .X(_07741_));
 sky130_fd_sc_hd__o21ai_2 _15258_ (.A1(_07041_),
    .A2(_07740_),
    .B1(_07741_),
    .Y(_07742_));
 sky130_fd_sc_hd__nand2_1 _15259_ (.A(_06604_),
    .B(_06996_),
    .Y(_07743_));
 sky130_fd_sc_hd__xnor2_1 _15260_ (.A(_07742_),
    .B(_07743_),
    .Y(_07744_));
 sky130_fd_sc_hd__a22oi_1 _15261_ (.A1(_06544_),
    .A2(_07493_),
    .B1(_06989_),
    .B2(_06549_),
    .Y(_07745_));
 sky130_fd_sc_hd__or2_1 _15262_ (.A(_07708_),
    .B(_07745_),
    .X(_07746_));
 sky130_fd_sc_hd__nor2_1 _15263_ (.A(_07744_),
    .B(_07746_),
    .Y(_07747_));
 sky130_fd_sc_hd__a21o_1 _15264_ (.A1(_07715_),
    .A2(_07709_),
    .B1(_07714_),
    .X(_07748_));
 sky130_fd_sc_hd__and3_1 _15265_ (.A(_07739_),
    .B(_07747_),
    .C(_07748_),
    .X(_07749_));
 sky130_fd_sc_hd__o2bb2a_1 _15266_ (.A1_N(_07710_),
    .A2_N(_07712_),
    .B1(_07711_),
    .B2(_07324_),
    .X(_07750_));
 sky130_fd_sc_hd__xor2_1 _15267_ (.A(_07749_),
    .B(_07750_),
    .X(_07751_));
 sky130_fd_sc_hd__nand2_1 _15268_ (.A(\wfg_stim_sine_top.gain_val_q[3] ),
    .B(_07007_),
    .Y(_07752_));
 sky130_fd_sc_hd__xor2_1 _15269_ (.A(_07751_),
    .B(_07752_),
    .X(_07753_));
 sky130_fd_sc_hd__o21a_1 _15270_ (.A1(_07717_),
    .A2(_07727_),
    .B1(_07726_),
    .X(_07754_));
 sky130_fd_sc_hd__nor2_1 _15271_ (.A(_07728_),
    .B(_07754_),
    .Y(_07755_));
 sky130_fd_sc_hd__nand2_1 _15272_ (.A(_07753_),
    .B(_07755_),
    .Y(_07756_));
 sky130_fd_sc_hd__a21oi_1 _15273_ (.A1(_07732_),
    .A2(_07729_),
    .B1(_07731_),
    .Y(_07757_));
 sky130_fd_sc_hd__or3_1 _15274_ (.A(_07738_),
    .B(_07756_),
    .C(_07757_),
    .X(_07758_));
 sky130_fd_sc_hd__or2b_1 _15275_ (.A(_07750_),
    .B_N(_07749_),
    .X(_07759_));
 sky130_fd_sc_hd__o21ai_1 _15276_ (.A1(_07751_),
    .A2(_07752_),
    .B1(_07759_),
    .Y(_07760_));
 sky130_fd_sc_hd__o21ai_1 _15277_ (.A1(_07738_),
    .A2(_07757_),
    .B1(_07756_),
    .Y(_07761_));
 sky130_fd_sc_hd__nand3_1 _15278_ (.A(_07758_),
    .B(_07760_),
    .C(_07761_),
    .Y(_07762_));
 sky130_fd_sc_hd__a21o_1 _15279_ (.A1(_07758_),
    .A2(_07761_),
    .B1(_07760_),
    .X(_07763_));
 sky130_fd_sc_hd__nand2_2 _15280_ (.A(_06895_),
    .B(\wfg_stim_sine_top.wfg_stim_sine.sin_17[3] ),
    .Y(_07764_));
 sky130_fd_sc_hd__a22o_1 _15281_ (.A1(_07043_),
    .A2(_07007_),
    .B1(_06996_),
    .B2(_07044_),
    .X(_07765_));
 sky130_fd_sc_hd__o21a_1 _15282_ (.A1(_07324_),
    .A2(_07764_),
    .B1(_07765_),
    .X(_07766_));
 sky130_fd_sc_hd__nand2_1 _15283_ (.A(_06604_),
    .B(_06972_),
    .Y(_07767_));
 sky130_fd_sc_hd__xnor2_1 _15284_ (.A(_07766_),
    .B(_07767_),
    .Y(_07768_));
 sky130_fd_sc_hd__nand3_1 _15285_ (.A(_06551_),
    .B(_07689_),
    .C(_07768_),
    .Y(_07769_));
 sky130_fd_sc_hd__xnor2_1 _15286_ (.A(_07744_),
    .B(_07746_),
    .Y(_07770_));
 sky130_fd_sc_hd__nor2_1 _15287_ (.A(_07769_),
    .B(_07770_),
    .Y(_07771_));
 sky130_fd_sc_hd__o22ai_2 _15288_ (.A1(_07324_),
    .A2(_07740_),
    .B1(_07742_),
    .B2(_07743_),
    .Y(_07772_));
 sky130_fd_sc_hd__xor2_1 _15289_ (.A(_07771_),
    .B(_07772_),
    .X(_07773_));
 sky130_fd_sc_hd__and2_1 _15290_ (.A(_07771_),
    .B(_07772_),
    .X(_07774_));
 sky130_fd_sc_hd__a31o_1 _15291_ (.A1(_07200_),
    .A2(_06996_),
    .A3(_07773_),
    .B1(_07774_),
    .X(_07775_));
 sky130_fd_sc_hd__xnor2_1 _15292_ (.A(_07753_),
    .B(_07755_),
    .Y(_07776_));
 sky130_fd_sc_hd__nand2_1 _15293_ (.A(\wfg_stim_sine_top.gain_val_q[3] ),
    .B(_06996_),
    .Y(_07777_));
 sky130_fd_sc_hd__xor2_1 _15294_ (.A(_07773_),
    .B(_07777_),
    .X(_07778_));
 sky130_fd_sc_hd__a21oi_1 _15295_ (.A1(_07739_),
    .A2(_07748_),
    .B1(_07747_),
    .Y(_07779_));
 sky130_fd_sc_hd__or3_1 _15296_ (.A(_07749_),
    .B(_07778_),
    .C(_07779_),
    .X(_07780_));
 sky130_fd_sc_hd__xor2_1 _15297_ (.A(_07776_),
    .B(_07780_),
    .X(_07781_));
 sky130_fd_sc_hd__nor2_1 _15298_ (.A(_07776_),
    .B(_07780_),
    .Y(_07782_));
 sky130_fd_sc_hd__a21o_1 _15299_ (.A1(_07775_),
    .A2(_07781_),
    .B1(_07782_),
    .X(_07783_));
 sky130_fd_sc_hd__nand2_1 _15300_ (.A(_07758_),
    .B(_07762_),
    .Y(_07784_));
 sky130_fd_sc_hd__xnor2_1 _15301_ (.A(_07723_),
    .B(_07733_),
    .Y(_07785_));
 sky130_fd_sc_hd__xnor2_1 _15302_ (.A(_07721_),
    .B(_07785_),
    .Y(_07786_));
 sky130_fd_sc_hd__a32o_1 _15303_ (.A1(_07762_),
    .A2(_07763_),
    .A3(_07783_),
    .B1(_07784_),
    .B2(_07786_),
    .X(_07787_));
 sky130_fd_sc_hd__nand2_1 _15304_ (.A(_07775_),
    .B(_07781_),
    .Y(_07788_));
 sky130_fd_sc_hd__a21o_1 _15305_ (.A1(_07762_),
    .A2(_07763_),
    .B1(_07783_),
    .X(_07789_));
 sky130_fd_sc_hd__nor2_1 _15306_ (.A(_07324_),
    .B(_07764_),
    .Y(_07790_));
 sky130_fd_sc_hd__a31o_1 _15307_ (.A1(_06605_),
    .A2(_06972_),
    .A3(_07765_),
    .B1(_07790_),
    .X(_07791_));
 sky130_fd_sc_hd__nand2_1 _15308_ (.A(_06599_),
    .B(_06972_),
    .Y(_07792_));
 sky130_fd_sc_hd__xor2_1 _15309_ (.A(_07791_),
    .B(_07792_),
    .X(_07793_));
 sky130_fd_sc_hd__and2_1 _15310_ (.A(_07769_),
    .B(_07770_),
    .X(_07794_));
 sky130_fd_sc_hd__or2_1 _15311_ (.A(_07771_),
    .B(_07794_),
    .X(_07795_));
 sky130_fd_sc_hd__nor2_1 _15312_ (.A(_07793_),
    .B(_07795_),
    .Y(_07796_));
 sky130_fd_sc_hd__and2_1 _15313_ (.A(_07793_),
    .B(_07795_),
    .X(_07797_));
 sky130_fd_sc_hd__nor2_1 _15314_ (.A(_07796_),
    .B(_07797_),
    .Y(_07798_));
 sky130_fd_sc_hd__a22o_1 _15315_ (.A1(_07043_),
    .A2(_06996_),
    .B1(_06972_),
    .B2(_07044_),
    .X(_07799_));
 sky130_fd_sc_hd__and2_2 _15316_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[3] ),
    .B(_06970_),
    .X(_07800_));
 sky130_fd_sc_hd__a32o_1 _15317_ (.A1(_06604_),
    .A2(_07493_),
    .A3(_07799_),
    .B1(_07800_),
    .B2(_07565_),
    .X(_07801_));
 sky130_fd_sc_hd__nand2_1 _15318_ (.A(\wfg_stim_sine_top.gain_val_q[3] ),
    .B(_07493_),
    .Y(_07802_));
 sky130_fd_sc_hd__xor2_1 _15319_ (.A(_07801_),
    .B(_07802_),
    .X(_07803_));
 sky130_fd_sc_hd__a21o_1 _15320_ (.A1(_06551_),
    .A2(_07689_),
    .B1(_07768_),
    .X(_07804_));
 sky130_fd_sc_hd__nand2_1 _15321_ (.A(_07769_),
    .B(_07804_),
    .Y(_07805_));
 sky130_fd_sc_hd__nor2_1 _15322_ (.A(_07803_),
    .B(_07805_),
    .Y(_07806_));
 sky130_fd_sc_hd__a31o_1 _15323_ (.A1(_07200_),
    .A2(_07493_),
    .A3(_07801_),
    .B1(_07806_),
    .X(_07807_));
 sky130_fd_sc_hd__nor2_1 _15324_ (.A(_07749_),
    .B(_07779_),
    .Y(_07808_));
 sky130_fd_sc_hd__xnor2_1 _15325_ (.A(_07778_),
    .B(_07808_),
    .Y(_07809_));
 sky130_fd_sc_hd__a31o_1 _15326_ (.A1(_07200_),
    .A2(_06972_),
    .A3(_07791_),
    .B1(_07796_),
    .X(_07810_));
 sky130_fd_sc_hd__a22o_1 _15327_ (.A1(_07043_),
    .A2(_06972_),
    .B1(_07493_),
    .B2(_07044_),
    .X(_07811_));
 sky130_fd_sc_hd__and2_1 _15328_ (.A(_06970_),
    .B(\wfg_stim_sine_top.wfg_stim_sine.sin_17[1] ),
    .X(_07812_));
 sky130_fd_sc_hd__a32o_1 _15329_ (.A1(_06604_),
    .A2(_06989_),
    .A3(_07811_),
    .B1(_07812_),
    .B2(_07565_),
    .X(_07813_));
 sky130_fd_sc_hd__and3_1 _15330_ (.A(\wfg_stim_sine_top.gain_val_q[3] ),
    .B(_07689_),
    .C(_07813_),
    .X(_07814_));
 sky130_fd_sc_hd__a21oi_1 _15331_ (.A1(\wfg_stim_sine_top.gain_val_q[3] ),
    .A2(_07689_),
    .B1(_07813_),
    .Y(_07815_));
 sky130_fd_sc_hd__or2_1 _15332_ (.A(_07814_),
    .B(_07815_),
    .X(_07816_));
 sky130_fd_sc_hd__nand2_1 _15333_ (.A(_06605_),
    .B(_07493_),
    .Y(_07817_));
 sky130_fd_sc_hd__a21boi_1 _15334_ (.A1(_07565_),
    .A2(_07800_),
    .B1_N(_07799_),
    .Y(_07818_));
 sky130_fd_sc_hd__xor2_1 _15335_ (.A(_07817_),
    .B(_07818_),
    .X(_07819_));
 sky130_fd_sc_hd__nor2_1 _15336_ (.A(_07816_),
    .B(_07819_),
    .Y(_07820_));
 sky130_fd_sc_hd__and2_1 _15337_ (.A(_07803_),
    .B(_07805_),
    .X(_07821_));
 sky130_fd_sc_hd__nor2_1 _15338_ (.A(_07806_),
    .B(_07821_),
    .Y(_07822_));
 sky130_fd_sc_hd__o21ai_1 _15339_ (.A1(_07814_),
    .A2(_07820_),
    .B1(_07822_),
    .Y(_07823_));
 sky130_fd_sc_hd__nor2_1 _15340_ (.A(_07822_),
    .B(_07814_),
    .Y(_07824_));
 sky130_fd_sc_hd__or2_1 _15341_ (.A(_06605_),
    .B(_06972_),
    .X(_07825_));
 sky130_fd_sc_hd__a221o_1 _15342_ (.A1(_07816_),
    .A2(_07819_),
    .B1(_07825_),
    .B2(_07767_),
    .C1(_07001_),
    .X(_07826_));
 sky130_fd_sc_hd__or4_1 _15343_ (.A(_07324_),
    .B(_07824_),
    .C(_07820_),
    .D(_07826_),
    .X(_07827_));
 sky130_fd_sc_hd__o2bb2a_1 _15344_ (.A1_N(_07823_),
    .A2_N(_07827_),
    .B1(_07798_),
    .B2(_07807_),
    .X(_07828_));
 sky130_fd_sc_hd__a221o_1 _15345_ (.A1(_07798_),
    .A2(_07807_),
    .B1(_07809_),
    .B2(_07810_),
    .C1(_07828_),
    .X(_07829_));
 sky130_fd_sc_hd__o22a_1 _15346_ (.A1(_07775_),
    .A2(_07781_),
    .B1(_07810_),
    .B2(_07809_),
    .X(_07830_));
 sky130_fd_sc_hd__and4_1 _15347_ (.A(_07788_),
    .B(_07789_),
    .C(_07829_),
    .D(_07830_),
    .X(_07831_));
 sky130_fd_sc_hd__or2_1 _15348_ (.A(_07786_),
    .B(_07784_),
    .X(_07832_));
 sky130_fd_sc_hd__o221a_1 _15349_ (.A1(_07703_),
    .A2(_07736_),
    .B1(_07787_),
    .B2(_07831_),
    .C1(_07832_),
    .X(_07833_));
 sky130_fd_sc_hd__a211o_1 _15350_ (.A1(_07586_),
    .A2(_07589_),
    .B1(_07587_),
    .C1(_07588_),
    .X(_07834_));
 sky130_fd_sc_hd__a21oi_1 _15351_ (.A1(_07634_),
    .A2(_07637_),
    .B1(_07655_),
    .Y(_07835_));
 sky130_fd_sc_hd__a31o_1 _15352_ (.A1(_07200_),
    .A2(_06748_),
    .A3(_07656_),
    .B1(_07835_),
    .X(_07836_));
 sky130_fd_sc_hd__o21a_1 _15353_ (.A1(_07576_),
    .A2(_07582_),
    .B1(_07581_),
    .X(_07837_));
 sky130_fd_sc_hd__nand3_1 _15354_ (.A(_07653_),
    .B(_07658_),
    .C(_07659_),
    .Y(_07838_));
 sky130_fd_sc_hd__o211ai_1 _15355_ (.A1(_07583_),
    .A2(_07837_),
    .B1(_07653_),
    .C1(_07838_),
    .Y(_07839_));
 sky130_fd_sc_hd__a211oi_1 _15356_ (.A1(_07653_),
    .A2(_07838_),
    .B1(_07583_),
    .C1(_07837_),
    .Y(_07840_));
 sky130_fd_sc_hd__a21o_1 _15357_ (.A1(_07836_),
    .A2(_07839_),
    .B1(_07840_),
    .X(_07841_));
 sky130_fd_sc_hd__a21o_1 _15358_ (.A1(_07590_),
    .A2(_07834_),
    .B1(_07841_),
    .X(_07842_));
 sky130_fd_sc_hd__nand3_1 _15359_ (.A(_07590_),
    .B(_07834_),
    .C(_07841_),
    .Y(_07843_));
 sky130_fd_sc_hd__o211a_1 _15360_ (.A1(_07665_),
    .A2(_07701_),
    .B1(_07842_),
    .C1(_07843_),
    .X(_07844_));
 sky130_fd_sc_hd__or2b_1 _15361_ (.A(_07840_),
    .B_N(_07839_),
    .X(_07845_));
 sky130_fd_sc_hd__xnor2_1 _15362_ (.A(_07836_),
    .B(_07845_),
    .Y(_07846_));
 sky130_fd_sc_hd__a21o_1 _15363_ (.A1(_07628_),
    .A2(_07664_),
    .B1(_07662_),
    .X(_07847_));
 sky130_fd_sc_hd__xor2_1 _15364_ (.A(_07846_),
    .B(_07847_),
    .X(_07848_));
 sky130_fd_sc_hd__o211ai_4 _15365_ (.A1(_07737_),
    .A2(_07833_),
    .B1(_07844_),
    .C1(_07848_),
    .Y(_07849_));
 sky130_fd_sc_hd__nand2_1 _15366_ (.A(_07846_),
    .B(_07847_),
    .Y(_07850_));
 sky130_fd_sc_hd__a21bo_1 _15367_ (.A1(_07843_),
    .A2(_07850_),
    .B1_N(_07842_),
    .X(_07851_));
 sky130_fd_sc_hd__o211a_1 _15368_ (.A1(_07536_),
    .A2(_07591_),
    .B1(_07586_),
    .C1(_07590_),
    .X(_07852_));
 sky130_fd_sc_hd__o21a_1 _15369_ (.A1(_07336_),
    .A2(_07483_),
    .B1(_07537_),
    .X(_07853_));
 sky130_fd_sc_hd__a311o_1 _15370_ (.A1(_07593_),
    .A2(_07849_),
    .A3(_07851_),
    .B1(_07852_),
    .C1(_07853_),
    .X(_07854_));
 sky130_fd_sc_hd__xnor2_1 _15371_ (.A(_07339_),
    .B(_07337_),
    .Y(_07855_));
 sky130_fd_sc_hd__nor2_1 _15372_ (.A(_07280_),
    .B(_07341_),
    .Y(_07856_));
 sky130_fd_sc_hd__nand2_1 _15373_ (.A(_07855_),
    .B(_07856_),
    .Y(_07857_));
 sky130_fd_sc_hd__a211o_1 _15374_ (.A1(_07539_),
    .A2(_07854_),
    .B1(_07857_),
    .C1(_07477_),
    .X(_07858_));
 sky130_fd_sc_hd__a21oi_1 _15375_ (.A1(_07449_),
    .A2(_07457_),
    .B1(_07459_),
    .Y(_07859_));
 sky130_fd_sc_hd__or2_1 _15376_ (.A(_06607_),
    .B(_07859_),
    .X(_07860_));
 sky130_fd_sc_hd__xnor2_1 _15377_ (.A(_06606_),
    .B(_07859_),
    .Y(_07861_));
 sky130_fd_sc_hd__or2_1 _15378_ (.A(_06602_),
    .B(_07861_),
    .X(_07862_));
 sky130_fd_sc_hd__xnor2_1 _15379_ (.A(_06903_),
    .B(_06909_),
    .Y(_07863_));
 sky130_fd_sc_hd__a21o_2 _15380_ (.A1(_07421_),
    .A2(_07428_),
    .B1(_07863_),
    .X(_07864_));
 sky130_fd_sc_hd__nand3_1 _15381_ (.A(_07863_),
    .B(_07421_),
    .C(_07428_),
    .Y(_07865_));
 sky130_fd_sc_hd__or2b_1 _15382_ (.A(_07434_),
    .B_N(_07437_),
    .X(_07866_));
 sky130_fd_sc_hd__a32o_1 _15383_ (.A1(_06468_),
    .A2(_06430_),
    .A3(_07424_),
    .B1(_07423_),
    .B2(_06748_),
    .X(_07867_));
 sky130_fd_sc_hd__o21ai_1 _15384_ (.A1(_06914_),
    .A2(_06915_),
    .B1(_06916_),
    .Y(_07868_));
 sky130_fd_sc_hd__nand2_1 _15385_ (.A(_06917_),
    .B(_07868_),
    .Y(_07869_));
 sky130_fd_sc_hd__xnor2_1 _15386_ (.A(_07867_),
    .B(_07869_),
    .Y(_07870_));
 sky130_fd_sc_hd__xor2_2 _15387_ (.A(_07866_),
    .B(_07870_),
    .X(_07871_));
 sky130_fd_sc_hd__nand3_4 _15388_ (.A(_07864_),
    .B(_07865_),
    .C(_07871_),
    .Y(_07872_));
 sky130_fd_sc_hd__a21o_1 _15389_ (.A1(_07864_),
    .A2(_07865_),
    .B1(_07871_),
    .X(_07873_));
 sky130_fd_sc_hd__o211ai_4 _15390_ (.A1(_07431_),
    .A2(_07444_),
    .B1(_07872_),
    .C1(_07873_),
    .Y(_07874_));
 sky130_fd_sc_hd__a211o_1 _15391_ (.A1(_07872_),
    .A2(_07873_),
    .B1(_07431_),
    .C1(_07444_),
    .X(_07875_));
 sky130_fd_sc_hd__nand2_1 _15392_ (.A(_07454_),
    .B(_07455_),
    .Y(_07876_));
 sky130_fd_sc_hd__nand2_1 _15393_ (.A(_06648_),
    .B(_07456_),
    .Y(_07877_));
 sky130_fd_sc_hd__o21bai_2 _15394_ (.A1(_07433_),
    .A2(_07441_),
    .B1_N(_07440_),
    .Y(_07878_));
 sky130_fd_sc_hd__xnor2_1 _15395_ (.A(_06545_),
    .B(_06933_),
    .Y(_07879_));
 sky130_fd_sc_hd__a31o_1 _15396_ (.A1(_06551_),
    .A2(_06453_),
    .A3(_07451_),
    .B1(_07450_),
    .X(_07880_));
 sky130_fd_sc_hd__xor2_1 _15397_ (.A(_07879_),
    .B(_07880_),
    .X(_07881_));
 sky130_fd_sc_hd__xnor2_1 _15398_ (.A(_06543_),
    .B(_07881_),
    .Y(_07882_));
 sky130_fd_sc_hd__xnor2_1 _15399_ (.A(_07878_),
    .B(_07882_),
    .Y(_07883_));
 sky130_fd_sc_hd__a21o_1 _15400_ (.A1(_07876_),
    .A2(_07877_),
    .B1(_07883_),
    .X(_07884_));
 sky130_fd_sc_hd__nand3_1 _15401_ (.A(_07876_),
    .B(_07877_),
    .C(_07883_),
    .Y(_07885_));
 sky130_fd_sc_hd__nand4_2 _15402_ (.A(_07874_),
    .B(_07875_),
    .C(_07884_),
    .D(_07885_),
    .Y(_07886_));
 sky130_fd_sc_hd__a22o_1 _15403_ (.A1(_07874_),
    .A2(_07875_),
    .B1(_07884_),
    .B2(_07885_),
    .X(_07887_));
 sky130_fd_sc_hd__o211ai_4 _15404_ (.A1(_07446_),
    .A2(_07461_),
    .B1(_07886_),
    .C1(_07887_),
    .Y(_07888_));
 sky130_fd_sc_hd__a211o_1 _15405_ (.A1(_07886_),
    .A2(_07887_),
    .B1(_07446_),
    .C1(_07461_),
    .X(_07889_));
 sky130_fd_sc_hd__xor2_1 _15406_ (.A(_06601_),
    .B(_07861_),
    .X(_07890_));
 sky130_fd_sc_hd__nand3_1 _15407_ (.A(_07888_),
    .B(_07889_),
    .C(_07890_),
    .Y(_07891_));
 sky130_fd_sc_hd__inv_2 _15408_ (.A(_07874_),
    .Y(_07892_));
 sky130_fd_sc_hd__and4_1 _15409_ (.A(_07874_),
    .B(_07875_),
    .C(_07884_),
    .D(_07885_),
    .X(_07893_));
 sky130_fd_sc_hd__and3_1 _15410_ (.A(_06912_),
    .B(_06913_),
    .C(_06923_),
    .X(_07894_));
 sky130_fd_sc_hd__a21oi_2 _15411_ (.A1(_06912_),
    .A2(_06913_),
    .B1(_06923_),
    .Y(_07895_));
 sky130_fd_sc_hd__a211o_2 _15412_ (.A1(_07864_),
    .A2(_07872_),
    .B1(_07894_),
    .C1(_07895_),
    .X(_07896_));
 sky130_fd_sc_hd__o211ai_4 _15413_ (.A1(_07894_),
    .A2(_07895_),
    .B1(_07864_),
    .C1(_07872_),
    .Y(_07897_));
 sky130_fd_sc_hd__nand2_1 _15414_ (.A(_07879_),
    .B(_07880_),
    .Y(_07898_));
 sky130_fd_sc_hd__nand2_1 _15415_ (.A(_06648_),
    .B(_07881_),
    .Y(_07899_));
 sky130_fd_sc_hd__a32o_1 _15416_ (.A1(_06917_),
    .A2(_07867_),
    .A3(_07868_),
    .B1(_07870_),
    .B2(_07866_),
    .X(_07900_));
 sky130_fd_sc_hd__xnor2_1 _15417_ (.A(_06648_),
    .B(_06937_),
    .Y(_07901_));
 sky130_fd_sc_hd__xnor2_1 _15418_ (.A(_07900_),
    .B(_07901_),
    .Y(_07902_));
 sky130_fd_sc_hd__a21o_1 _15419_ (.A1(_07898_),
    .A2(_07899_),
    .B1(_07902_),
    .X(_07903_));
 sky130_fd_sc_hd__nand3_1 _15420_ (.A(_07898_),
    .B(_07899_),
    .C(_07902_),
    .Y(_07904_));
 sky130_fd_sc_hd__nand4_4 _15421_ (.A(_07896_),
    .B(_07897_),
    .C(_07903_),
    .D(_07904_),
    .Y(_07905_));
 sky130_fd_sc_hd__a22o_1 _15422_ (.A1(_07896_),
    .A2(_07897_),
    .B1(_07903_),
    .B2(_07904_),
    .X(_07906_));
 sky130_fd_sc_hd__o211ai_4 _15423_ (.A1(_07892_),
    .A2(_07893_),
    .B1(_07905_),
    .C1(_07906_),
    .Y(_07907_));
 sky130_fd_sc_hd__a211o_1 _15424_ (.A1(_07905_),
    .A2(_07906_),
    .B1(_07892_),
    .C1(_07893_),
    .X(_07908_));
 sky130_fd_sc_hd__a21boi_1 _15425_ (.A1(_07878_),
    .A2(_07882_),
    .B1_N(_07884_),
    .Y(_07909_));
 sky130_fd_sc_hd__xnor2_1 _15426_ (.A(_06606_),
    .B(_07909_),
    .Y(_07910_));
 sky130_fd_sc_hd__xor2_1 _15427_ (.A(_06601_),
    .B(_07910_),
    .X(_07911_));
 sky130_fd_sc_hd__and3_1 _15428_ (.A(_07907_),
    .B(_07908_),
    .C(_07911_),
    .X(_07912_));
 sky130_fd_sc_hd__a21oi_1 _15429_ (.A1(_07907_),
    .A2(_07908_),
    .B1(_07911_),
    .Y(_07913_));
 sky130_fd_sc_hd__a211oi_2 _15430_ (.A1(_07888_),
    .A2(_07891_),
    .B1(_07912_),
    .C1(_07913_),
    .Y(_07914_));
 sky130_fd_sc_hd__o211a_1 _15431_ (.A1(_07912_),
    .A2(_07913_),
    .B1(_07888_),
    .C1(_07891_),
    .X(_07915_));
 sky130_fd_sc_hd__a211oi_2 _15432_ (.A1(_07860_),
    .A2(_07862_),
    .B1(_07914_),
    .C1(_07915_),
    .Y(_07916_));
 sky130_fd_sc_hd__o211a_1 _15433_ (.A1(_07914_),
    .A2(_07915_),
    .B1(_07860_),
    .C1(_07862_),
    .X(_07917_));
 sky130_fd_sc_hd__nand3_1 _15434_ (.A(_07463_),
    .B(_07464_),
    .C(_07467_),
    .Y(_07918_));
 sky130_fd_sc_hd__and3_1 _15435_ (.A(_07888_),
    .B(_07889_),
    .C(_07890_),
    .X(_07919_));
 sky130_fd_sc_hd__a21oi_1 _15436_ (.A1(_07888_),
    .A2(_07889_),
    .B1(_07890_),
    .Y(_07920_));
 sky130_fd_sc_hd__a211o_1 _15437_ (.A1(_07463_),
    .A2(_07918_),
    .B1(_07919_),
    .C1(_07920_),
    .X(_07921_));
 sky130_fd_sc_hd__nor2_1 _15438_ (.A(_06653_),
    .B(_07465_),
    .Y(_07922_));
 sky130_fd_sc_hd__nor2_1 _15439_ (.A(_06602_),
    .B(_07466_),
    .Y(_07923_));
 sky130_fd_sc_hd__o211ai_1 _15440_ (.A1(_07919_),
    .A2(_07920_),
    .B1(_07463_),
    .C1(_07918_),
    .Y(_07924_));
 sky130_fd_sc_hd__o211ai_2 _15441_ (.A1(_07922_),
    .A2(_07923_),
    .B1(_07921_),
    .C1(_07924_),
    .Y(_07925_));
 sky130_fd_sc_hd__o211a_1 _15442_ (.A1(_07916_),
    .A2(_07917_),
    .B1(_07921_),
    .C1(_07925_),
    .X(_07926_));
 sky130_fd_sc_hd__a211o_1 _15443_ (.A1(_07921_),
    .A2(_07925_),
    .B1(_07916_),
    .C1(_07917_),
    .X(_07927_));
 sky130_fd_sc_hd__or2b_1 _15444_ (.A(_07926_),
    .B_N(_07927_),
    .X(_07928_));
 sky130_fd_sc_hd__a211o_1 _15445_ (.A1(_07921_),
    .A2(_07924_),
    .B1(_07922_),
    .C1(_07923_),
    .X(_07929_));
 sky130_fd_sc_hd__and2_1 _15446_ (.A(_07925_),
    .B(_07929_),
    .X(_07930_));
 sky130_fd_sc_hd__nor2_1 _15447_ (.A(_07470_),
    .B(_07472_),
    .Y(_07931_));
 sky130_fd_sc_hd__xnor2_2 _15448_ (.A(_07930_),
    .B(_07931_),
    .Y(_07932_));
 sky130_fd_sc_hd__or2b_1 _15449_ (.A(_07928_),
    .B_N(_07932_),
    .X(_07933_));
 sky130_fd_sc_hd__a21o_1 _15450_ (.A1(_07481_),
    .A2(_07858_),
    .B1(_07933_),
    .X(_07934_));
 sky130_fd_sc_hd__or2b_1 _15451_ (.A(_07931_),
    .B_N(_07930_),
    .X(_07935_));
 sky130_fd_sc_hd__a21o_1 _15452_ (.A1(_07927_),
    .A2(_07935_),
    .B1(_07926_),
    .X(_07936_));
 sky130_fd_sc_hd__nand3_1 _15453_ (.A(_07907_),
    .B(_07908_),
    .C(_07911_),
    .Y(_07937_));
 sky130_fd_sc_hd__a21oi_1 _15454_ (.A1(_06927_),
    .A2(_06928_),
    .B1(_06944_),
    .Y(_07938_));
 sky130_fd_sc_hd__and3_1 _15455_ (.A(_06927_),
    .B(_06928_),
    .C(_06944_),
    .X(_07939_));
 sky130_fd_sc_hd__a211o_2 _15456_ (.A1(_07896_),
    .A2(_07905_),
    .B1(_07938_),
    .C1(_07939_),
    .X(_07940_));
 sky130_fd_sc_hd__o211ai_1 _15457_ (.A1(_07939_),
    .A2(_07938_),
    .B1(_07905_),
    .C1(_07896_),
    .Y(_07941_));
 sky130_fd_sc_hd__a21boi_1 _15458_ (.A1(_07900_),
    .A2(_07901_),
    .B1_N(_07903_),
    .Y(_07942_));
 sky130_fd_sc_hd__xnor2_1 _15459_ (.A(_06606_),
    .B(_07942_),
    .Y(_07943_));
 sky130_fd_sc_hd__xor2_1 _15460_ (.A(_06601_),
    .B(_07943_),
    .X(_07944_));
 sky130_fd_sc_hd__and3_1 _15461_ (.A(_07940_),
    .B(_07941_),
    .C(_07944_),
    .X(_07945_));
 sky130_fd_sc_hd__a21oi_1 _15462_ (.A1(_07940_),
    .A2(_07941_),
    .B1(_07944_),
    .Y(_07946_));
 sky130_fd_sc_hd__a211o_1 _15463_ (.A1(_07907_),
    .A2(_07937_),
    .B1(_07945_),
    .C1(_07946_),
    .X(_07947_));
 sky130_fd_sc_hd__nor2_1 _15464_ (.A(_06653_),
    .B(_07909_),
    .Y(_07948_));
 sky130_fd_sc_hd__nor2_1 _15465_ (.A(_06603_),
    .B(_07910_),
    .Y(_07949_));
 sky130_fd_sc_hd__o211ai_2 _15466_ (.A1(_07945_),
    .A2(_07946_),
    .B1(_07907_),
    .C1(_07937_),
    .Y(_07950_));
 sky130_fd_sc_hd__o211ai_2 _15467_ (.A1(_07948_),
    .A2(_07949_),
    .B1(_07947_),
    .C1(_07950_),
    .Y(_07951_));
 sky130_fd_sc_hd__or2_1 _15468_ (.A(_06653_),
    .B(_07942_),
    .X(_07952_));
 sky130_fd_sc_hd__or2_1 _15469_ (.A(_06603_),
    .B(_07943_),
    .X(_07953_));
 sky130_fd_sc_hd__nand3_1 _15470_ (.A(_07940_),
    .B(_07941_),
    .C(_07944_),
    .Y(_07954_));
 sky130_fd_sc_hd__o21ba_1 _15471_ (.A1(_06947_),
    .A2(_06948_),
    .B1_N(_06953_),
    .X(_07955_));
 sky130_fd_sc_hd__a211oi_4 _15472_ (.A1(_07940_),
    .A2(_07954_),
    .B1(_06954_),
    .C1(_07955_),
    .Y(_07956_));
 sky130_fd_sc_hd__o211a_1 _15473_ (.A1(_06954_),
    .A2(_07955_),
    .B1(_07940_),
    .C1(_07954_),
    .X(_07957_));
 sky130_fd_sc_hd__a211oi_4 _15474_ (.A1(_07952_),
    .A2(_07953_),
    .B1(_07956_),
    .C1(_07957_),
    .Y(_07958_));
 sky130_fd_sc_hd__o211a_1 _15475_ (.A1(_07956_),
    .A2(_07957_),
    .B1(_07952_),
    .C1(_07953_),
    .X(_07959_));
 sky130_fd_sc_hd__a211oi_1 _15476_ (.A1(_07947_),
    .A2(_07951_),
    .B1(_07958_),
    .C1(_07959_),
    .Y(_07960_));
 sky130_fd_sc_hd__a211o_1 _15477_ (.A1(_07947_),
    .A2(_07950_),
    .B1(_07948_),
    .C1(_07949_),
    .X(_07961_));
 sky130_fd_sc_hd__o211ai_1 _15478_ (.A1(_07914_),
    .A2(_07916_),
    .B1(_07951_),
    .C1(_07961_),
    .Y(_07962_));
 sky130_fd_sc_hd__inv_2 _15479_ (.A(_07962_),
    .Y(_07963_));
 sky130_fd_sc_hd__o211a_1 _15480_ (.A1(_07958_),
    .A2(_07959_),
    .B1(_07947_),
    .C1(_07951_),
    .X(_07964_));
 sky130_fd_sc_hd__o21bai_1 _15481_ (.A1(_07960_),
    .A2(_07963_),
    .B1_N(_07964_),
    .Y(_07965_));
 sky130_fd_sc_hd__or2_1 _15482_ (.A(_07960_),
    .B(_07964_),
    .X(_07966_));
 sky130_fd_sc_hd__a211o_1 _15483_ (.A1(_07951_),
    .A2(_07961_),
    .B1(_07914_),
    .C1(_07916_),
    .X(_07967_));
 sky130_fd_sc_hd__nand2_1 _15484_ (.A(_07962_),
    .B(_07967_),
    .Y(_07968_));
 sky130_fd_sc_hd__o21a_1 _15485_ (.A1(_07966_),
    .A2(_07968_),
    .B1(_07965_),
    .X(_07969_));
 sky130_fd_sc_hd__a31o_2 _15486_ (.A1(_07934_),
    .A2(_07936_),
    .A3(_07965_),
    .B1(_07969_),
    .X(_07970_));
 sky130_fd_sc_hd__nand2_1 _15487_ (.A(_06958_),
    .B(_06960_),
    .Y(_07971_));
 sky130_fd_sc_hd__and2_1 _15488_ (.A(_06961_),
    .B(_07971_),
    .X(_07972_));
 sky130_fd_sc_hd__o21ai_1 _15489_ (.A1(_07956_),
    .A2(_07958_),
    .B1(_07972_),
    .Y(_07973_));
 sky130_fd_sc_hd__or3_1 _15490_ (.A(_07956_),
    .B(_07958_),
    .C(_07972_),
    .X(_07974_));
 sky130_fd_sc_hd__nand2_1 _15491_ (.A(_07973_),
    .B(_07974_),
    .Y(_07975_));
 sky130_fd_sc_hd__or3_2 _15492_ (.A(_06964_),
    .B(_07970_),
    .C(_07975_),
    .X(_07976_));
 sky130_fd_sc_hd__a21o_1 _15493_ (.A1(_06963_),
    .A2(_07973_),
    .B1(_06962_),
    .X(_07977_));
 sky130_fd_sc_hd__nor3_2 _15494_ (.A(_06876_),
    .B(_06877_),
    .C(_06885_),
    .Y(_07978_));
 sky130_fd_sc_hd__nor3_1 _15495_ (.A(_06868_),
    .B(_06869_),
    .C(_06873_),
    .Y(_07979_));
 sky130_fd_sc_hd__nand3_2 _15496_ (.A(_06860_),
    .B(_06861_),
    .C(_06865_),
    .Y(_07980_));
 sky130_fd_sc_hd__and3_1 _15497_ (.A(_06482_),
    .B(_06483_),
    .C(_06502_),
    .X(_07981_));
 sky130_fd_sc_hd__a21oi_2 _15498_ (.A1(_06482_),
    .A2(_06483_),
    .B1(_06502_),
    .Y(_07982_));
 sky130_fd_sc_hd__a211oi_4 _15499_ (.A1(_06860_),
    .A2(_07980_),
    .B1(_07981_),
    .C1(_07982_),
    .Y(_07983_));
 sky130_fd_sc_hd__o211a_1 _15500_ (.A1(_07981_),
    .A2(_07982_),
    .B1(_06860_),
    .C1(_07980_),
    .X(_07984_));
 sky130_fd_sc_hd__o21ai_1 _15501_ (.A1(_06822_),
    .A2(_06825_),
    .B1(_06495_),
    .Y(_07985_));
 sky130_fd_sc_hd__a21bo_1 _15502_ (.A1(_06862_),
    .A2(_06864_),
    .B1_N(_07985_),
    .X(_07986_));
 sky130_fd_sc_hd__xnor2_1 _15503_ (.A(_06557_),
    .B(_07986_),
    .Y(_07987_));
 sky130_fd_sc_hd__xnor2_1 _15504_ (.A(_06555_),
    .B(_07987_),
    .Y(_07988_));
 sky130_fd_sc_hd__or3_1 _15505_ (.A(_07983_),
    .B(_07984_),
    .C(_07988_),
    .X(_07989_));
 sky130_fd_sc_hd__o21ai_1 _15506_ (.A1(_07983_),
    .A2(_07984_),
    .B1(_07988_),
    .Y(_07990_));
 sky130_fd_sc_hd__o211a_1 _15507_ (.A1(_06868_),
    .A2(_07979_),
    .B1(_07989_),
    .C1(_07990_),
    .X(_07991_));
 sky130_fd_sc_hd__a211oi_1 _15508_ (.A1(_07989_),
    .A2(_07990_),
    .B1(_06868_),
    .C1(_07979_),
    .Y(_07992_));
 sky130_fd_sc_hd__and2_1 _15509_ (.A(_06649_),
    .B(_06871_),
    .X(_07993_));
 sky130_fd_sc_hd__a21oi_1 _15510_ (.A1(_06555_),
    .A2(_06872_),
    .B1(_07993_),
    .Y(_07994_));
 sky130_fd_sc_hd__xnor2_1 _15511_ (.A(_06607_),
    .B(_07994_),
    .Y(_07995_));
 sky130_fd_sc_hd__or2_1 _15512_ (.A(_06601_),
    .B(_07995_),
    .X(_07996_));
 sky130_fd_sc_hd__nand2_1 _15513_ (.A(_06602_),
    .B(_07995_),
    .Y(_07997_));
 sky130_fd_sc_hd__nand2_1 _15514_ (.A(_07996_),
    .B(_07997_),
    .Y(_07998_));
 sky130_fd_sc_hd__o21ai_2 _15515_ (.A1(_07991_),
    .A2(_07992_),
    .B1(_07998_),
    .Y(_07999_));
 sky130_fd_sc_hd__or3_2 _15516_ (.A(_07991_),
    .B(_07992_),
    .C(_07998_),
    .X(_08000_));
 sky130_fd_sc_hd__o211ai_4 _15517_ (.A1(_06876_),
    .A2(_07978_),
    .B1(_07999_),
    .C1(_08000_),
    .Y(_08001_));
 sky130_fd_sc_hd__a211o_1 _15518_ (.A1(_08000_),
    .A2(_07999_),
    .B1(_07978_),
    .C1(_06876_),
    .X(_08002_));
 sky130_fd_sc_hd__o211ai_2 _15519_ (.A1(_06880_),
    .A2(_06883_),
    .B1(_08001_),
    .C1(_08002_),
    .Y(_08003_));
 sky130_fd_sc_hd__or2_1 _15520_ (.A(_06653_),
    .B(_07994_),
    .X(_08004_));
 sky130_fd_sc_hd__inv_2 _15521_ (.A(_07991_),
    .Y(_08005_));
 sky130_fd_sc_hd__nor3_1 _15522_ (.A(_07983_),
    .B(_07984_),
    .C(_07988_),
    .Y(_08006_));
 sky130_fd_sc_hd__o21ai_1 _15523_ (.A1(_06533_),
    .A2(_06535_),
    .B1(_06561_),
    .Y(_08007_));
 sky130_fd_sc_hd__o211a_1 _15524_ (.A1(_07983_),
    .A2(_08006_),
    .B1(_06562_),
    .C1(_08007_),
    .X(_08008_));
 sky130_fd_sc_hd__a211oi_1 _15525_ (.A1(_06562_),
    .A2(_08007_),
    .B1(_07983_),
    .C1(_08006_),
    .Y(_08009_));
 sky130_fd_sc_hd__and2_1 _15526_ (.A(_06649_),
    .B(_07986_),
    .X(_08010_));
 sky130_fd_sc_hd__a21oi_1 _15527_ (.A1(_06556_),
    .A2(_07987_),
    .B1(_08010_),
    .Y(_08011_));
 sky130_fd_sc_hd__nor2_1 _15528_ (.A(_06607_),
    .B(_08011_),
    .Y(_08012_));
 sky130_fd_sc_hd__and2_1 _15529_ (.A(_06607_),
    .B(_08011_),
    .X(_08013_));
 sky130_fd_sc_hd__or2_1 _15530_ (.A(_08012_),
    .B(_08013_),
    .X(_08014_));
 sky130_fd_sc_hd__nor2_1 _15531_ (.A(_06602_),
    .B(_08014_),
    .Y(_08015_));
 sky130_fd_sc_hd__and2_1 _15532_ (.A(_06602_),
    .B(_08014_),
    .X(_08016_));
 sky130_fd_sc_hd__or2_1 _15533_ (.A(_08015_),
    .B(_08016_),
    .X(_08017_));
 sky130_fd_sc_hd__nor3_1 _15534_ (.A(_08008_),
    .B(_08009_),
    .C(_08017_),
    .Y(_08018_));
 sky130_fd_sc_hd__o21a_1 _15535_ (.A1(_08008_),
    .A2(_08009_),
    .B1(_08017_),
    .X(_08019_));
 sky130_fd_sc_hd__a211oi_2 _15536_ (.A1(_08005_),
    .A2(_08000_),
    .B1(_08018_),
    .C1(_08019_),
    .Y(_08020_));
 sky130_fd_sc_hd__o211a_1 _15537_ (.A1(_08018_),
    .A2(_08019_),
    .B1(_08005_),
    .C1(_08000_),
    .X(_08021_));
 sky130_fd_sc_hd__a211oi_2 _15538_ (.A1(_08004_),
    .A2(_07996_),
    .B1(_08020_),
    .C1(_08021_),
    .Y(_08022_));
 sky130_fd_sc_hd__o211a_1 _15539_ (.A1(_08020_),
    .A2(_08021_),
    .B1(_08004_),
    .C1(_07996_),
    .X(_08023_));
 sky130_fd_sc_hd__a211o_1 _15540_ (.A1(_08001_),
    .A2(_08003_),
    .B1(_08022_),
    .C1(_08023_),
    .X(_08024_));
 sky130_fd_sc_hd__o211ai_1 _15541_ (.A1(_08022_),
    .A2(_08023_),
    .B1(_08001_),
    .C1(_08003_),
    .Y(_08025_));
 sky130_fd_sc_hd__nor2_1 _15542_ (.A(_06888_),
    .B(_06890_),
    .Y(_08026_));
 sky130_fd_sc_hd__a211o_1 _15543_ (.A1(_08001_),
    .A2(_08002_),
    .B1(_06880_),
    .C1(_06883_),
    .X(_08027_));
 sky130_fd_sc_hd__and2_1 _15544_ (.A(_08003_),
    .B(_08027_),
    .X(_08028_));
 sky130_fd_sc_hd__and2b_1 _15545_ (.A_N(_08026_),
    .B(_08028_),
    .X(_08029_));
 sky130_fd_sc_hd__nand2_1 _15546_ (.A(_08025_),
    .B(_08029_),
    .Y(_08030_));
 sky130_fd_sc_hd__and2_1 _15547_ (.A(_08024_),
    .B(_08030_),
    .X(_08031_));
 sky130_fd_sc_hd__and2_1 _15548_ (.A(_07977_),
    .B(_08031_),
    .X(_08032_));
 sky130_fd_sc_hd__nand2_1 _15549_ (.A(_08024_),
    .B(_08025_),
    .Y(_08033_));
 sky130_fd_sc_hd__xor2_1 _15550_ (.A(_08028_),
    .B(_08026_),
    .X(_08034_));
 sky130_fd_sc_hd__or2_1 _15551_ (.A(_08033_),
    .B(_08034_),
    .X(_08035_));
 sky130_fd_sc_hd__o21a_1 _15552_ (.A1(_06597_),
    .A2(_06598_),
    .B1(_06612_),
    .X(_08036_));
 sky130_fd_sc_hd__nor2_1 _15553_ (.A(_06613_),
    .B(_08036_),
    .Y(_08037_));
 sky130_fd_sc_hd__nor2_1 _15554_ (.A(_08008_),
    .B(_08018_),
    .Y(_08038_));
 sky130_fd_sc_hd__xnor2_1 _15555_ (.A(_08037_),
    .B(_08038_),
    .Y(_08039_));
 sky130_fd_sc_hd__o21a_1 _15556_ (.A1(_08012_),
    .A2(_08015_),
    .B1(_08039_),
    .X(_08040_));
 sky130_fd_sc_hd__nor3_1 _15557_ (.A(_08012_),
    .B(_08015_),
    .C(_08039_),
    .Y(_08041_));
 sky130_fd_sc_hd__or2_1 _15558_ (.A(_08040_),
    .B(_08041_),
    .X(_08042_));
 sky130_fd_sc_hd__nor2_1 _15559_ (.A(_08020_),
    .B(_08022_),
    .Y(_08043_));
 sky130_fd_sc_hd__nor2_1 _15560_ (.A(_08042_),
    .B(_08043_),
    .Y(_08044_));
 sky130_fd_sc_hd__and2_1 _15561_ (.A(_08042_),
    .B(_08043_),
    .X(_08045_));
 sky130_fd_sc_hd__or2_1 _15562_ (.A(_08044_),
    .B(_08045_),
    .X(_08046_));
 sky130_fd_sc_hd__a221oi_4 _15563_ (.A1(_07976_),
    .A2(_08032_),
    .B1(_08035_),
    .B2(_08031_),
    .C1(_08046_),
    .Y(_08047_));
 sky130_fd_sc_hd__and2b_1 _15564_ (.A_N(_08038_),
    .B(_08037_),
    .X(_08048_));
 sky130_fd_sc_hd__xnor2_1 _15565_ (.A(_06662_),
    .B(_06660_),
    .Y(_08049_));
 sky130_fd_sc_hd__o21ai_1 _15566_ (.A1(_08048_),
    .A2(_08040_),
    .B1(_08049_),
    .Y(_08050_));
 sky130_fd_sc_hd__o21ai_1 _15567_ (.A1(_08042_),
    .A2(_08043_),
    .B1(_08050_),
    .Y(_08051_));
 sky130_fd_sc_hd__or3_1 _15568_ (.A(_06704_),
    .B(_06659_),
    .C(_06663_),
    .X(_08052_));
 sky130_fd_sc_hd__and2b_1 _15569_ (.A_N(_06705_),
    .B(_08052_),
    .X(_08053_));
 sky130_fd_sc_hd__or3_1 _15570_ (.A(_08049_),
    .B(_08048_),
    .C(_08040_),
    .X(_08054_));
 sky130_fd_sc_hd__o211a_1 _15571_ (.A1(_08047_),
    .A2(_08051_),
    .B1(_08053_),
    .C1(_08054_),
    .X(_08055_));
 sky130_fd_sc_hd__or2_1 _15572_ (.A(_06705_),
    .B(_08055_),
    .X(_08056_));
 sky130_fd_sc_hd__a21o_1 _15573_ (.A1(_06702_),
    .A2(_06703_),
    .B1(_06700_),
    .X(_08057_));
 sky130_fd_sc_hd__a21o_1 _15574_ (.A1(_06556_),
    .A2(_06668_),
    .B1(_06666_),
    .X(_08058_));
 sky130_fd_sc_hd__a21oi_1 _15575_ (.A1(_06568_),
    .A2(_06680_),
    .B1(_06678_),
    .Y(_08059_));
 sky130_fd_sc_hd__xnor2_1 _15576_ (.A(_08058_),
    .B(_08059_),
    .Y(_08060_));
 sky130_fd_sc_hd__xnor2_1 _15577_ (.A(_06669_),
    .B(_06621_),
    .Y(_08061_));
 sky130_fd_sc_hd__o21a_1 _15578_ (.A1(_06621_),
    .A2(_06684_),
    .B1(_06682_),
    .X(_08062_));
 sky130_fd_sc_hd__nor2_1 _15579_ (.A(_06505_),
    .B(_06509_),
    .Y(_08063_));
 sky130_fd_sc_hd__a211o_1 _15580_ (.A1(_06672_),
    .A2(_06674_),
    .B1(_08063_),
    .C1(_06407_),
    .X(_08064_));
 sky130_fd_sc_hd__buf_2 _15581_ (.A(_06600_),
    .X(_08065_));
 sky130_fd_sc_hd__clkbuf_4 _15582_ (.A(_08065_),
    .X(_08066_));
 sky130_fd_sc_hd__o211a_1 _15583_ (.A1(_06406_),
    .A2(_06675_),
    .B1(_08064_),
    .C1(_08066_),
    .X(_08067_));
 sky130_fd_sc_hd__xnor2_1 _15584_ (.A(_06568_),
    .B(_08067_),
    .Y(_08068_));
 sky130_fd_sc_hd__xnor2_1 _15585_ (.A(_08062_),
    .B(_08068_),
    .Y(_08069_));
 sky130_fd_sc_hd__xnor2_1 _15586_ (.A(_08061_),
    .B(_08069_),
    .Y(_08070_));
 sky130_fd_sc_hd__xnor2_1 _15587_ (.A(_08060_),
    .B(_08070_),
    .Y(_08071_));
 sky130_fd_sc_hd__o21ai_1 _15588_ (.A1(_06669_),
    .A2(_06689_),
    .B1(_06687_),
    .Y(_08072_));
 sky130_fd_sc_hd__o21a_1 _15589_ (.A1(_06603_),
    .A2(_06697_),
    .B1(_06695_),
    .X(_08073_));
 sky130_fd_sc_hd__xnor2_1 _15590_ (.A(_08072_),
    .B(_08073_),
    .Y(_08074_));
 sky130_fd_sc_hd__xnor2_1 _15591_ (.A(_08071_),
    .B(_08074_),
    .Y(_08075_));
 sky130_fd_sc_hd__a21boi_1 _15592_ (.A1(_06692_),
    .A2(_06698_),
    .B1_N(_06691_),
    .Y(_08076_));
 sky130_fd_sc_hd__xnor2_1 _15593_ (.A(_06603_),
    .B(_06653_),
    .Y(_08077_));
 sky130_fd_sc_hd__xnor2_1 _15594_ (.A(_08076_),
    .B(_08077_),
    .Y(_08078_));
 sky130_fd_sc_hd__xnor2_1 _15595_ (.A(_08075_),
    .B(_08078_),
    .Y(_08079_));
 sky130_fd_sc_hd__xnor2_2 _15596_ (.A(_08057_),
    .B(_08079_),
    .Y(_08080_));
 sky130_fd_sc_hd__buf_6 _15597_ (.A(_06406_),
    .X(_08081_));
 sky130_fd_sc_hd__clkbuf_8 _15598_ (.A(_08081_),
    .X(_08082_));
 sky130_fd_sc_hd__a21oi_1 _15599_ (.A1(_08056_),
    .A2(_08080_),
    .B1(_08082_),
    .Y(_08083_));
 sky130_fd_sc_hd__o21a_2 _15600_ (.A1(_08056_),
    .A2(_08080_),
    .B1(_08083_),
    .X(_08084_));
 sky130_fd_sc_hd__o22a_1 _15601_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.temp[31] ),
    .A2(_06404_),
    .B1(_06411_),
    .B2(_08084_),
    .X(_00961_));
 sky130_fd_sc_hd__buf_4 _15602_ (.A(_08066_),
    .X(_08085_));
 sky130_fd_sc_hd__or2_1 _15603_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[13] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.sin_17[12] ),
    .X(_08086_));
 sky130_fd_sc_hd__and3_1 _15604_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[14] ),
    .B(_07042_),
    .C(_08086_),
    .X(_08087_));
 sky130_fd_sc_hd__a21oi_1 _15605_ (.A1(_07042_),
    .A2(_08086_),
    .B1(\wfg_stim_sine_top.wfg_stim_sine.sin_17[14] ),
    .Y(_08088_));
 sky130_fd_sc_hd__or2_1 _15606_ (.A(_08087_),
    .B(_08088_),
    .X(_08089_));
 sky130_fd_sc_hd__buf_4 _15607_ (.A(_08089_),
    .X(_08090_));
 sky130_fd_sc_hd__or2_1 _15608_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[12] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.sin_17[11] ),
    .X(_08091_));
 sky130_fd_sc_hd__and3_1 _15609_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[13] ),
    .B(_07307_),
    .C(_08091_),
    .X(_08092_));
 sky130_fd_sc_hd__a21oi_4 _15610_ (.A1(_06421_),
    .A2(_06413_),
    .B1(_08092_),
    .Y(_08093_));
 sky130_fd_sc_hd__xor2_4 _15611_ (.A(_08090_),
    .B(_08093_),
    .X(_08094_));
 sky130_fd_sc_hd__nor2_1 _15612_ (.A(_08090_),
    .B(_08093_),
    .Y(_08095_));
 sky130_fd_sc_hd__a21oi_4 _15613_ (.A1(_06454_),
    .A2(_08094_),
    .B1(_08095_),
    .Y(_08096_));
 sky130_fd_sc_hd__inv_2 _15614_ (.A(_08096_),
    .Y(_08097_));
 sky130_fd_sc_hd__xor2_2 _15615_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[14] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.sin_17[13] ),
    .X(_08098_));
 sky130_fd_sc_hd__xnor2_4 _15616_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[15] ),
    .B(_08098_),
    .Y(_08099_));
 sky130_fd_sc_hd__a21boi_2 _15617_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.sin_17[14] ),
    .A2(_08086_),
    .B1_N(_07042_),
    .Y(_08100_));
 sky130_fd_sc_hd__nand2_1 _15618_ (.A(_08099_),
    .B(_08100_),
    .Y(_08101_));
 sky130_fd_sc_hd__or2_1 _15619_ (.A(_08099_),
    .B(_08100_),
    .X(_08102_));
 sky130_fd_sc_hd__nand2_2 _15620_ (.A(_08101_),
    .B(_08102_),
    .Y(_08103_));
 sky130_fd_sc_hd__mux2_1 _15621_ (.A0(_08097_),
    .A1(_06600_),
    .S(_08103_),
    .X(_08104_));
 sky130_fd_sc_hd__nor2_1 _15622_ (.A(_08099_),
    .B(_08100_),
    .Y(_08105_));
 sky130_fd_sc_hd__a21oi_2 _15623_ (.A1(_06525_),
    .A2(_08101_),
    .B1(_08105_),
    .Y(_08106_));
 sky130_fd_sc_hd__o21a_1 _15624_ (.A1(_06473_),
    .A2(_06463_),
    .B1(_06454_),
    .X(_08107_));
 sky130_fd_sc_hd__a21o_2 _15625_ (.A1(_06510_),
    .A2(_06513_),
    .B1(_08107_),
    .X(_08108_));
 sky130_fd_sc_hd__and2_1 _15626_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[15] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.sin_17[14] ),
    .X(_08109_));
 sky130_fd_sc_hd__nor2_2 _15627_ (.A(_06452_),
    .B(_06440_),
    .Y(_08110_));
 sky130_fd_sc_hd__or3_2 _15628_ (.A(_06410_),
    .B(_08109_),
    .C(_08110_),
    .X(_08111_));
 sky130_fd_sc_hd__o21ai_2 _15629_ (.A1(_08109_),
    .A2(_08110_),
    .B1(_06410_),
    .Y(_08112_));
 sky130_fd_sc_hd__nand2_4 _15630_ (.A(_08111_),
    .B(_08112_),
    .Y(_08113_));
 sky130_fd_sc_hd__xor2_1 _15631_ (.A(_08108_),
    .B(_08113_),
    .X(_08114_));
 sky130_fd_sc_hd__xor2_1 _15632_ (.A(_08106_),
    .B(_08114_),
    .X(_08115_));
 sky130_fd_sc_hd__and2_1 _15633_ (.A(_08104_),
    .B(_08115_),
    .X(_08116_));
 sky130_fd_sc_hd__nor2_1 _15634_ (.A(_08104_),
    .B(_08115_),
    .Y(_08117_));
 sky130_fd_sc_hd__nor2_1 _15635_ (.A(_08116_),
    .B(_08117_),
    .Y(_08118_));
 sky130_fd_sc_hd__xnor2_4 _15636_ (.A(_06472_),
    .B(_08094_),
    .Y(_08119_));
 sky130_fd_sc_hd__a21oi_1 _15637_ (.A1(_07307_),
    .A2(_08091_),
    .B1(_06442_),
    .Y(_08120_));
 sky130_fd_sc_hd__or2_1 _15638_ (.A(_08092_),
    .B(_08120_),
    .X(_08121_));
 sky130_fd_sc_hd__buf_4 _15639_ (.A(_08121_),
    .X(_08122_));
 sky130_fd_sc_hd__xor2_4 _15640_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[11] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.sin_17[10] ),
    .X(_08123_));
 sky130_fd_sc_hd__a21boi_4 _15641_ (.A1(_06422_),
    .A2(_08123_),
    .B1_N(_07511_),
    .Y(_08124_));
 sky130_fd_sc_hd__xnor2_2 _15642_ (.A(_08122_),
    .B(_08124_),
    .Y(_08125_));
 sky130_fd_sc_hd__or2_1 _15643_ (.A(_08122_),
    .B(_08124_),
    .X(_08126_));
 sky130_fd_sc_hd__o21a_4 _15644_ (.A1(_08113_),
    .A2(_08125_),
    .B1(_08126_),
    .X(_08127_));
 sky130_fd_sc_hd__xnor2_1 _15645_ (.A(_08119_),
    .B(_08127_),
    .Y(_08128_));
 sky130_fd_sc_hd__nand2_2 _15646_ (.A(_06453_),
    .B(_06473_),
    .Y(_08129_));
 sky130_fd_sc_hd__nand2_4 _15647_ (.A(_08129_),
    .B(_08111_),
    .Y(_08130_));
 sky130_fd_sc_hd__or2b_1 _15648_ (.A(_08128_),
    .B_N(_08130_),
    .X(_08131_));
 sky130_fd_sc_hd__o21a_1 _15649_ (.A1(_08119_),
    .A2(_08127_),
    .B1(_08131_),
    .X(_08132_));
 sky130_fd_sc_hd__clkinv_2 _15650_ (.A(_08132_),
    .Y(_08133_));
 sky130_fd_sc_hd__xnor2_2 _15651_ (.A(_06410_),
    .B(_08103_),
    .Y(_08134_));
 sky130_fd_sc_hd__xnor2_1 _15652_ (.A(_08134_),
    .B(_08096_),
    .Y(_08135_));
 sky130_fd_sc_hd__mux2_1 _15653_ (.A0(_08133_),
    .A1(_08065_),
    .S(_08135_),
    .X(_08136_));
 sky130_fd_sc_hd__xor2_1 _15654_ (.A(_08118_),
    .B(_08136_),
    .X(_08137_));
 sky130_fd_sc_hd__xor2_1 _15655_ (.A(_08135_),
    .B(_08132_),
    .X(_08138_));
 sky130_fd_sc_hd__or2b_1 _15656_ (.A(_08130_),
    .B_N(_08128_),
    .X(_08139_));
 sky130_fd_sc_hd__nand2_1 _15657_ (.A(_08131_),
    .B(_08139_),
    .Y(_08140_));
 sky130_fd_sc_hd__xor2_4 _15658_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[10] ),
    .B(_06426_),
    .X(_08141_));
 sky130_fd_sc_hd__a21oi_4 _15659_ (.A1(_06413_),
    .A2(_08141_),
    .B1(_07566_),
    .Y(_08142_));
 sky130_fd_sc_hd__xnor2_4 _15660_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[12] ),
    .B(_08123_),
    .Y(_08143_));
 sky130_fd_sc_hd__xnor2_2 _15661_ (.A(_08142_),
    .B(_08143_),
    .Y(_08144_));
 sky130_fd_sc_hd__or2_1 _15662_ (.A(_08142_),
    .B(_08143_),
    .X(_08145_));
 sky130_fd_sc_hd__o21ai_2 _15663_ (.A1(_08099_),
    .A2(_08144_),
    .B1(_08145_),
    .Y(_08146_));
 sky130_fd_sc_hd__xor2_2 _15664_ (.A(_08113_),
    .B(_08125_),
    .X(_08147_));
 sky130_fd_sc_hd__and2_1 _15665_ (.A(_08146_),
    .B(_08147_),
    .X(_08148_));
 sky130_fd_sc_hd__nor2_1 _15666_ (.A(_08146_),
    .B(_08147_),
    .Y(_08149_));
 sky130_fd_sc_hd__nor2_1 _15667_ (.A(_08148_),
    .B(_08149_),
    .Y(_08150_));
 sky130_fd_sc_hd__a21oi_1 _15668_ (.A1(_08108_),
    .A2(_08150_),
    .B1(_08148_),
    .Y(_08151_));
 sky130_fd_sc_hd__nor2_1 _15669_ (.A(_08140_),
    .B(_08151_),
    .Y(_08152_));
 sky130_fd_sc_hd__and2_1 _15670_ (.A(_08140_),
    .B(_08151_),
    .X(_08153_));
 sky130_fd_sc_hd__nor2_1 _15671_ (.A(_08152_),
    .B(_08153_),
    .Y(_08154_));
 sky130_fd_sc_hd__a21o_1 _15672_ (.A1(_06600_),
    .A2(_08154_),
    .B1(_08152_),
    .X(_08155_));
 sky130_fd_sc_hd__nand2_1 _15673_ (.A(_08138_),
    .B(_08155_),
    .Y(_08156_));
 sky130_fd_sc_hd__or2_1 _15674_ (.A(_08138_),
    .B(_08155_),
    .X(_08157_));
 sky130_fd_sc_hd__nand2_1 _15675_ (.A(_08156_),
    .B(_08157_),
    .Y(_08158_));
 sky130_fd_sc_hd__o21ai_1 _15676_ (.A1(_06410_),
    .A2(_08158_),
    .B1(_08156_),
    .Y(_08159_));
 sky130_fd_sc_hd__nand2_1 _15677_ (.A(_08137_),
    .B(_08159_),
    .Y(_08160_));
 sky130_fd_sc_hd__or2_1 _15678_ (.A(_08137_),
    .B(_08159_),
    .X(_08161_));
 sky130_fd_sc_hd__and2_1 _15679_ (.A(_08160_),
    .B(_08161_),
    .X(_08162_));
 sky130_fd_sc_hd__nand2_1 _15680_ (.A(_08085_),
    .B(_08162_),
    .Y(_08163_));
 sky130_fd_sc_hd__or2_1 _15681_ (.A(_08085_),
    .B(_08162_),
    .X(_08164_));
 sky130_fd_sc_hd__xor2_4 _15682_ (.A(_06426_),
    .B(_06744_),
    .X(_08165_));
 sky130_fd_sc_hd__a21oi_4 _15683_ (.A1(_06415_),
    .A2(_08165_),
    .B1(_07601_),
    .Y(_08166_));
 sky130_fd_sc_hd__xnor2_4 _15684_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[11] ),
    .B(_08141_),
    .Y(_08167_));
 sky130_fd_sc_hd__nor2_1 _15685_ (.A(_08166_),
    .B(_08167_),
    .Y(_08168_));
 sky130_fd_sc_hd__xnor2_1 _15686_ (.A(_08166_),
    .B(_08167_),
    .Y(_08169_));
 sky130_fd_sc_hd__nor2_1 _15687_ (.A(_08090_),
    .B(_08169_),
    .Y(_08170_));
 sky130_fd_sc_hd__or2_1 _15688_ (.A(_08168_),
    .B(_08170_),
    .X(_08171_));
 sky130_fd_sc_hd__xor2_2 _15689_ (.A(_08099_),
    .B(_08144_),
    .X(_08172_));
 sky130_fd_sc_hd__nand2_1 _15690_ (.A(_08171_),
    .B(_08172_),
    .Y(_08173_));
 sky130_fd_sc_hd__a21o_1 _15691_ (.A1(_06513_),
    .A2(_06423_),
    .B1(_08087_),
    .X(_08174_));
 sky130_fd_sc_hd__nor2_1 _15692_ (.A(_08168_),
    .B(_08170_),
    .Y(_08175_));
 sky130_fd_sc_hd__xnor2_1 _15693_ (.A(_08175_),
    .B(_08172_),
    .Y(_08176_));
 sky130_fd_sc_hd__nand2_1 _15694_ (.A(_08174_),
    .B(_08176_),
    .Y(_08177_));
 sky130_fd_sc_hd__xnor2_1 _15695_ (.A(_08108_),
    .B(_08150_),
    .Y(_08178_));
 sky130_fd_sc_hd__a21o_1 _15696_ (.A1(_08173_),
    .A2(_08177_),
    .B1(_08178_),
    .X(_08179_));
 sky130_fd_sc_hd__nand3_1 _15697_ (.A(_08178_),
    .B(_08173_),
    .C(_08177_),
    .Y(_08180_));
 sky130_fd_sc_hd__nand2_1 _15698_ (.A(_08179_),
    .B(_08180_),
    .Y(_08181_));
 sky130_fd_sc_hd__o21a_1 _15699_ (.A1(_06410_),
    .A2(_08181_),
    .B1(_08179_),
    .X(_08182_));
 sky130_fd_sc_hd__clkinv_2 _15700_ (.A(_08182_),
    .Y(_08183_));
 sky130_fd_sc_hd__mux2_1 _15701_ (.A0(_08085_),
    .A1(_08183_),
    .S(_08154_),
    .X(_08184_));
 sky130_fd_sc_hd__mux2_1 _15702_ (.A0(_08184_),
    .A1(_08085_),
    .S(_08158_),
    .X(_08185_));
 sky130_fd_sc_hd__nand3_1 _15703_ (.A(_08163_),
    .B(_08164_),
    .C(_08185_),
    .Y(_08186_));
 sky130_fd_sc_hd__a21o_1 _15704_ (.A1(_08066_),
    .A2(_08118_),
    .B1(_08116_),
    .X(_08187_));
 sky130_fd_sc_hd__mux2_1 _15705_ (.A0(_08106_),
    .A1(_06410_),
    .S(_08114_),
    .X(_08188_));
 sky130_fd_sc_hd__a21oi_1 _15706_ (.A1(_06510_),
    .A2(_06513_),
    .B1(_06672_),
    .Y(_08189_));
 sky130_fd_sc_hd__nor2_1 _15707_ (.A(_08107_),
    .B(_08189_),
    .Y(_08190_));
 sky130_fd_sc_hd__xnor2_1 _15708_ (.A(_08188_),
    .B(_08190_),
    .Y(_08191_));
 sky130_fd_sc_hd__nand2_1 _15709_ (.A(_08187_),
    .B(_08191_),
    .Y(_08192_));
 sky130_fd_sc_hd__or2_1 _15710_ (.A(_08187_),
    .B(_08191_),
    .X(_08193_));
 sky130_fd_sc_hd__and2_1 _15711_ (.A(_08192_),
    .B(_08193_),
    .X(_08194_));
 sky130_fd_sc_hd__mux2_1 _15712_ (.A0(_08085_),
    .A1(_08136_),
    .S(_08118_),
    .X(_08195_));
 sky130_fd_sc_hd__xnor2_1 _15713_ (.A(_08194_),
    .B(_08195_),
    .Y(_08196_));
 sky130_fd_sc_hd__a21o_1 _15714_ (.A1(_08160_),
    .A2(_08163_),
    .B1(_08196_),
    .X(_08197_));
 sky130_fd_sc_hd__or2_1 _15715_ (.A(_08174_),
    .B(_08176_),
    .X(_08198_));
 sky130_fd_sc_hd__nand2_1 _15716_ (.A(_08177_),
    .B(_08198_),
    .Y(_08199_));
 sky130_fd_sc_hd__xnor2_4 _15717_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[10] ),
    .B(_08165_),
    .Y(_08200_));
 sky130_fd_sc_hd__xor2_4 _15718_ (.A(_06744_),
    .B(_06736_),
    .X(_08201_));
 sky130_fd_sc_hd__a21boi_4 _15719_ (.A1(_06426_),
    .A2(_08201_),
    .B1_N(_07609_),
    .Y(_08202_));
 sky130_fd_sc_hd__nor2_1 _15720_ (.A(_08200_),
    .B(_08202_),
    .Y(_08203_));
 sky130_fd_sc_hd__xnor2_2 _15721_ (.A(_08200_),
    .B(_08202_),
    .Y(_08204_));
 sky130_fd_sc_hd__nor2_1 _15722_ (.A(_08122_),
    .B(_08204_),
    .Y(_08205_));
 sky130_fd_sc_hd__nor2_1 _15723_ (.A(_08203_),
    .B(_08205_),
    .Y(_08206_));
 sky130_fd_sc_hd__xor2_2 _15724_ (.A(_08090_),
    .B(_08169_),
    .X(_08207_));
 sky130_fd_sc_hd__xnor2_1 _15725_ (.A(_08206_),
    .B(_08207_),
    .Y(_08208_));
 sky130_fd_sc_hd__and2b_1 _15726_ (.A_N(_06454_),
    .B(_08093_),
    .X(_08209_));
 sky130_fd_sc_hd__and2b_1 _15727_ (.A_N(_08093_),
    .B(_06454_),
    .X(_08210_));
 sky130_fd_sc_hd__nor2_1 _15728_ (.A(_08209_),
    .B(_08210_),
    .Y(_08211_));
 sky130_fd_sc_hd__xor2_1 _15729_ (.A(_08130_),
    .B(_08211_),
    .X(_08212_));
 sky130_fd_sc_hd__or2_1 _15730_ (.A(_08203_),
    .B(_08205_),
    .X(_08213_));
 sky130_fd_sc_hd__and2_1 _15731_ (.A(_08213_),
    .B(_08207_),
    .X(_08214_));
 sky130_fd_sc_hd__a21oi_1 _15732_ (.A1(_08208_),
    .A2(_08212_),
    .B1(_08214_),
    .Y(_08215_));
 sky130_fd_sc_hd__xnor2_1 _15733_ (.A(_08199_),
    .B(_08215_),
    .Y(_08216_));
 sky130_fd_sc_hd__a21oi_1 _15734_ (.A1(_08130_),
    .A2(_08211_),
    .B1(_08210_),
    .Y(_08217_));
 sky130_fd_sc_hd__xnor2_1 _15735_ (.A(_08216_),
    .B(_08217_),
    .Y(_08218_));
 sky130_fd_sc_hd__xnor2_1 _15736_ (.A(_08208_),
    .B(_08212_),
    .Y(_08219_));
 sky130_fd_sc_hd__xnor2_4 _15737_ (.A(_06426_),
    .B(_08201_),
    .Y(_08220_));
 sky130_fd_sc_hd__xor2_4 _15738_ (.A(_06736_),
    .B(\wfg_stim_sine_top.wfg_stim_sine.sin_17[6] ),
    .X(_08221_));
 sky130_fd_sc_hd__a21boi_4 _15739_ (.A1(_06747_),
    .A2(_08221_),
    .B1_N(_07668_),
    .Y(_08222_));
 sky130_fd_sc_hd__xnor2_2 _15740_ (.A(_08220_),
    .B(_08222_),
    .Y(_08223_));
 sky130_fd_sc_hd__or2_1 _15741_ (.A(_08220_),
    .B(_08222_),
    .X(_08224_));
 sky130_fd_sc_hd__o21ai_4 _15742_ (.A1(_08143_),
    .A2(_08223_),
    .B1(_08224_),
    .Y(_08225_));
 sky130_fd_sc_hd__xor2_4 _15743_ (.A(_08122_),
    .B(_08204_),
    .X(_08226_));
 sky130_fd_sc_hd__xnor2_1 _15744_ (.A(_08225_),
    .B(_08226_),
    .Y(_08227_));
 sky130_fd_sc_hd__xnor2_1 _15745_ (.A(_08113_),
    .B(_08124_),
    .Y(_08228_));
 sky130_fd_sc_hd__or2b_1 _15746_ (.A(_08228_),
    .B_N(_08108_),
    .X(_08229_));
 sky130_fd_sc_hd__or2b_1 _15747_ (.A(_08108_),
    .B_N(_08228_),
    .X(_08230_));
 sky130_fd_sc_hd__nand2_1 _15748_ (.A(_08229_),
    .B(_08230_),
    .Y(_08231_));
 sky130_fd_sc_hd__nand2_1 _15749_ (.A(_08225_),
    .B(_08226_),
    .Y(_08232_));
 sky130_fd_sc_hd__o21a_1 _15750_ (.A1(_08227_),
    .A2(_08231_),
    .B1(_08232_),
    .X(_08233_));
 sky130_fd_sc_hd__o21a_1 _15751_ (.A1(_08113_),
    .A2(_08124_),
    .B1(_08229_),
    .X(_08234_));
 sky130_fd_sc_hd__xor2_1 _15752_ (.A(_08219_),
    .B(_08233_),
    .X(_08235_));
 sky130_fd_sc_hd__or2b_1 _15753_ (.A(_08234_),
    .B_N(_08235_),
    .X(_08236_));
 sky130_fd_sc_hd__o21a_1 _15754_ (.A1(_08219_),
    .A2(_08233_),
    .B1(_08236_),
    .X(_08237_));
 sky130_fd_sc_hd__or2_1 _15755_ (.A(_08218_),
    .B(_08237_),
    .X(_08238_));
 sky130_fd_sc_hd__nand2_1 _15756_ (.A(_08218_),
    .B(_08237_),
    .Y(_08239_));
 sky130_fd_sc_hd__and2_1 _15757_ (.A(_08238_),
    .B(_08239_),
    .X(_08240_));
 sky130_fd_sc_hd__nand2_1 _15758_ (.A(_08065_),
    .B(_08240_),
    .Y(_08241_));
 sky130_fd_sc_hd__or2_1 _15759_ (.A(_08199_),
    .B(_08215_),
    .X(_08242_));
 sky130_fd_sc_hd__o21ai_1 _15760_ (.A1(_08216_),
    .A2(_08217_),
    .B1(_08242_),
    .Y(_08243_));
 sky130_fd_sc_hd__xor2_1 _15761_ (.A(_08181_),
    .B(_08243_),
    .X(_08244_));
 sky130_fd_sc_hd__a21o_1 _15762_ (.A1(_08238_),
    .A2(_08241_),
    .B1(_08244_),
    .X(_08245_));
 sky130_fd_sc_hd__nand3_1 _15763_ (.A(_08244_),
    .B(_08238_),
    .C(_08241_),
    .Y(_08246_));
 sky130_fd_sc_hd__and2_1 _15764_ (.A(_08245_),
    .B(_08246_),
    .X(_08247_));
 sky130_fd_sc_hd__nand2_1 _15765_ (.A(_08085_),
    .B(_08247_),
    .Y(_08248_));
 sky130_fd_sc_hd__xnor2_1 _15766_ (.A(_08154_),
    .B(_08182_),
    .Y(_08249_));
 sky130_fd_sc_hd__mux2_1 _15767_ (.A0(_08243_),
    .A1(_08065_),
    .S(_08181_),
    .X(_08250_));
 sky130_fd_sc_hd__nand2_1 _15768_ (.A(_08249_),
    .B(_08250_),
    .Y(_08251_));
 sky130_fd_sc_hd__or2_1 _15769_ (.A(_08249_),
    .B(_08250_),
    .X(_08252_));
 sky130_fd_sc_hd__and2_1 _15770_ (.A(_08251_),
    .B(_08252_),
    .X(_08253_));
 sky130_fd_sc_hd__nand2_1 _15771_ (.A(_08066_),
    .B(_08253_),
    .Y(_08254_));
 sky130_fd_sc_hd__or2_1 _15772_ (.A(_08066_),
    .B(_08253_),
    .X(_08255_));
 sky130_fd_sc_hd__nand2_1 _15773_ (.A(_08254_),
    .B(_08255_),
    .Y(_08256_));
 sky130_fd_sc_hd__a21o_1 _15774_ (.A1(_08245_),
    .A2(_08248_),
    .B1(_08256_),
    .X(_08257_));
 sky130_fd_sc_hd__xor2_1 _15775_ (.A(_08158_),
    .B(_08184_),
    .X(_08258_));
 sky130_fd_sc_hd__a21o_1 _15776_ (.A1(_08251_),
    .A2(_08254_),
    .B1(_08258_),
    .X(_08259_));
 sky130_fd_sc_hd__and2_1 _15777_ (.A(_08257_),
    .B(_08259_),
    .X(_08260_));
 sky130_fd_sc_hd__xnor2_4 _15778_ (.A(_06744_),
    .B(_08221_),
    .Y(_08261_));
 sky130_fd_sc_hd__xor2_4 _15779_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[6] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.sin_17[5] ),
    .X(_08262_));
 sky130_fd_sc_hd__a21boi_4 _15780_ (.A1(_06737_),
    .A2(_08262_),
    .B1_N(_07711_),
    .Y(_08263_));
 sky130_fd_sc_hd__xnor2_1 _15781_ (.A(_08261_),
    .B(_08263_),
    .Y(_08264_));
 sky130_fd_sc_hd__or2_1 _15782_ (.A(_08261_),
    .B(_08263_),
    .X(_08265_));
 sky130_fd_sc_hd__o21a_2 _15783_ (.A1(_08167_),
    .A2(_08264_),
    .B1(_08265_),
    .X(_08266_));
 sky130_fd_sc_hd__xor2_2 _15784_ (.A(_08143_),
    .B(_08223_),
    .X(_08267_));
 sky130_fd_sc_hd__xor2_1 _15785_ (.A(_08266_),
    .B(_08267_),
    .X(_08268_));
 sky130_fd_sc_hd__xnor2_1 _15786_ (.A(_08103_),
    .B(_08142_),
    .Y(_08269_));
 sky130_fd_sc_hd__xnor2_1 _15787_ (.A(_08268_),
    .B(_08269_),
    .Y(_08270_));
 sky130_fd_sc_hd__xnor2_4 _15788_ (.A(_06736_),
    .B(_08262_),
    .Y(_08271_));
 sky130_fd_sc_hd__xor2_4 _15789_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[5] ),
    .B(_06895_),
    .X(_08272_));
 sky130_fd_sc_hd__a21boi_4 _15790_ (.A1(_06738_),
    .A2(_08272_),
    .B1_N(_07740_),
    .Y(_08273_));
 sky130_fd_sc_hd__xnor2_1 _15791_ (.A(_08271_),
    .B(_08273_),
    .Y(_08274_));
 sky130_fd_sc_hd__or2_1 _15792_ (.A(_08271_),
    .B(_08273_),
    .X(_08275_));
 sky130_fd_sc_hd__o21a_1 _15793_ (.A1(_08200_),
    .A2(_08274_),
    .B1(_08275_),
    .X(_08276_));
 sky130_fd_sc_hd__xor2_2 _15794_ (.A(_08167_),
    .B(_08264_),
    .X(_08277_));
 sky130_fd_sc_hd__xnor2_1 _15795_ (.A(_08276_),
    .B(_08277_),
    .Y(_08278_));
 sky130_fd_sc_hd__xnor2_1 _15796_ (.A(_08090_),
    .B(_08166_),
    .Y(_08279_));
 sky130_fd_sc_hd__xor2_1 _15797_ (.A(_08093_),
    .B(_08279_),
    .X(_08280_));
 sky130_fd_sc_hd__and2b_1 _15798_ (.A_N(_08276_),
    .B(_08277_),
    .X(_08281_));
 sky130_fd_sc_hd__a21oi_1 _15799_ (.A1(_08278_),
    .A2(_08280_),
    .B1(_08281_),
    .Y(_08282_));
 sky130_fd_sc_hd__nor2_1 _15800_ (.A(_08270_),
    .B(_08282_),
    .Y(_08283_));
 sky130_fd_sc_hd__nand2_1 _15801_ (.A(_08270_),
    .B(_08282_),
    .Y(_08284_));
 sky130_fd_sc_hd__or2b_1 _15802_ (.A(_08283_),
    .B_N(_08284_),
    .X(_08285_));
 sky130_fd_sc_hd__or2_1 _15803_ (.A(_08090_),
    .B(_08166_),
    .X(_08286_));
 sky130_fd_sc_hd__o21a_1 _15804_ (.A1(_08093_),
    .A2(_08279_),
    .B1(_08286_),
    .X(_08287_));
 sky130_fd_sc_hd__xnor2_1 _15805_ (.A(_06600_),
    .B(_08287_),
    .Y(_08288_));
 sky130_fd_sc_hd__xor2_1 _15806_ (.A(_08130_),
    .B(_08288_),
    .X(_08289_));
 sky130_fd_sc_hd__xnor2_1 _15807_ (.A(_08285_),
    .B(_08289_),
    .Y(_08290_));
 sky130_fd_sc_hd__xnor2_1 _15808_ (.A(_08278_),
    .B(_08280_),
    .Y(_08291_));
 sky130_fd_sc_hd__xor2_2 _15809_ (.A(_08200_),
    .B(_08274_),
    .X(_08292_));
 sky130_fd_sc_hd__xnor2_4 _15810_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[6] ),
    .B(_08272_),
    .Y(_08293_));
 sky130_fd_sc_hd__xor2_4 _15811_ (.A(_06895_),
    .B(\wfg_stim_sine_top.wfg_stim_sine.sin_17[3] ),
    .X(_08294_));
 sky130_fd_sc_hd__a21boi_4 _15812_ (.A1(_06750_),
    .A2(_08294_),
    .B1_N(_07764_),
    .Y(_08295_));
 sky130_fd_sc_hd__xnor2_2 _15813_ (.A(_08293_),
    .B(_08295_),
    .Y(_08296_));
 sky130_fd_sc_hd__or2_1 _15814_ (.A(_08293_),
    .B(_08295_),
    .X(_08297_));
 sky130_fd_sc_hd__o21a_2 _15815_ (.A1(_08220_),
    .A2(_08296_),
    .B1(_08297_),
    .X(_08298_));
 sky130_fd_sc_hd__xnor2_1 _15816_ (.A(_08292_),
    .B(_08298_),
    .Y(_08299_));
 sky130_fd_sc_hd__xnor2_1 _15817_ (.A(_08122_),
    .B(_08202_),
    .Y(_08300_));
 sky130_fd_sc_hd__xor2_1 _15818_ (.A(_08124_),
    .B(_08300_),
    .X(_08301_));
 sky130_fd_sc_hd__and2b_1 _15819_ (.A_N(_08298_),
    .B(_08292_),
    .X(_08302_));
 sky130_fd_sc_hd__a21oi_1 _15820_ (.A1(_08299_),
    .A2(_08301_),
    .B1(_08302_),
    .Y(_08303_));
 sky130_fd_sc_hd__or2_1 _15821_ (.A(_08291_),
    .B(_08303_),
    .X(_08304_));
 sky130_fd_sc_hd__nand2_1 _15822_ (.A(_08291_),
    .B(_08303_),
    .Y(_08305_));
 sky130_fd_sc_hd__nand2_1 _15823_ (.A(_08304_),
    .B(_08305_),
    .Y(_08306_));
 sky130_fd_sc_hd__o31a_1 _15824_ (.A1(_06513_),
    .A2(_08109_),
    .A3(_08110_),
    .B1(_08112_),
    .X(_08307_));
 sky130_fd_sc_hd__nor2_1 _15825_ (.A(_08122_),
    .B(_08202_),
    .Y(_08308_));
 sky130_fd_sc_hd__nor2_1 _15826_ (.A(_08124_),
    .B(_08300_),
    .Y(_08309_));
 sky130_fd_sc_hd__a21bo_1 _15827_ (.A1(_06525_),
    .A2(_06454_),
    .B1_N(_06510_),
    .X(_08310_));
 sky130_fd_sc_hd__o21a_1 _15828_ (.A1(_06525_),
    .A2(_06454_),
    .B1(_08310_),
    .X(_08311_));
 sky130_fd_sc_hd__o21a_1 _15829_ (.A1(_08308_),
    .A2(_08309_),
    .B1(_08311_),
    .X(_08312_));
 sky130_fd_sc_hd__nor3_1 _15830_ (.A(_08311_),
    .B(_08308_),
    .C(_08309_),
    .Y(_08313_));
 sky130_fd_sc_hd__nor2_1 _15831_ (.A(_08312_),
    .B(_08313_),
    .Y(_08314_));
 sky130_fd_sc_hd__xnor2_1 _15832_ (.A(_08307_),
    .B(_08314_),
    .Y(_08315_));
 sky130_fd_sc_hd__o21a_1 _15833_ (.A1(_08306_),
    .A2(_08315_),
    .B1(_08304_),
    .X(_08316_));
 sky130_fd_sc_hd__xor2_1 _15834_ (.A(_08290_),
    .B(_08316_),
    .X(_08317_));
 sky130_fd_sc_hd__a21oi_1 _15835_ (.A1(_08307_),
    .A2(_08314_),
    .B1(_08312_),
    .Y(_08318_));
 sky130_fd_sc_hd__xnor2_1 _15836_ (.A(_08317_),
    .B(_08318_),
    .Y(_08319_));
 sky130_fd_sc_hd__xor2_1 _15837_ (.A(_08306_),
    .B(_08315_),
    .X(_08320_));
 sky130_fd_sc_hd__xnor2_1 _15838_ (.A(_08299_),
    .B(_08301_),
    .Y(_08321_));
 sky130_fd_sc_hd__xor2_4 _15839_ (.A(_08220_),
    .B(_08296_),
    .X(_08322_));
 sky130_fd_sc_hd__xnor2_4 _15840_ (.A(_06750_),
    .B(_08294_),
    .Y(_08323_));
 sky130_fd_sc_hd__xor2_4 _15841_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[3] ),
    .B(_06970_),
    .X(_08324_));
 sky130_fd_sc_hd__a21oi_4 _15842_ (.A1(_06965_),
    .A2(_08324_),
    .B1(_07800_),
    .Y(_08325_));
 sky130_fd_sc_hd__and2_1 _15843_ (.A(_08323_),
    .B(_08325_),
    .X(_08326_));
 sky130_fd_sc_hd__or2_1 _15844_ (.A(_08323_),
    .B(_08325_),
    .X(_08327_));
 sky130_fd_sc_hd__o21a_2 _15845_ (.A1(_08261_),
    .A2(_08326_),
    .B1(_08327_),
    .X(_08328_));
 sky130_fd_sc_hd__xnor2_1 _15846_ (.A(_08322_),
    .B(_08328_),
    .Y(_08329_));
 sky130_fd_sc_hd__clkinv_2 _15847_ (.A(_08142_),
    .Y(_08330_));
 sky130_fd_sc_hd__nand2_1 _15848_ (.A(_08143_),
    .B(_08222_),
    .Y(_08331_));
 sky130_fd_sc_hd__or2_1 _15849_ (.A(_08143_),
    .B(_08222_),
    .X(_08332_));
 sky130_fd_sc_hd__nand2_1 _15850_ (.A(_08331_),
    .B(_08332_),
    .Y(_08333_));
 sky130_fd_sc_hd__xnor2_1 _15851_ (.A(_08330_),
    .B(_08333_),
    .Y(_08334_));
 sky130_fd_sc_hd__and2b_1 _15852_ (.A_N(_08328_),
    .B(_08322_),
    .X(_08335_));
 sky130_fd_sc_hd__a21oi_1 _15853_ (.A1(_08329_),
    .A2(_08334_),
    .B1(_08335_),
    .Y(_08336_));
 sky130_fd_sc_hd__xnor2_1 _15854_ (.A(_08321_),
    .B(_08336_),
    .Y(_08337_));
 sky130_fd_sc_hd__a21oi_2 _15855_ (.A1(_06463_),
    .A2(_08129_),
    .B1(_08110_),
    .Y(_08338_));
 sky130_fd_sc_hd__o21ai_1 _15856_ (.A1(_08142_),
    .A2(_08333_),
    .B1(_08332_),
    .Y(_08339_));
 sky130_fd_sc_hd__xnor2_1 _15857_ (.A(_08338_),
    .B(_08339_),
    .Y(_08340_));
 sky130_fd_sc_hd__xnor2_1 _15858_ (.A(_08106_),
    .B(_08340_),
    .Y(_08341_));
 sky130_fd_sc_hd__or2_1 _15859_ (.A(_08337_),
    .B(_08341_),
    .X(_08342_));
 sky130_fd_sc_hd__o21a_1 _15860_ (.A1(_08321_),
    .A2(_08336_),
    .B1(_08342_),
    .X(_08343_));
 sky130_fd_sc_hd__xnor2_1 _15861_ (.A(_08320_),
    .B(_08343_),
    .Y(_08344_));
 sky130_fd_sc_hd__nand2_1 _15862_ (.A(_08338_),
    .B(_08339_),
    .Y(_08345_));
 sky130_fd_sc_hd__o21a_1 _15863_ (.A1(_08106_),
    .A2(_08340_),
    .B1(_08345_),
    .X(_08346_));
 sky130_fd_sc_hd__inv_2 _15864_ (.A(_08346_),
    .Y(_08347_));
 sky130_fd_sc_hd__and2b_1 _15865_ (.A_N(_08343_),
    .B(_08320_),
    .X(_08348_));
 sky130_fd_sc_hd__a21o_1 _15866_ (.A1(_08344_),
    .A2(_08347_),
    .B1(_08348_),
    .X(_08349_));
 sky130_fd_sc_hd__xnor2_1 _15867_ (.A(_08319_),
    .B(_08349_),
    .Y(_08350_));
 sky130_fd_sc_hd__nand2_1 _15868_ (.A(_08065_),
    .B(_08350_),
    .Y(_08351_));
 sky130_fd_sc_hd__or2_1 _15869_ (.A(_08065_),
    .B(_08350_),
    .X(_08352_));
 sky130_fd_sc_hd__nand2_1 _15870_ (.A(_08351_),
    .B(_08352_),
    .Y(_08353_));
 sky130_fd_sc_hd__xnor2_1 _15871_ (.A(_08329_),
    .B(_08334_),
    .Y(_08354_));
 sky130_fd_sc_hd__xor2_1 _15872_ (.A(_08323_),
    .B(_08325_),
    .X(_08355_));
 sky130_fd_sc_hd__xnor2_2 _15873_ (.A(_08261_),
    .B(_08355_),
    .Y(_08356_));
 sky130_fd_sc_hd__inv_2 _15874_ (.A(_08271_),
    .Y(_08357_));
 sky130_fd_sc_hd__xor2_4 _15875_ (.A(_06970_),
    .B(\wfg_stim_sine_top.wfg_stim_sine.sin_17[1] ),
    .X(_08358_));
 sky130_fd_sc_hd__a21oi_4 _15876_ (.A1(_06995_),
    .A2(_08358_),
    .B1(_07812_),
    .Y(_08359_));
 sky130_fd_sc_hd__xnor2_4 _15877_ (.A(_06895_),
    .B(_08324_),
    .Y(_08360_));
 sky130_fd_sc_hd__xor2_4 _15878_ (.A(_08359_),
    .B(_08360_),
    .X(_08361_));
 sky130_fd_sc_hd__nor2_2 _15879_ (.A(_08359_),
    .B(_08360_),
    .Y(_08362_));
 sky130_fd_sc_hd__a21oi_2 _15880_ (.A1(_08357_),
    .A2(_08361_),
    .B1(_08362_),
    .Y(_08363_));
 sky130_fd_sc_hd__xnor2_4 _15881_ (.A(_08356_),
    .B(_08363_),
    .Y(_08364_));
 sky130_fd_sc_hd__inv_2 _15882_ (.A(_08166_),
    .Y(_08365_));
 sky130_fd_sc_hd__nand2_1 _15883_ (.A(_08167_),
    .B(_08263_),
    .Y(_08366_));
 sky130_fd_sc_hd__or2_1 _15884_ (.A(_08167_),
    .B(_08263_),
    .X(_08367_));
 sky130_fd_sc_hd__nand2_1 _15885_ (.A(_08366_),
    .B(_08367_),
    .Y(_08368_));
 sky130_fd_sc_hd__xnor2_1 _15886_ (.A(_08365_),
    .B(_08368_),
    .Y(_08369_));
 sky130_fd_sc_hd__or2b_1 _15887_ (.A(_08363_),
    .B_N(_08356_),
    .X(_08370_));
 sky130_fd_sc_hd__a21boi_2 _15888_ (.A1(_08364_),
    .A2(_08369_),
    .B1_N(_08370_),
    .Y(_08371_));
 sky130_fd_sc_hd__nand2_1 _15889_ (.A(_08354_),
    .B(_08371_),
    .Y(_08372_));
 sky130_fd_sc_hd__o21a_1 _15890_ (.A1(_08166_),
    .A2(_08368_),
    .B1(_08367_),
    .X(_08373_));
 sky130_fd_sc_hd__xnor2_1 _15891_ (.A(_08134_),
    .B(_08373_),
    .Y(_08374_));
 sky130_fd_sc_hd__xor2_2 _15892_ (.A(_08096_),
    .B(_08374_),
    .X(_08375_));
 sky130_fd_sc_hd__nor2_1 _15893_ (.A(_08354_),
    .B(_08371_),
    .Y(_08376_));
 sky130_fd_sc_hd__a21oi_2 _15894_ (.A1(_08372_),
    .A2(_08375_),
    .B1(_08376_),
    .Y(_08377_));
 sky130_fd_sc_hd__xor2_1 _15895_ (.A(_08337_),
    .B(_08341_),
    .X(_08378_));
 sky130_fd_sc_hd__or2b_1 _15896_ (.A(_08377_),
    .B_N(_08378_),
    .X(_08379_));
 sky130_fd_sc_hd__or2_1 _15897_ (.A(_08096_),
    .B(_08374_),
    .X(_08380_));
 sky130_fd_sc_hd__o21a_2 _15898_ (.A1(_08134_),
    .A2(_08373_),
    .B1(_08380_),
    .X(_08381_));
 sky130_fd_sc_hd__xnor2_2 _15899_ (.A(_08378_),
    .B(_08377_),
    .Y(_08382_));
 sky130_fd_sc_hd__or2b_1 _15900_ (.A(_08381_),
    .B_N(_08382_),
    .X(_08383_));
 sky130_fd_sc_hd__xnor2_1 _15901_ (.A(_08344_),
    .B(_08347_),
    .Y(_08384_));
 sky130_fd_sc_hd__a21o_1 _15902_ (.A1(_08379_),
    .A2(_08383_),
    .B1(_08384_),
    .X(_08385_));
 sky130_fd_sc_hd__nand3_1 _15903_ (.A(_08384_),
    .B(_08379_),
    .C(_08383_),
    .Y(_08386_));
 sky130_fd_sc_hd__and2_1 _15904_ (.A(_08385_),
    .B(_08386_),
    .X(_08387_));
 sky130_fd_sc_hd__nand2_1 _15905_ (.A(_08065_),
    .B(_08387_),
    .Y(_08388_));
 sky130_fd_sc_hd__nand3_1 _15906_ (.A(_08353_),
    .B(_08385_),
    .C(_08388_),
    .Y(_08389_));
 sky130_fd_sc_hd__inv_2 _15907_ (.A(_08389_),
    .Y(_08390_));
 sky130_fd_sc_hd__a21oi_1 _15908_ (.A1(_08385_),
    .A2(_08388_),
    .B1(_08353_),
    .Y(_08391_));
 sky130_fd_sc_hd__nor2_1 _15909_ (.A(_08390_),
    .B(_08391_),
    .Y(_08392_));
 sky130_fd_sc_hd__xnor2_4 _15910_ (.A(_08382_),
    .B(_08381_),
    .Y(_08393_));
 sky130_fd_sc_hd__xnor2_1 _15911_ (.A(_08354_),
    .B(_08371_),
    .Y(_08394_));
 sky130_fd_sc_hd__xnor2_1 _15912_ (.A(_08394_),
    .B(_08375_),
    .Y(_08395_));
 sky130_fd_sc_hd__xnor2_1 _15913_ (.A(_08364_),
    .B(_08369_),
    .Y(_08396_));
 sky130_fd_sc_hd__xnor2_2 _15914_ (.A(_08271_),
    .B(_08361_),
    .Y(_08397_));
 sky130_fd_sc_hd__inv_2 _15915_ (.A(_08293_),
    .Y(_08398_));
 sky130_fd_sc_hd__xor2_4 _15916_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[1] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.sin_17[0] ),
    .X(_08399_));
 sky130_fd_sc_hd__and2_2 _15917_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[1] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.sin_17[0] ),
    .X(_08400_));
 sky130_fd_sc_hd__a21oi_4 _15918_ (.A1(_06991_),
    .A2(_08399_),
    .B1(_08400_),
    .Y(_08401_));
 sky130_fd_sc_hd__xnor2_4 _15919_ (.A(_06995_),
    .B(_08358_),
    .Y(_08402_));
 sky130_fd_sc_hd__xor2_2 _15920_ (.A(_08401_),
    .B(_08402_),
    .X(_08403_));
 sky130_fd_sc_hd__nor2_2 _15921_ (.A(_08401_),
    .B(_08402_),
    .Y(_08404_));
 sky130_fd_sc_hd__a21oi_2 _15922_ (.A1(_08398_),
    .A2(_08403_),
    .B1(_08404_),
    .Y(_08405_));
 sky130_fd_sc_hd__xnor2_4 _15923_ (.A(_08397_),
    .B(_08405_),
    .Y(_08406_));
 sky130_fd_sc_hd__inv_2 _15924_ (.A(_08202_),
    .Y(_08407_));
 sky130_fd_sc_hd__nand2_1 _15925_ (.A(_08200_),
    .B(_08273_),
    .Y(_08408_));
 sky130_fd_sc_hd__or2_1 _15926_ (.A(_08200_),
    .B(_08273_),
    .X(_08409_));
 sky130_fd_sc_hd__nand2_1 _15927_ (.A(_08408_),
    .B(_08409_),
    .Y(_08410_));
 sky130_fd_sc_hd__xnor2_2 _15928_ (.A(_08407_),
    .B(_08410_),
    .Y(_08411_));
 sky130_fd_sc_hd__or2b_1 _15929_ (.A(_08405_),
    .B_N(_08397_),
    .X(_08412_));
 sky130_fd_sc_hd__a21boi_2 _15930_ (.A1(_08406_),
    .A2(_08411_),
    .B1_N(_08412_),
    .Y(_08413_));
 sky130_fd_sc_hd__nand2_1 _15931_ (.A(_08396_),
    .B(_08413_),
    .Y(_08414_));
 sky130_fd_sc_hd__o21a_1 _15932_ (.A1(_08202_),
    .A2(_08410_),
    .B1(_08409_),
    .X(_08415_));
 sky130_fd_sc_hd__xnor2_2 _15933_ (.A(_08119_),
    .B(_08415_),
    .Y(_08416_));
 sky130_fd_sc_hd__xor2_2 _15934_ (.A(_08127_),
    .B(_08416_),
    .X(_08417_));
 sky130_fd_sc_hd__nor2_1 _15935_ (.A(_08396_),
    .B(_08413_),
    .Y(_08418_));
 sky130_fd_sc_hd__a21oi_2 _15936_ (.A1(_08414_),
    .A2(_08417_),
    .B1(_08418_),
    .Y(_08419_));
 sky130_fd_sc_hd__xnor2_2 _15937_ (.A(_08395_),
    .B(_08419_),
    .Y(_08420_));
 sky130_fd_sc_hd__or2_1 _15938_ (.A(_08119_),
    .B(_08415_),
    .X(_08421_));
 sky130_fd_sc_hd__o21ai_2 _15939_ (.A1(_08127_),
    .A2(_08416_),
    .B1(_08421_),
    .Y(_08422_));
 sky130_fd_sc_hd__and2b_1 _15940_ (.A_N(_08419_),
    .B(_08395_),
    .X(_08423_));
 sky130_fd_sc_hd__a21o_1 _15941_ (.A1(_08420_),
    .A2(_08422_),
    .B1(_08423_),
    .X(_08424_));
 sky130_fd_sc_hd__xor2_4 _15942_ (.A(_08393_),
    .B(_08424_),
    .X(_08425_));
 sky130_fd_sc_hd__xnor2_2 _15943_ (.A(_06600_),
    .B(_08425_),
    .Y(_08426_));
 sky130_fd_sc_hd__xnor2_2 _15944_ (.A(_08420_),
    .B(_08422_),
    .Y(_08427_));
 sky130_fd_sc_hd__xnor2_1 _15945_ (.A(_08396_),
    .B(_08413_),
    .Y(_08428_));
 sky130_fd_sc_hd__xnor2_2 _15946_ (.A(_08428_),
    .B(_08417_),
    .Y(_08429_));
 sky130_fd_sc_hd__xnor2_2 _15947_ (.A(_08406_),
    .B(_08411_),
    .Y(_08430_));
 sky130_fd_sc_hd__xnor2_1 _15948_ (.A(_08293_),
    .B(_08403_),
    .Y(_08431_));
 sky130_fd_sc_hd__inv_2 _15949_ (.A(_08323_),
    .Y(_08432_));
 sky130_fd_sc_hd__xnor2_4 _15950_ (.A(_06970_),
    .B(_08399_),
    .Y(_08433_));
 sky130_fd_sc_hd__xnor2_4 _15951_ (.A(_08400_),
    .B(_08433_),
    .Y(_08434_));
 sky130_fd_sc_hd__nor2_1 _15952_ (.A(_07001_),
    .B(_08433_),
    .Y(_08435_));
 sky130_fd_sc_hd__a21oi_1 _15953_ (.A1(_08432_),
    .A2(_08434_),
    .B1(_08435_),
    .Y(_08436_));
 sky130_fd_sc_hd__xnor2_2 _15954_ (.A(_08431_),
    .B(_08436_),
    .Y(_08437_));
 sky130_fd_sc_hd__nand2_1 _15955_ (.A(_08220_),
    .B(_08295_),
    .Y(_08438_));
 sky130_fd_sc_hd__or2_1 _15956_ (.A(_08220_),
    .B(_08295_),
    .X(_08439_));
 sky130_fd_sc_hd__nand2_1 _15957_ (.A(_08438_),
    .B(_08439_),
    .Y(_08440_));
 sky130_fd_sc_hd__xor2_1 _15958_ (.A(_08222_),
    .B(_08440_),
    .X(_08441_));
 sky130_fd_sc_hd__and2b_1 _15959_ (.A_N(_08436_),
    .B(_08431_),
    .X(_08442_));
 sky130_fd_sc_hd__a21oi_2 _15960_ (.A1(_08437_),
    .A2(_08441_),
    .B1(_08442_),
    .Y(_08443_));
 sky130_fd_sc_hd__nand2_1 _15961_ (.A(_08430_),
    .B(_08443_),
    .Y(_08444_));
 sky130_fd_sc_hd__o21a_1 _15962_ (.A1(_08222_),
    .A2(_08440_),
    .B1(_08439_),
    .X(_08445_));
 sky130_fd_sc_hd__xnor2_1 _15963_ (.A(_08147_),
    .B(_08445_),
    .Y(_08446_));
 sky130_fd_sc_hd__xor2_1 _15964_ (.A(_08146_),
    .B(_08446_),
    .X(_08447_));
 sky130_fd_sc_hd__nor2_1 _15965_ (.A(_08430_),
    .B(_08443_),
    .Y(_08448_));
 sky130_fd_sc_hd__a21oi_1 _15966_ (.A1(_08444_),
    .A2(_08447_),
    .B1(_08448_),
    .Y(_08449_));
 sky130_fd_sc_hd__xnor2_2 _15967_ (.A(_08429_),
    .B(_08449_),
    .Y(_08450_));
 sky130_fd_sc_hd__and2b_1 _15968_ (.A_N(_08445_),
    .B(_08147_),
    .X(_08451_));
 sky130_fd_sc_hd__a21o_1 _15969_ (.A1(_08146_),
    .A2(_08446_),
    .B1(_08451_),
    .X(_08452_));
 sky130_fd_sc_hd__or2b_1 _15970_ (.A(_08449_),
    .B_N(_08429_),
    .X(_08453_));
 sky130_fd_sc_hd__a21bo_1 _15971_ (.A1(_08450_),
    .A2(_08452_),
    .B1_N(_08453_),
    .X(_08454_));
 sky130_fd_sc_hd__xnor2_2 _15972_ (.A(_08427_),
    .B(_08454_),
    .Y(_08455_));
 sky130_fd_sc_hd__or2b_1 _15973_ (.A(_08427_),
    .B_N(_08454_),
    .X(_08456_));
 sky130_fd_sc_hd__a21boi_2 _15974_ (.A1(_06600_),
    .A2(_08455_),
    .B1_N(_08456_),
    .Y(_08457_));
 sky130_fd_sc_hd__nand2_1 _15975_ (.A(_08426_),
    .B(_08457_),
    .Y(_08458_));
 sky130_fd_sc_hd__xnor2_1 _15976_ (.A(_06600_),
    .B(_08455_),
    .Y(_08459_));
 sky130_fd_sc_hd__xnor2_2 _15977_ (.A(_08450_),
    .B(_08452_),
    .Y(_08460_));
 sky130_fd_sc_hd__xnor2_1 _15978_ (.A(_08430_),
    .B(_08443_),
    .Y(_08461_));
 sky130_fd_sc_hd__xnor2_1 _15979_ (.A(_08461_),
    .B(_08447_),
    .Y(_08462_));
 sky130_fd_sc_hd__xnor2_1 _15980_ (.A(_08437_),
    .B(_08441_),
    .Y(_08463_));
 sky130_fd_sc_hd__xnor2_2 _15981_ (.A(_08323_),
    .B(_08434_),
    .Y(_08464_));
 sky130_fd_sc_hd__and2b_1 _15982_ (.A_N(_08360_),
    .B(_08399_),
    .X(_08465_));
 sky130_fd_sc_hd__nand2_2 _15983_ (.A(_08464_),
    .B(_08465_),
    .Y(_08466_));
 sky130_fd_sc_hd__xnor2_1 _15984_ (.A(_08464_),
    .B(_08465_),
    .Y(_08467_));
 sky130_fd_sc_hd__xnor2_1 _15985_ (.A(_08261_),
    .B(_08325_),
    .Y(_08468_));
 sky130_fd_sc_hd__nor2_1 _15986_ (.A(_08263_),
    .B(_08468_),
    .Y(_08469_));
 sky130_fd_sc_hd__and2_1 _15987_ (.A(_08263_),
    .B(_08468_),
    .X(_08470_));
 sky130_fd_sc_hd__or2_1 _15988_ (.A(_08469_),
    .B(_08470_),
    .X(_08471_));
 sky130_fd_sc_hd__or2_1 _15989_ (.A(_08467_),
    .B(_08471_),
    .X(_08472_));
 sky130_fd_sc_hd__nand3_1 _15990_ (.A(_08463_),
    .B(_08466_),
    .C(_08472_),
    .Y(_08473_));
 sky130_fd_sc_hd__nor2_1 _15991_ (.A(_08261_),
    .B(_08325_),
    .Y(_08474_));
 sky130_fd_sc_hd__o21a_1 _15992_ (.A1(_08474_),
    .A2(_08469_),
    .B1(_08172_),
    .X(_08475_));
 sky130_fd_sc_hd__or3_1 _15993_ (.A(_08172_),
    .B(_08474_),
    .C(_08469_),
    .X(_08476_));
 sky130_fd_sc_hd__and2b_1 _15994_ (.A_N(_08475_),
    .B(_08476_),
    .X(_08477_));
 sky130_fd_sc_hd__xnor2_2 _15995_ (.A(_08175_),
    .B(_08477_),
    .Y(_08478_));
 sky130_fd_sc_hd__a21oi_1 _15996_ (.A1(_08466_),
    .A2(_08472_),
    .B1(_08463_),
    .Y(_08479_));
 sky130_fd_sc_hd__a21oi_1 _15997_ (.A1(_08473_),
    .A2(_08478_),
    .B1(_08479_),
    .Y(_08480_));
 sky130_fd_sc_hd__xnor2_1 _15998_ (.A(_08462_),
    .B(_08480_),
    .Y(_08481_));
 sky130_fd_sc_hd__a21o_1 _15999_ (.A1(_08171_),
    .A2(_08476_),
    .B1(_08475_),
    .X(_08482_));
 sky130_fd_sc_hd__or2b_1 _16000_ (.A(_08480_),
    .B_N(_08462_),
    .X(_08483_));
 sky130_fd_sc_hd__a21bo_1 _16001_ (.A1(_08481_),
    .A2(_08482_),
    .B1_N(_08483_),
    .X(_08484_));
 sky130_fd_sc_hd__xnor2_1 _16002_ (.A(_08460_),
    .B(_08484_),
    .Y(_08485_));
 sky130_fd_sc_hd__or2b_1 _16003_ (.A(_08460_),
    .B_N(_08484_),
    .X(_08486_));
 sky130_fd_sc_hd__a21boi_1 _16004_ (.A1(_08130_),
    .A2(_08485_),
    .B1_N(_08486_),
    .Y(_08487_));
 sky130_fd_sc_hd__nor2_1 _16005_ (.A(_08459_),
    .B(_08487_),
    .Y(_08488_));
 sky130_fd_sc_hd__nor2_1 _16006_ (.A(_08426_),
    .B(_08457_),
    .Y(_08489_));
 sky130_fd_sc_hd__a21o_1 _16007_ (.A1(_08458_),
    .A2(_08488_),
    .B1(_08489_),
    .X(_08490_));
 sky130_fd_sc_hd__xnor2_1 _16008_ (.A(_08481_),
    .B(_08482_),
    .Y(_08491_));
 sky130_fd_sc_hd__or2b_1 _16009_ (.A(_08479_),
    .B_N(_08473_),
    .X(_08492_));
 sky130_fd_sc_hd__xnor2_1 _16010_ (.A(_08492_),
    .B(_08478_),
    .Y(_08493_));
 sky130_fd_sc_hd__xor2_1 _16011_ (.A(_08467_),
    .B(_08471_),
    .X(_08494_));
 sky130_fd_sc_hd__inv_2 _16012_ (.A(\wfg_stim_sine_top.wfg_stim_sine.sin_17[0] ),
    .Y(_08495_));
 sky130_fd_sc_hd__or2_1 _16013_ (.A(_08495_),
    .B(_08402_),
    .X(_08496_));
 sky130_fd_sc_hd__xnor2_1 _16014_ (.A(_08360_),
    .B(_08399_),
    .Y(_08497_));
 sky130_fd_sc_hd__xnor2_1 _16015_ (.A(_08496_),
    .B(_08497_),
    .Y(_08498_));
 sky130_fd_sc_hd__xnor2_1 _16016_ (.A(_08271_),
    .B(_08359_),
    .Y(_08499_));
 sky130_fd_sc_hd__xor2_1 _16017_ (.A(_08273_),
    .B(_08499_),
    .X(_08500_));
 sky130_fd_sc_hd__and2b_1 _16018_ (.A_N(_08496_),
    .B(_08497_),
    .X(_08501_));
 sky130_fd_sc_hd__a21oi_1 _16019_ (.A1(_08498_),
    .A2(_08500_),
    .B1(_08501_),
    .Y(_08502_));
 sky130_fd_sc_hd__xnor2_1 _16020_ (.A(_08494_),
    .B(_08502_),
    .Y(_08503_));
 sky130_fd_sc_hd__nor2_1 _16021_ (.A(_08271_),
    .B(_08359_),
    .Y(_08504_));
 sky130_fd_sc_hd__nor2_1 _16022_ (.A(_08273_),
    .B(_08499_),
    .Y(_08505_));
 sky130_fd_sc_hd__o21a_1 _16023_ (.A1(_08504_),
    .A2(_08505_),
    .B1(_08207_),
    .X(_08506_));
 sky130_fd_sc_hd__nor3_1 _16024_ (.A(_08207_),
    .B(_08504_),
    .C(_08505_),
    .Y(_08507_));
 sky130_fd_sc_hd__nor2_1 _16025_ (.A(_08506_),
    .B(_08507_),
    .Y(_08508_));
 sky130_fd_sc_hd__xnor2_1 _16026_ (.A(_08206_),
    .B(_08508_),
    .Y(_08509_));
 sky130_fd_sc_hd__and2b_1 _16027_ (.A_N(_08502_),
    .B(_08494_),
    .X(_08510_));
 sky130_fd_sc_hd__a21o_1 _16028_ (.A1(_08503_),
    .A2(_08509_),
    .B1(_08510_),
    .X(_08511_));
 sky130_fd_sc_hd__xor2_1 _16029_ (.A(_08493_),
    .B(_08511_),
    .X(_08512_));
 sky130_fd_sc_hd__a21o_1 _16030_ (.A1(_08213_),
    .A2(_08508_),
    .B1(_08506_),
    .X(_08513_));
 sky130_fd_sc_hd__and2_1 _16031_ (.A(_08493_),
    .B(_08511_),
    .X(_08514_));
 sky130_fd_sc_hd__a21o_1 _16032_ (.A1(_08512_),
    .A2(_08513_),
    .B1(_08514_),
    .X(_08515_));
 sky130_fd_sc_hd__or2b_1 _16033_ (.A(_08491_),
    .B_N(_08515_),
    .X(_08516_));
 sky130_fd_sc_hd__xnor2_1 _16034_ (.A(_08491_),
    .B(_08515_),
    .Y(_08517_));
 sky130_fd_sc_hd__nand2_1 _16035_ (.A(_08108_),
    .B(_08517_),
    .Y(_08518_));
 sky130_fd_sc_hd__xnor2_1 _16036_ (.A(_08130_),
    .B(_08485_),
    .Y(_08519_));
 sky130_fd_sc_hd__a21oi_1 _16037_ (.A1(_08516_),
    .A2(_08518_),
    .B1(_08519_),
    .Y(_08520_));
 sky130_fd_sc_hd__xnor2_1 _16038_ (.A(_08108_),
    .B(_08517_),
    .Y(_08521_));
 sky130_fd_sc_hd__xor2_1 _16039_ (.A(_08512_),
    .B(_08513_),
    .X(_08522_));
 sky130_fd_sc_hd__xnor2_1 _16040_ (.A(_08503_),
    .B(_08509_),
    .Y(_08523_));
 sky130_fd_sc_hd__xnor2_1 _16041_ (.A(_08498_),
    .B(_08500_),
    .Y(_08524_));
 sky130_fd_sc_hd__xnor2_1 _16042_ (.A(_08293_),
    .B(_08401_),
    .Y(_08525_));
 sky130_fd_sc_hd__xnor2_1 _16043_ (.A(_08295_),
    .B(_08525_),
    .Y(_08526_));
 sky130_fd_sc_hd__nand2_1 _16044_ (.A(_08495_),
    .B(_08402_),
    .Y(_08527_));
 sky130_fd_sc_hd__nand2_1 _16045_ (.A(_08496_),
    .B(_08527_),
    .Y(_08528_));
 sky130_fd_sc_hd__or2_2 _16046_ (.A(_08526_),
    .B(_08528_),
    .X(_08529_));
 sky130_fd_sc_hd__or2_1 _16047_ (.A(_08293_),
    .B(_08401_),
    .X(_08530_));
 sky130_fd_sc_hd__o21a_1 _16048_ (.A1(_08295_),
    .A2(_08525_),
    .B1(_08530_),
    .X(_08531_));
 sky130_fd_sc_hd__xnor2_1 _16049_ (.A(_08226_),
    .B(_08531_),
    .Y(_08532_));
 sky130_fd_sc_hd__xor2_1 _16050_ (.A(_08225_),
    .B(_08532_),
    .X(_08533_));
 sky130_fd_sc_hd__xor2_1 _16051_ (.A(_08524_),
    .B(_08529_),
    .X(_08534_));
 sky130_fd_sc_hd__nand2_1 _16052_ (.A(_08533_),
    .B(_08534_),
    .Y(_08535_));
 sky130_fd_sc_hd__o21ai_1 _16053_ (.A1(_08524_),
    .A2(_08529_),
    .B1(_08535_),
    .Y(_08536_));
 sky130_fd_sc_hd__xor2_1 _16054_ (.A(_08523_),
    .B(_08536_),
    .X(_08537_));
 sky130_fd_sc_hd__or2b_1 _16055_ (.A(_08531_),
    .B_N(_08226_),
    .X(_08538_));
 sky130_fd_sc_hd__a21boi_1 _16056_ (.A1(_08225_),
    .A2(_08532_),
    .B1_N(_08538_),
    .Y(_08539_));
 sky130_fd_sc_hd__and2b_1 _16057_ (.A_N(_08523_),
    .B(_08536_),
    .X(_08540_));
 sky130_fd_sc_hd__o21ba_1 _16058_ (.A1(_08537_),
    .A2(_08539_),
    .B1_N(_08540_),
    .X(_08541_));
 sky130_fd_sc_hd__xnor2_1 _16059_ (.A(_08522_),
    .B(_08541_),
    .Y(_08542_));
 sky130_fd_sc_hd__or2b_1 _16060_ (.A(_08541_),
    .B_N(_08522_),
    .X(_08543_));
 sky130_fd_sc_hd__a21bo_1 _16061_ (.A1(_08174_),
    .A2(_08542_),
    .B1_N(_08543_),
    .X(_08544_));
 sky130_fd_sc_hd__and2b_1 _16062_ (.A_N(_08521_),
    .B(_08544_),
    .X(_08545_));
 sky130_fd_sc_hd__xor2_1 _16063_ (.A(_08459_),
    .B(_08487_),
    .X(_08546_));
 sky130_fd_sc_hd__xor2_2 _16064_ (.A(_08426_),
    .B(_08457_),
    .X(_08547_));
 sky130_fd_sc_hd__and2_1 _16065_ (.A(_08546_),
    .B(_08547_),
    .X(_08548_));
 sky130_fd_sc_hd__nand3_1 _16066_ (.A(_08519_),
    .B(_08516_),
    .C(_08518_),
    .Y(_08549_));
 sky130_fd_sc_hd__o211a_1 _16067_ (.A1(_08520_),
    .A2(_08545_),
    .B1(_08548_),
    .C1(_08549_),
    .X(_08550_));
 sky130_fd_sc_hd__xnor2_1 _16068_ (.A(_08537_),
    .B(_08539_),
    .Y(_08551_));
 sky130_fd_sc_hd__xnor2_1 _16069_ (.A(_08533_),
    .B(_08534_),
    .Y(_08552_));
 sky130_fd_sc_hd__nand2_1 _16070_ (.A(_08526_),
    .B(_08528_),
    .Y(_08553_));
 sky130_fd_sc_hd__xnor2_1 _16071_ (.A(_07001_),
    .B(_08323_),
    .Y(_08554_));
 sky130_fd_sc_hd__xnor2_1 _16072_ (.A(_08325_),
    .B(_08554_),
    .Y(_08555_));
 sky130_fd_sc_hd__nor2_2 _16073_ (.A(_08433_),
    .B(_08555_),
    .Y(_08556_));
 sky130_fd_sc_hd__or2_1 _16074_ (.A(_07001_),
    .B(_08323_),
    .X(_08557_));
 sky130_fd_sc_hd__o21a_1 _16075_ (.A1(_08325_),
    .A2(_08554_),
    .B1(_08557_),
    .X(_08558_));
 sky130_fd_sc_hd__xnor2_1 _16076_ (.A(_08267_),
    .B(_08558_),
    .Y(_08559_));
 sky130_fd_sc_hd__xnor2_2 _16077_ (.A(_08266_),
    .B(_08559_),
    .Y(_08560_));
 sky130_fd_sc_hd__xnor2_1 _16078_ (.A(_08526_),
    .B(_08528_),
    .Y(_08561_));
 sky130_fd_sc_hd__xnor2_2 _16079_ (.A(_08561_),
    .B(_08556_),
    .Y(_08562_));
 sky130_fd_sc_hd__a32oi_4 _16080_ (.A1(_08529_),
    .A2(_08553_),
    .A3(_08556_),
    .B1(_08560_),
    .B2(_08562_),
    .Y(_08563_));
 sky130_fd_sc_hd__xnor2_1 _16081_ (.A(_08552_),
    .B(_08563_),
    .Y(_08564_));
 sky130_fd_sc_hd__or2b_1 _16082_ (.A(_08558_),
    .B_N(_08267_),
    .X(_08565_));
 sky130_fd_sc_hd__or2b_1 _16083_ (.A(_08266_),
    .B_N(_08559_),
    .X(_08566_));
 sky130_fd_sc_hd__nand2_1 _16084_ (.A(_08565_),
    .B(_08566_),
    .Y(_08567_));
 sky130_fd_sc_hd__or2b_1 _16085_ (.A(_08564_),
    .B_N(_08567_),
    .X(_08568_));
 sky130_fd_sc_hd__o21ai_1 _16086_ (.A1(_08552_),
    .A2(_08563_),
    .B1(_08568_),
    .Y(_08569_));
 sky130_fd_sc_hd__and2b_1 _16087_ (.A_N(_08551_),
    .B(_08569_),
    .X(_08570_));
 sky130_fd_sc_hd__xor2_1 _16088_ (.A(_08551_),
    .B(_08569_),
    .X(_08571_));
 sky130_fd_sc_hd__nor2_1 _16089_ (.A(_08093_),
    .B(_08571_),
    .Y(_08572_));
 sky130_fd_sc_hd__xnor2_1 _16090_ (.A(_08100_),
    .B(_08542_),
    .Y(_08573_));
 sky130_fd_sc_hd__o21a_1 _16091_ (.A1(_08570_),
    .A2(_08572_),
    .B1(_08573_),
    .X(_08574_));
 sky130_fd_sc_hd__inv_2 _16092_ (.A(_08574_),
    .Y(_08575_));
 sky130_fd_sc_hd__xor2_1 _16093_ (.A(_08567_),
    .B(_08564_),
    .X(_08576_));
 sky130_fd_sc_hd__xnor2_1 _16094_ (.A(_08277_),
    .B(_08362_),
    .Y(_08577_));
 sky130_fd_sc_hd__nand2_1 _16095_ (.A(_08277_),
    .B(_08362_),
    .Y(_08578_));
 sky130_fd_sc_hd__o21ai_1 _16096_ (.A1(_08276_),
    .A2(_08577_),
    .B1(_08578_),
    .Y(_08579_));
 sky130_fd_sc_hd__xnor2_1 _16097_ (.A(_08560_),
    .B(_08562_),
    .Y(_08580_));
 sky130_fd_sc_hd__xnor2_1 _16098_ (.A(_08276_),
    .B(_08577_),
    .Y(_08581_));
 sky130_fd_sc_hd__xor2_1 _16099_ (.A(_08433_),
    .B(_08555_),
    .X(_08582_));
 sky130_fd_sc_hd__and2_1 _16100_ (.A(_08361_),
    .B(_08399_),
    .X(_08583_));
 sky130_fd_sc_hd__xnor2_1 _16101_ (.A(_08582_),
    .B(_08583_),
    .Y(_08584_));
 sky130_fd_sc_hd__nand2_1 _16102_ (.A(_08582_),
    .B(_08583_),
    .Y(_08585_));
 sky130_fd_sc_hd__o21a_1 _16103_ (.A1(_08581_),
    .A2(_08584_),
    .B1(_08585_),
    .X(_08586_));
 sky130_fd_sc_hd__xor2_1 _16104_ (.A(_08580_),
    .B(_08586_),
    .X(_08587_));
 sky130_fd_sc_hd__nor2_1 _16105_ (.A(_08580_),
    .B(_08586_),
    .Y(_08588_));
 sky130_fd_sc_hd__a21oi_1 _16106_ (.A1(_08579_),
    .A2(_08587_),
    .B1(_08588_),
    .Y(_08589_));
 sky130_fd_sc_hd__or2_1 _16107_ (.A(_08576_),
    .B(_08589_),
    .X(_08590_));
 sky130_fd_sc_hd__nand2_1 _16108_ (.A(_08576_),
    .B(_08589_),
    .Y(_08591_));
 sky130_fd_sc_hd__and2_1 _16109_ (.A(_08590_),
    .B(_08591_),
    .X(_08592_));
 sky130_fd_sc_hd__or2b_1 _16110_ (.A(_08124_),
    .B_N(_08592_),
    .X(_08593_));
 sky130_fd_sc_hd__and2_1 _16111_ (.A(_08093_),
    .B(_08571_),
    .X(_08594_));
 sky130_fd_sc_hd__or2_1 _16112_ (.A(_08572_),
    .B(_08594_),
    .X(_08595_));
 sky130_fd_sc_hd__a21o_1 _16113_ (.A1(_08590_),
    .A2(_08593_),
    .B1(_08595_),
    .X(_08596_));
 sky130_fd_sc_hd__xnor2_1 _16114_ (.A(_08124_),
    .B(_08592_),
    .Y(_08597_));
 sky130_fd_sc_hd__xnor2_1 _16115_ (.A(_08579_),
    .B(_08587_),
    .Y(_08598_));
 sky130_fd_sc_hd__xnor2_1 _16116_ (.A(_08292_),
    .B(_08404_),
    .Y(_08599_));
 sky130_fd_sc_hd__nand2_1 _16117_ (.A(_08292_),
    .B(_08404_),
    .Y(_08600_));
 sky130_fd_sc_hd__o21ai_1 _16118_ (.A1(_08298_),
    .A2(_08599_),
    .B1(_08600_),
    .Y(_08601_));
 sky130_fd_sc_hd__xnor2_1 _16119_ (.A(_08581_),
    .B(_08584_),
    .Y(_08602_));
 sky130_fd_sc_hd__nand2_1 _16120_ (.A(_06989_),
    .B(_08403_),
    .Y(_08603_));
 sky130_fd_sc_hd__xnor2_1 _16121_ (.A(_08361_),
    .B(_08399_),
    .Y(_08604_));
 sky130_fd_sc_hd__nand2_1 _16122_ (.A(_08603_),
    .B(_08604_),
    .Y(_08605_));
 sky130_fd_sc_hd__xor2_1 _16123_ (.A(_08298_),
    .B(_08599_),
    .X(_08606_));
 sky130_fd_sc_hd__nor2_1 _16124_ (.A(_08603_),
    .B(_08604_),
    .Y(_08607_));
 sky130_fd_sc_hd__a21oi_1 _16125_ (.A1(_08605_),
    .A2(_08606_),
    .B1(_08607_),
    .Y(_08608_));
 sky130_fd_sc_hd__nand2_1 _16126_ (.A(_08602_),
    .B(_08608_),
    .Y(_08609_));
 sky130_fd_sc_hd__nor2_1 _16127_ (.A(_08602_),
    .B(_08608_),
    .Y(_08610_));
 sky130_fd_sc_hd__a21oi_1 _16128_ (.A1(_08601_),
    .A2(_08609_),
    .B1(_08610_),
    .Y(_08611_));
 sky130_fd_sc_hd__xor2_1 _16129_ (.A(_08598_),
    .B(_08611_),
    .X(_08612_));
 sky130_fd_sc_hd__nor2_1 _16130_ (.A(_08598_),
    .B(_08611_),
    .Y(_08613_));
 sky130_fd_sc_hd__a21o_1 _16131_ (.A1(_08330_),
    .A2(_08612_),
    .B1(_08613_),
    .X(_08614_));
 sky130_fd_sc_hd__xnor2_1 _16132_ (.A(_08330_),
    .B(_08612_),
    .Y(_08615_));
 sky130_fd_sc_hd__xnor2_1 _16133_ (.A(_08602_),
    .B(_08608_),
    .Y(_08616_));
 sky130_fd_sc_hd__xnor2_1 _16134_ (.A(_08601_),
    .B(_08616_),
    .Y(_08617_));
 sky130_fd_sc_hd__xnor2_1 _16135_ (.A(_08322_),
    .B(_08435_),
    .Y(_08618_));
 sky130_fd_sc_hd__xnor2_1 _16136_ (.A(_08328_),
    .B(_08618_),
    .Y(_08619_));
 sky130_fd_sc_hd__or2_1 _16137_ (.A(_07689_),
    .B(_08403_),
    .X(_08620_));
 sky130_fd_sc_hd__nand2_1 _16138_ (.A(_08603_),
    .B(_08620_),
    .Y(_08621_));
 sky130_fd_sc_hd__and2b_1 _16139_ (.A_N(_08607_),
    .B(_08605_),
    .X(_08622_));
 sky130_fd_sc_hd__xnor2_1 _16140_ (.A(_08622_),
    .B(_08606_),
    .Y(_08623_));
 sky130_fd_sc_hd__nand2_1 _16141_ (.A(_08322_),
    .B(_08435_),
    .Y(_08624_));
 sky130_fd_sc_hd__o21ai_1 _16142_ (.A1(_08328_),
    .A2(_08618_),
    .B1(_08624_),
    .Y(_08625_));
 sky130_fd_sc_hd__inv_2 _16143_ (.A(_08625_),
    .Y(_08626_));
 sky130_fd_sc_hd__or2_1 _16144_ (.A(_08619_),
    .B(_08621_),
    .X(_08627_));
 sky130_fd_sc_hd__xnor2_1 _16145_ (.A(_08627_),
    .B(_08623_),
    .Y(_08628_));
 sky130_fd_sc_hd__o32a_1 _16146_ (.A1(_08619_),
    .A2(_08621_),
    .A3(_08623_),
    .B1(_08626_),
    .B2(_08628_),
    .X(_08629_));
 sky130_fd_sc_hd__xnor2_1 _16147_ (.A(_08617_),
    .B(_08629_),
    .Y(_08630_));
 sky130_fd_sc_hd__and2b_1 _16148_ (.A_N(_08629_),
    .B(_08617_),
    .X(_08631_));
 sky130_fd_sc_hd__a21oi_1 _16149_ (.A1(_08365_),
    .A2(_08630_),
    .B1(_08631_),
    .Y(_08632_));
 sky130_fd_sc_hd__o2bb2a_1 _16150_ (.A1_N(_08597_),
    .A2_N(_08614_),
    .B1(_08615_),
    .B2(_08632_),
    .X(_08633_));
 sky130_fd_sc_hd__xnor2_1 _16151_ (.A(_08166_),
    .B(_08630_),
    .Y(_08634_));
 sky130_fd_sc_hd__xnor2_1 _16152_ (.A(_08619_),
    .B(_08621_),
    .Y(_08635_));
 sky130_fd_sc_hd__a21bo_1 _16153_ (.A1(_08364_),
    .A2(_08434_),
    .B1_N(_08370_),
    .X(_08636_));
 sky130_fd_sc_hd__or2b_1 _16154_ (.A(_08635_),
    .B_N(_08636_),
    .X(_08637_));
 sky130_fd_sc_hd__xnor2_1 _16155_ (.A(_08625_),
    .B(_08628_),
    .Y(_08638_));
 sky130_fd_sc_hd__xnor2_1 _16156_ (.A(_08637_),
    .B(_08638_),
    .Y(_08639_));
 sky130_fd_sc_hd__and2b_1 _16157_ (.A_N(_08637_),
    .B(_08638_),
    .X(_08640_));
 sky130_fd_sc_hd__a21o_1 _16158_ (.A1(_08407_),
    .A2(_08639_),
    .B1(_08640_),
    .X(_08641_));
 sky130_fd_sc_hd__xnor2_1 _16159_ (.A(_08202_),
    .B(_08639_),
    .Y(_08642_));
 sky130_fd_sc_hd__xnor2_1 _16160_ (.A(_08364_),
    .B(_08434_),
    .Y(_08643_));
 sky130_fd_sc_hd__a21bo_1 _16161_ (.A1(_08399_),
    .A2(_08406_),
    .B1_N(_08412_),
    .X(_08644_));
 sky130_fd_sc_hd__and2b_1 _16162_ (.A_N(_08643_),
    .B(_08644_),
    .X(_08645_));
 sky130_fd_sc_hd__xnor2_1 _16163_ (.A(_08635_),
    .B(_08636_),
    .Y(_08646_));
 sky130_fd_sc_hd__xnor2_1 _16164_ (.A(_08645_),
    .B(_08646_),
    .Y(_08647_));
 sky130_fd_sc_hd__nand2_1 _16165_ (.A(_08645_),
    .B(_08646_),
    .Y(_08648_));
 sky130_fd_sc_hd__o21ai_1 _16166_ (.A1(_08222_),
    .A2(_08647_),
    .B1(_08648_),
    .Y(_08649_));
 sky130_fd_sc_hd__a22o_1 _16167_ (.A1(_08634_),
    .A2(_08641_),
    .B1(_08642_),
    .B2(_08649_),
    .X(_08650_));
 sky130_fd_sc_hd__xor2_1 _16168_ (.A(_08222_),
    .B(_08647_),
    .X(_08651_));
 sky130_fd_sc_hd__xor2_1 _16169_ (.A(_08643_),
    .B(_08644_),
    .X(_08652_));
 sky130_fd_sc_hd__xnor2_2 _16170_ (.A(_08399_),
    .B(_08406_),
    .Y(_08653_));
 sky130_fd_sc_hd__a21oi_1 _16171_ (.A1(_07689_),
    .A2(_08437_),
    .B1(_08442_),
    .Y(_08654_));
 sky130_fd_sc_hd__nor2_1 _16172_ (.A(_08653_),
    .B(_08654_),
    .Y(_08655_));
 sky130_fd_sc_hd__xnor2_1 _16173_ (.A(_08652_),
    .B(_08655_),
    .Y(_08656_));
 sky130_fd_sc_hd__or2b_1 _16174_ (.A(_08263_),
    .B_N(_08656_),
    .X(_08657_));
 sky130_fd_sc_hd__o31ai_1 _16175_ (.A1(_08652_),
    .A2(_08653_),
    .A3(_08654_),
    .B1(_08657_),
    .Y(_08658_));
 sky130_fd_sc_hd__or2_1 _16176_ (.A(_08651_),
    .B(_08658_),
    .X(_08659_));
 sky130_fd_sc_hd__xor2_1 _16177_ (.A(_08263_),
    .B(_08656_),
    .X(_08660_));
 sky130_fd_sc_hd__xnor2_1 _16178_ (.A(_07689_),
    .B(_08437_),
    .Y(_08661_));
 sky130_fd_sc_hd__nor2_1 _16179_ (.A(_08466_),
    .B(_08661_),
    .Y(_08662_));
 sky130_fd_sc_hd__xor2_1 _16180_ (.A(_08653_),
    .B(_08654_),
    .X(_08663_));
 sky130_fd_sc_hd__xnor2_1 _16181_ (.A(_08662_),
    .B(_08663_),
    .Y(_08664_));
 sky130_fd_sc_hd__nand2_1 _16182_ (.A(_08662_),
    .B(_08663_),
    .Y(_08665_));
 sky130_fd_sc_hd__o21a_1 _16183_ (.A1(_08273_),
    .A2(_08664_),
    .B1(_08665_),
    .X(_08666_));
 sky130_fd_sc_hd__nand2_1 _16184_ (.A(_08660_),
    .B(_08666_),
    .Y(_08667_));
 sky130_fd_sc_hd__or2_1 _16185_ (.A(_08273_),
    .B(_08664_),
    .X(_08668_));
 sky130_fd_sc_hd__xor2_1 _16186_ (.A(_08466_),
    .B(_08661_),
    .X(_08669_));
 sky130_fd_sc_hd__nand2_1 _16187_ (.A(_08464_),
    .B(_08501_),
    .Y(_08670_));
 sky130_fd_sc_hd__nor2_1 _16188_ (.A(_08295_),
    .B(_08670_),
    .Y(_08671_));
 sky130_fd_sc_hd__nand2_1 _16189_ (.A(_08295_),
    .B(_08670_),
    .Y(_08672_));
 sky130_fd_sc_hd__o21ai_1 _16190_ (.A1(_08669_),
    .A2(_08671_),
    .B1(_08672_),
    .Y(_08673_));
 sky130_fd_sc_hd__nand2_1 _16191_ (.A(_07668_),
    .B(_08673_),
    .Y(_08674_));
 sky130_fd_sc_hd__nand2_1 _16192_ (.A(_08273_),
    .B(_08664_),
    .Y(_08675_));
 sky130_fd_sc_hd__nor2_1 _16193_ (.A(_07668_),
    .B(_08673_),
    .Y(_08676_));
 sky130_fd_sc_hd__a31o_1 _16194_ (.A1(_08668_),
    .A2(_08674_),
    .A3(_08675_),
    .B1(_08676_),
    .X(_08677_));
 sky130_fd_sc_hd__nor2_1 _16195_ (.A(_08660_),
    .B(_08666_),
    .Y(_08678_));
 sky130_fd_sc_hd__a221o_1 _16196_ (.A1(_08651_),
    .A2(_08658_),
    .B1(_08667_),
    .B2(_08677_),
    .C1(_08678_),
    .X(_08679_));
 sky130_fd_sc_hd__o211a_1 _16197_ (.A1(_08642_),
    .A2(_08649_),
    .B1(_08659_),
    .C1(_08679_),
    .X(_08680_));
 sky130_fd_sc_hd__o2bb2a_1 _16198_ (.A1_N(_08615_),
    .A2_N(_08632_),
    .B1(_08634_),
    .B2(_08641_),
    .X(_08681_));
 sky130_fd_sc_hd__o21ai_1 _16199_ (.A1(_08650_),
    .A2(_08680_),
    .B1(_08681_),
    .Y(_08682_));
 sky130_fd_sc_hd__a2bb2o_2 _16200_ (.A1_N(_08597_),
    .A2_N(_08614_),
    .B1(_08633_),
    .B2(_08682_),
    .X(_08683_));
 sky130_fd_sc_hd__and3_1 _16201_ (.A(_08595_),
    .B(_08590_),
    .C(_08593_),
    .X(_08684_));
 sky130_fd_sc_hd__a21o_1 _16202_ (.A1(_08596_),
    .A2(_08683_),
    .B1(_08684_),
    .X(_08685_));
 sky130_fd_sc_hd__xor2_1 _16203_ (.A(_08521_),
    .B(_08544_),
    .X(_08686_));
 sky130_fd_sc_hd__or3b_1 _16204_ (.A(_08520_),
    .B(_08686_),
    .C_N(_08549_),
    .X(_08687_));
 sky130_fd_sc_hd__inv_2 _16205_ (.A(_08548_),
    .Y(_08688_));
 sky130_fd_sc_hd__nor3_2 _16206_ (.A(_08573_),
    .B(_08570_),
    .C(_08572_),
    .Y(_08689_));
 sky130_fd_sc_hd__a2111oi_2 _16207_ (.A1(_08575_),
    .A2(_08685_),
    .B1(_08687_),
    .C1(_08688_),
    .D1(_08689_),
    .Y(_08690_));
 sky130_fd_sc_hd__or2_1 _16208_ (.A(_08065_),
    .B(_08387_),
    .X(_08691_));
 sky130_fd_sc_hd__nand2_1 _16209_ (.A(_08388_),
    .B(_08691_),
    .Y(_08692_));
 sky130_fd_sc_hd__nand2_1 _16210_ (.A(_08393_),
    .B(_08424_),
    .Y(_08693_));
 sky130_fd_sc_hd__a21bo_1 _16211_ (.A1(_08065_),
    .A2(_08425_),
    .B1_N(_08693_),
    .X(_08694_));
 sky130_fd_sc_hd__xnor2_2 _16212_ (.A(_08692_),
    .B(_08694_),
    .Y(_08695_));
 sky130_fd_sc_hd__o31a_1 _16213_ (.A1(_08490_),
    .A2(_08550_),
    .A3(_08690_),
    .B1(_08695_),
    .X(_08696_));
 sky130_fd_sc_hd__and2_1 _16214_ (.A(_08392_),
    .B(_08696_),
    .X(_08697_));
 sky130_fd_sc_hd__and3_1 _16215_ (.A(_08388_),
    .B(_08691_),
    .C(_08694_),
    .X(_08698_));
 sky130_fd_sc_hd__o21a_1 _16216_ (.A1(_08391_),
    .A2(_08698_),
    .B1(_08389_),
    .X(_08699_));
 sky130_fd_sc_hd__or2b_1 _16217_ (.A(_08266_),
    .B_N(_08267_),
    .X(_08700_));
 sky130_fd_sc_hd__o21a_1 _16218_ (.A1(_08268_),
    .A2(_08269_),
    .B1(_08700_),
    .X(_08701_));
 sky130_fd_sc_hd__xor2_1 _16219_ (.A(_08227_),
    .B(_08231_),
    .X(_08702_));
 sky130_fd_sc_hd__and2b_1 _16220_ (.A_N(_08701_),
    .B(_08702_),
    .X(_08703_));
 sky130_fd_sc_hd__and2b_1 _16221_ (.A_N(_08702_),
    .B(_08701_),
    .X(_08704_));
 sky130_fd_sc_hd__nor2_1 _16222_ (.A(_08703_),
    .B(_08704_),
    .Y(_08705_));
 sky130_fd_sc_hd__a21oi_1 _16223_ (.A1(_08101_),
    .A2(_08330_),
    .B1(_08105_),
    .Y(_08706_));
 sky130_fd_sc_hd__inv_2 _16224_ (.A(_08706_),
    .Y(_08707_));
 sky130_fd_sc_hd__a21oi_1 _16225_ (.A1(_08705_),
    .A2(_08707_),
    .B1(_08703_),
    .Y(_08708_));
 sky130_fd_sc_hd__xnor2_1 _16226_ (.A(_08235_),
    .B(_08234_),
    .Y(_08709_));
 sky130_fd_sc_hd__and2b_1 _16227_ (.A_N(_08708_),
    .B(_08709_),
    .X(_08710_));
 sky130_fd_sc_hd__and2b_1 _16228_ (.A_N(_08709_),
    .B(_08708_),
    .X(_08711_));
 sky130_fd_sc_hd__nor2_1 _16229_ (.A(_08710_),
    .B(_08711_),
    .Y(_08712_));
 sky130_fd_sc_hd__xnor2_1 _16230_ (.A(_08705_),
    .B(_08707_),
    .Y(_08713_));
 sky130_fd_sc_hd__a21oi_1 _16231_ (.A1(_08284_),
    .A2(_08289_),
    .B1(_08283_),
    .Y(_08714_));
 sky130_fd_sc_hd__or2_1 _16232_ (.A(_08713_),
    .B(_08714_),
    .X(_08715_));
 sky130_fd_sc_hd__nand2_1 _16233_ (.A(_08713_),
    .B(_08714_),
    .Y(_08716_));
 sky130_fd_sc_hd__nand2_1 _16234_ (.A(_08715_),
    .B(_08716_),
    .Y(_08717_));
 sky130_fd_sc_hd__nor2_1 _16235_ (.A(_06410_),
    .B(_08287_),
    .Y(_08718_));
 sky130_fd_sc_hd__a21oi_1 _16236_ (.A1(_08130_),
    .A2(_08288_),
    .B1(_08718_),
    .Y(_08719_));
 sky130_fd_sc_hd__o21a_1 _16237_ (.A1(_08717_),
    .A2(_08719_),
    .B1(_08715_),
    .X(_08720_));
 sky130_fd_sc_hd__xor2_1 _16238_ (.A(_08712_),
    .B(_08720_),
    .X(_08721_));
 sky130_fd_sc_hd__or2b_1 _16239_ (.A(_08316_),
    .B_N(_08290_),
    .X(_08722_));
 sky130_fd_sc_hd__or2_1 _16240_ (.A(_08317_),
    .B(_08318_),
    .X(_08723_));
 sky130_fd_sc_hd__xnor2_1 _16241_ (.A(_08717_),
    .B(_08719_),
    .Y(_08724_));
 sky130_fd_sc_hd__a21o_1 _16242_ (.A1(_08722_),
    .A2(_08723_),
    .B1(_08724_),
    .X(_08725_));
 sky130_fd_sc_hd__nand3_1 _16243_ (.A(_08722_),
    .B(_08723_),
    .C(_08724_),
    .Y(_08726_));
 sky130_fd_sc_hd__and2_1 _16244_ (.A(_08725_),
    .B(_08726_),
    .X(_08727_));
 sky130_fd_sc_hd__nand2_1 _16245_ (.A(_08066_),
    .B(_08727_),
    .Y(_08728_));
 sky130_fd_sc_hd__nand3_1 _16246_ (.A(_08721_),
    .B(_08725_),
    .C(_08728_),
    .Y(_08729_));
 sky130_fd_sc_hd__or2b_1 _16247_ (.A(_08319_),
    .B_N(_08349_),
    .X(_08730_));
 sky130_fd_sc_hd__xnor2_1 _16248_ (.A(_08066_),
    .B(_08727_),
    .Y(_08731_));
 sky130_fd_sc_hd__a21oi_1 _16249_ (.A1(_08730_),
    .A2(_08351_),
    .B1(_08731_),
    .Y(_08732_));
 sky130_fd_sc_hd__a21oi_1 _16250_ (.A1(_08725_),
    .A2(_08728_),
    .B1(_08721_),
    .Y(_08733_));
 sky130_fd_sc_hd__a21o_1 _16251_ (.A1(_08729_),
    .A2(_08732_),
    .B1(_08733_),
    .X(_08734_));
 sky130_fd_sc_hd__nand3_1 _16252_ (.A(_08730_),
    .B(_08351_),
    .C(_08731_),
    .Y(_08735_));
 sky130_fd_sc_hd__o21a_1 _16253_ (.A1(_08733_),
    .A2(_08735_),
    .B1(_08729_),
    .X(_08736_));
 sky130_fd_sc_hd__a21oi_1 _16254_ (.A1(_08065_),
    .A2(_08712_),
    .B1(_08710_),
    .Y(_08737_));
 sky130_fd_sc_hd__xnor2_1 _16255_ (.A(_08240_),
    .B(_08737_),
    .Y(_08738_));
 sky130_fd_sc_hd__inv_2 _16256_ (.A(_08720_),
    .Y(_08739_));
 sky130_fd_sc_hd__mux2_1 _16257_ (.A0(_08066_),
    .A1(_08739_),
    .S(_08712_),
    .X(_08740_));
 sky130_fd_sc_hd__nand2_1 _16258_ (.A(_08738_),
    .B(_08740_),
    .Y(_08741_));
 sky130_fd_sc_hd__or2_1 _16259_ (.A(_08738_),
    .B(_08740_),
    .X(_08742_));
 sky130_fd_sc_hd__and2_1 _16260_ (.A(_08741_),
    .B(_08742_),
    .X(_08743_));
 sky130_fd_sc_hd__o311a_2 _16261_ (.A1(_08697_),
    .A2(_08699_),
    .A3(_08734_),
    .B1(_08736_),
    .C1(_08743_),
    .X(_08744_));
 sky130_fd_sc_hd__xnor2_1 _16262_ (.A(_08066_),
    .B(_08247_),
    .Y(_08745_));
 sky130_fd_sc_hd__clkinv_2 _16263_ (.A(_08737_),
    .Y(_08746_));
 sky130_fd_sc_hd__mux2_1 _16264_ (.A0(_08066_),
    .A1(_08746_),
    .S(_08240_),
    .X(_08747_));
 sky130_fd_sc_hd__or2b_1 _16265_ (.A(_08745_),
    .B_N(_08747_),
    .X(_08748_));
 sky130_fd_sc_hd__and2_1 _16266_ (.A(_08741_),
    .B(_08748_),
    .X(_08749_));
 sky130_fd_sc_hd__inv_2 _16267_ (.A(_08749_),
    .Y(_08750_));
 sky130_fd_sc_hd__nand3_1 _16268_ (.A(_08256_),
    .B(_08245_),
    .C(_08248_),
    .Y(_08751_));
 sky130_fd_sc_hd__nand2_1 _16269_ (.A(_08257_),
    .B(_08751_),
    .Y(_08752_));
 sky130_fd_sc_hd__inv_2 _16270_ (.A(_08752_),
    .Y(_08753_));
 sky130_fd_sc_hd__and2b_1 _16271_ (.A_N(_08747_),
    .B(_08745_),
    .X(_08754_));
 sky130_fd_sc_hd__inv_2 _16272_ (.A(_08754_),
    .Y(_08755_));
 sky130_fd_sc_hd__o211ai_4 _16273_ (.A1(_08744_),
    .A2(_08750_),
    .B1(_08753_),
    .C1(_08755_),
    .Y(_08756_));
 sky130_fd_sc_hd__a21o_1 _16274_ (.A1(_08163_),
    .A2(_08164_),
    .B1(_08185_),
    .X(_08757_));
 sky130_fd_sc_hd__nand2_1 _16275_ (.A(_08186_),
    .B(_08757_),
    .Y(_08758_));
 sky130_fd_sc_hd__and3_1 _16276_ (.A(_08258_),
    .B(_08251_),
    .C(_08254_),
    .X(_08759_));
 sky130_fd_sc_hd__a211o_1 _16277_ (.A1(_08260_),
    .A2(_08756_),
    .B1(_08758_),
    .C1(_08759_),
    .X(_08760_));
 sky130_fd_sc_hd__and3_1 _16278_ (.A(_08196_),
    .B(_08160_),
    .C(_08163_),
    .X(_08761_));
 sky130_fd_sc_hd__a31o_1 _16279_ (.A1(_08186_),
    .A2(_08197_),
    .A3(_08760_),
    .B1(_08761_),
    .X(_08762_));
 sky130_fd_sc_hd__mux2_1 _16280_ (.A0(_08085_),
    .A1(_08195_),
    .S(_08194_),
    .X(_08763_));
 sky130_fd_sc_hd__nand2_1 _16281_ (.A(_08085_),
    .B(_08194_),
    .Y(_08764_));
 sky130_fd_sc_hd__a22o_1 _16282_ (.A1(_08085_),
    .A2(_08189_),
    .B1(_08192_),
    .B2(_08764_),
    .X(_08765_));
 sky130_fd_sc_hd__a21boi_1 _16283_ (.A1(_06410_),
    .A2(_08107_),
    .B1_N(_08765_),
    .Y(_08766_));
 sky130_fd_sc_hd__xnor2_1 _16284_ (.A(_08763_),
    .B(_08766_),
    .Y(_08767_));
 sky130_fd_sc_hd__xnor2_1 _16285_ (.A(_08762_),
    .B(_08767_),
    .Y(_08768_));
 sky130_fd_sc_hd__o21a_1 _16286_ (.A1(_08047_),
    .A2(_08051_),
    .B1(_08054_),
    .X(_08769_));
 sky130_fd_sc_hd__or2_1 _16287_ (.A(_08053_),
    .B(_08769_),
    .X(_08770_));
 sky130_fd_sc_hd__nor2_1 _16288_ (.A(_08081_),
    .B(_08055_),
    .Y(_08771_));
 sky130_fd_sc_hd__a22o_2 _16289_ (.A1(_08082_),
    .A2(_08768_),
    .B1(_08770_),
    .B2(_08771_),
    .X(_08772_));
 sky130_fd_sc_hd__clkbuf_8 _16290_ (.A(_06403_),
    .X(_08773_));
 sky130_fd_sc_hd__mux2_1 _16291_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.temp[30] ),
    .A1(_08772_),
    .S(_08773_),
    .X(_08774_));
 sky130_fd_sc_hd__clkbuf_1 _16292_ (.A(_08774_),
    .X(_00960_));
 sky130_fd_sc_hd__or2b_1 _16293_ (.A(_08761_),
    .B_N(_08197_),
    .X(_08775_));
 sky130_fd_sc_hd__a21oi_1 _16294_ (.A1(_08186_),
    .A2(_08760_),
    .B1(_08775_),
    .Y(_08776_));
 sky130_fd_sc_hd__a31o_1 _16295_ (.A1(_08186_),
    .A2(_08760_),
    .A3(_08775_),
    .B1(_06407_),
    .X(_08777_));
 sky130_fd_sc_hd__nand2_1 _16296_ (.A(_08054_),
    .B(_08050_),
    .Y(_08778_));
 sky130_fd_sc_hd__or2_1 _16297_ (.A(_08044_),
    .B(_08047_),
    .X(_08779_));
 sky130_fd_sc_hd__xnor2_1 _16298_ (.A(_08778_),
    .B(_08779_),
    .Y(_08780_));
 sky130_fd_sc_hd__a2bb2o_2 _16299_ (.A1_N(_08776_),
    .A2_N(_08777_),
    .B1(_08780_),
    .B2(_06408_),
    .X(_08781_));
 sky130_fd_sc_hd__mux2_1 _16300_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.temp[29] ),
    .A1(_08781_),
    .S(_08773_),
    .X(_08782_));
 sky130_fd_sc_hd__clkbuf_1 _16301_ (.A(_08782_),
    .X(_00959_));
 sky130_fd_sc_hd__a21o_1 _16302_ (.A1(_08260_),
    .A2(_08756_),
    .B1(_08759_),
    .X(_08783_));
 sky130_fd_sc_hd__a21oi_1 _16303_ (.A1(_08758_),
    .A2(_08783_),
    .B1(_06408_),
    .Y(_08784_));
 sky130_fd_sc_hd__a22o_1 _16304_ (.A1(_07976_),
    .A2(_08032_),
    .B1(_08035_),
    .B2(_08031_),
    .X(_08785_));
 sky130_fd_sc_hd__or2_1 _16305_ (.A(_06406_),
    .B(_08047_),
    .X(_08786_));
 sky130_fd_sc_hd__a21o_1 _16306_ (.A1(_08046_),
    .A2(_08785_),
    .B1(_08786_),
    .X(_08787_));
 sky130_fd_sc_hd__a21bo_2 _16307_ (.A1(_08760_),
    .A2(_08784_),
    .B1_N(_08787_),
    .X(_08788_));
 sky130_fd_sc_hd__mux2_1 _16308_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.temp[28] ),
    .A1(_08788_),
    .S(_08773_),
    .X(_08789_));
 sky130_fd_sc_hd__clkbuf_1 _16309_ (.A(_08789_),
    .X(_00958_));
 sky130_fd_sc_hd__or2b_1 _16310_ (.A(_08759_),
    .B_N(_08259_),
    .X(_08790_));
 sky130_fd_sc_hd__nand3_1 _16311_ (.A(_08257_),
    .B(_08756_),
    .C(_08790_),
    .Y(_08791_));
 sky130_fd_sc_hd__a21o_1 _16312_ (.A1(_08257_),
    .A2(_08756_),
    .B1(_08790_),
    .X(_08792_));
 sky130_fd_sc_hd__a21oi_1 _16313_ (.A1(_07976_),
    .A2(_07977_),
    .B1(_08034_),
    .Y(_08793_));
 sky130_fd_sc_hd__nor2_1 _16314_ (.A(_08029_),
    .B(_08793_),
    .Y(_08794_));
 sky130_fd_sc_hd__nand2_1 _16315_ (.A(_08033_),
    .B(_08794_),
    .Y(_08795_));
 sky130_fd_sc_hd__o21a_1 _16316_ (.A1(_08033_),
    .A2(_08794_),
    .B1(_06407_),
    .X(_08796_));
 sky130_fd_sc_hd__a32o_2 _16317_ (.A1(_08082_),
    .A2(_08791_),
    .A3(_08792_),
    .B1(_08795_),
    .B2(_08796_),
    .X(_08797_));
 sky130_fd_sc_hd__mux2_1 _16318_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.temp[27] ),
    .A1(_08797_),
    .S(_08773_),
    .X(_08798_));
 sky130_fd_sc_hd__clkbuf_1 _16319_ (.A(_08798_),
    .X(_00957_));
 sky130_fd_sc_hd__o21a_1 _16320_ (.A1(_08744_),
    .A2(_08750_),
    .B1(_08755_),
    .X(_08799_));
 sky130_fd_sc_hd__nor2_1 _16321_ (.A(_08753_),
    .B(_08799_),
    .Y(_08800_));
 sky130_fd_sc_hd__nand2_1 _16322_ (.A(_08082_),
    .B(_08756_),
    .Y(_08801_));
 sky130_fd_sc_hd__and3_1 _16323_ (.A(_07976_),
    .B(_07977_),
    .C(_08034_),
    .X(_08802_));
 sky130_fd_sc_hd__or3_1 _16324_ (.A(_08081_),
    .B(_08793_),
    .C(_08802_),
    .X(_08803_));
 sky130_fd_sc_hd__o211a_1 _16325_ (.A1(_08800_),
    .A2(_08801_),
    .B1(_06404_),
    .C1(_08803_),
    .X(_08804_));
 sky130_fd_sc_hd__o21ba_1 _16326_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.temp[26] ),
    .A2(_06404_),
    .B1_N(_08804_),
    .X(_00956_));
 sky130_fd_sc_hd__o31a_1 _16327_ (.A1(_08697_),
    .A2(_08699_),
    .A3(_08734_),
    .B1(_08736_),
    .X(_08805_));
 sky130_fd_sc_hd__nand2_1 _16328_ (.A(_08743_),
    .B(_08805_),
    .Y(_08806_));
 sky130_fd_sc_hd__nand2_1 _16329_ (.A(_08755_),
    .B(_08748_),
    .Y(_08807_));
 sky130_fd_sc_hd__a31o_1 _16330_ (.A1(_08741_),
    .A2(_08806_),
    .A3(_08807_),
    .B1(_06407_),
    .X(_08808_));
 sky130_fd_sc_hd__a21oi_1 _16331_ (.A1(_08741_),
    .A2(_08806_),
    .B1(_08807_),
    .Y(_08809_));
 sky130_fd_sc_hd__o21a_1 _16332_ (.A1(_07970_),
    .A2(_07975_),
    .B1(_07973_),
    .X(_08810_));
 sky130_fd_sc_hd__o21a_1 _16333_ (.A1(_06964_),
    .A2(_08810_),
    .B1(_06407_),
    .X(_08811_));
 sky130_fd_sc_hd__nand2_1 _16334_ (.A(_06964_),
    .B(_08810_),
    .Y(_08812_));
 sky130_fd_sc_hd__a2bb2o_1 _16335_ (.A1_N(_08808_),
    .A2_N(_08809_),
    .B1(_08811_),
    .B2(_08812_),
    .X(_08813_));
 sky130_fd_sc_hd__mux2_1 _16336_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.temp[25] ),
    .A1(_08813_),
    .S(_08773_),
    .X(_08814_));
 sky130_fd_sc_hd__clkbuf_1 _16337_ (.A(_08814_),
    .X(_00955_));
 sky130_fd_sc_hd__nor2_1 _16338_ (.A(_08743_),
    .B(_08805_),
    .Y(_08815_));
 sky130_fd_sc_hd__nor2_1 _16339_ (.A(_07970_),
    .B(_07975_),
    .Y(_08816_));
 sky130_fd_sc_hd__nand2_1 _16340_ (.A(_07970_),
    .B(_07975_),
    .Y(_08817_));
 sky130_fd_sc_hd__or3b_2 _16341_ (.A(_08081_),
    .B(_08816_),
    .C_N(_08817_),
    .X(_08818_));
 sky130_fd_sc_hd__o31ai_4 _16342_ (.A1(_06408_),
    .A2(_08744_),
    .A3(_08815_),
    .B1(_08818_),
    .Y(_08819_));
 sky130_fd_sc_hd__mux2_1 _16343_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.temp[24] ),
    .A1(_08819_),
    .S(_08773_),
    .X(_08820_));
 sky130_fd_sc_hd__clkbuf_1 _16344_ (.A(_08820_),
    .X(_00954_));
 sky130_fd_sc_hd__a21oi_1 _16345_ (.A1(_07934_),
    .A2(_07936_),
    .B1(_07968_),
    .Y(_08821_));
 sky130_fd_sc_hd__nor2_1 _16346_ (.A(_07963_),
    .B(_08821_),
    .Y(_08822_));
 sky130_fd_sc_hd__xnor2_1 _16347_ (.A(_07966_),
    .B(_08822_),
    .Y(_08823_));
 sky130_fd_sc_hd__or2b_1 _16348_ (.A(_08733_),
    .B_N(_08729_),
    .X(_08824_));
 sky130_fd_sc_hd__and2b_1 _16349_ (.A_N(_08732_),
    .B(_08735_),
    .X(_08825_));
 sky130_fd_sc_hd__o21a_1 _16350_ (.A1(_08697_),
    .A2(_08699_),
    .B1(_08825_),
    .X(_08826_));
 sky130_fd_sc_hd__nor2_1 _16351_ (.A(_08732_),
    .B(_08826_),
    .Y(_08827_));
 sky130_fd_sc_hd__o21ai_1 _16352_ (.A1(_08824_),
    .A2(_08827_),
    .B1(_08081_),
    .Y(_08828_));
 sky130_fd_sc_hd__a21o_1 _16353_ (.A1(_08824_),
    .A2(_08827_),
    .B1(_08828_),
    .X(_08829_));
 sky130_fd_sc_hd__o211a_1 _16354_ (.A1(_08082_),
    .A2(_08823_),
    .B1(_08829_),
    .C1(_06404_),
    .X(_08830_));
 sky130_fd_sc_hd__o21ba_1 _16355_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.temp[23] ),
    .A2(_06404_),
    .B1_N(_08830_),
    .X(_00953_));
 sky130_fd_sc_hd__nor3_1 _16356_ (.A(_08697_),
    .B(_08699_),
    .C(_08825_),
    .Y(_08831_));
 sky130_fd_sc_hd__and3_1 _16357_ (.A(_07934_),
    .B(_07936_),
    .C(_07968_),
    .X(_08832_));
 sky130_fd_sc_hd__or3_4 _16358_ (.A(_08081_),
    .B(_08821_),
    .C(_08832_),
    .X(_08833_));
 sky130_fd_sc_hd__o31ai_4 _16359_ (.A1(_06408_),
    .A2(_08826_),
    .A3(_08831_),
    .B1(_08833_),
    .Y(_08834_));
 sky130_fd_sc_hd__mux2_1 _16360_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.temp[22] ),
    .A1(_08834_),
    .S(_08773_),
    .X(_08835_));
 sky130_fd_sc_hd__clkbuf_1 _16361_ (.A(_08835_),
    .X(_00952_));
 sky130_fd_sc_hd__nand2_1 _16362_ (.A(_07481_),
    .B(_07858_),
    .Y(_08836_));
 sky130_fd_sc_hd__a21boi_1 _16363_ (.A1(_08836_),
    .A2(_07932_),
    .B1_N(_07935_),
    .Y(_08837_));
 sky130_fd_sc_hd__xnor2_1 _16364_ (.A(_07928_),
    .B(_08837_),
    .Y(_08838_));
 sky130_fd_sc_hd__o21a_1 _16365_ (.A1(_08698_),
    .A2(_08696_),
    .B1(_08392_),
    .X(_08839_));
 sky130_fd_sc_hd__or3_1 _16366_ (.A(_08392_),
    .B(_08698_),
    .C(_08696_),
    .X(_08840_));
 sky130_fd_sc_hd__or3b_4 _16367_ (.A(_08839_),
    .B(_06408_),
    .C_N(_08840_),
    .X(_08841_));
 sky130_fd_sc_hd__o211a_1 _16368_ (.A1(_08082_),
    .A2(_08838_),
    .B1(_08841_),
    .C1(_06404_),
    .X(_08842_));
 sky130_fd_sc_hd__o21ba_1 _16369_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.temp[21] ),
    .A2(_06404_),
    .B1_N(_08842_),
    .X(_00951_));
 sky130_fd_sc_hd__o41ai_1 _16370_ (.A1(_08490_),
    .A2(_08550_),
    .A3(_08690_),
    .A4(_08695_),
    .B1(_08081_),
    .Y(_08843_));
 sky130_fd_sc_hd__xor2_2 _16371_ (.A(_08836_),
    .B(_07932_),
    .X(_08844_));
 sky130_fd_sc_hd__a2bb2o_2 _16372_ (.A1_N(_08843_),
    .A2_N(_08696_),
    .B1(_06408_),
    .B2(_08844_),
    .X(_08845_));
 sky130_fd_sc_hd__mux2_1 _16373_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.temp[20] ),
    .A1(_08845_),
    .S(_08773_),
    .X(_08846_));
 sky130_fd_sc_hd__clkbuf_1 _16374_ (.A(_08846_),
    .X(_00950_));
 sky130_fd_sc_hd__inv_2 _16375_ (.A(_07855_),
    .Y(_08847_));
 sky130_fd_sc_hd__a21o_1 _16376_ (.A1(_07539_),
    .A2(_07854_),
    .B1(_08847_),
    .X(_08848_));
 sky130_fd_sc_hd__o21ai_1 _16377_ (.A1(_07341_),
    .A2(_08848_),
    .B1(_07342_),
    .Y(_08849_));
 sky130_fd_sc_hd__a21oi_1 _16378_ (.A1(_07411_),
    .A2(_08849_),
    .B1(_07478_),
    .Y(_08850_));
 sky130_fd_sc_hd__xnor2_1 _16379_ (.A(_08850_),
    .B(_07476_),
    .Y(_08851_));
 sky130_fd_sc_hd__a21o_1 _16380_ (.A1(_08575_),
    .A2(_08685_),
    .B1(_08689_),
    .X(_08852_));
 sky130_fd_sc_hd__or2_2 _16381_ (.A(_08852_),
    .B(_08686_),
    .X(_08853_));
 sky130_fd_sc_hd__or2b_1 _16382_ (.A(_08545_),
    .B_N(_08853_),
    .X(_08854_));
 sky130_fd_sc_hd__a21o_1 _16383_ (.A1(_08549_),
    .A2(_08854_),
    .B1(_08520_),
    .X(_08855_));
 sky130_fd_sc_hd__and2_1 _16384_ (.A(_08546_),
    .B(_08855_),
    .X(_08856_));
 sky130_fd_sc_hd__or2_1 _16385_ (.A(_08488_),
    .B(_08856_),
    .X(_08857_));
 sky130_fd_sc_hd__xor2_2 _16386_ (.A(_08857_),
    .B(_08547_),
    .X(_08858_));
 sky130_fd_sc_hd__mux2_1 _16387_ (.A0(_08851_),
    .A1(_08858_),
    .S(_08081_),
    .X(_08859_));
 sky130_fd_sc_hd__mux2_1 _16388_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.temp[19] ),
    .A1(_08859_),
    .S(_08773_),
    .X(_08860_));
 sky130_fd_sc_hd__clkbuf_1 _16389_ (.A(_08860_),
    .X(_00949_));
 sky130_fd_sc_hd__xnor2_1 _16390_ (.A(_07411_),
    .B(_08849_),
    .Y(_08861_));
 sky130_fd_sc_hd__or2_2 _16391_ (.A(_08546_),
    .B(_08855_),
    .X(_08862_));
 sky130_fd_sc_hd__nor2_2 _16392_ (.A(_06407_),
    .B(_08856_),
    .Y(_08863_));
 sky130_fd_sc_hd__a2bb2o_1 _16393_ (.A1_N(_08082_),
    .A2_N(_08861_),
    .B1(_08862_),
    .B2(_08863_),
    .X(_08864_));
 sky130_fd_sc_hd__mux2_1 _16394_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.temp[18] ),
    .A1(_08864_),
    .S(_06403_),
    .X(_08865_));
 sky130_fd_sc_hd__clkbuf_1 _16395_ (.A(_08865_),
    .X(_00948_));
 sky130_fd_sc_hd__and2b_1 _16396_ (.A_N(_08520_),
    .B(_08549_),
    .X(_08866_));
 sky130_fd_sc_hd__nand2_1 _16397_ (.A(_08854_),
    .B(_08866_),
    .Y(_08867_));
 sky130_fd_sc_hd__or2_2 _16398_ (.A(_08854_),
    .B(_08866_),
    .X(_08868_));
 sky130_fd_sc_hd__nand2_1 _16399_ (.A(_07340_),
    .B(_08848_),
    .Y(_08869_));
 sky130_fd_sc_hd__nand2_1 _16400_ (.A(_08869_),
    .B(_07856_),
    .Y(_08870_));
 sky130_fd_sc_hd__o21a_1 _16401_ (.A1(_08869_),
    .A2(_07856_),
    .B1(_06407_),
    .X(_08871_));
 sky130_fd_sc_hd__a32o_1 _16402_ (.A1(_08082_),
    .A2(_08867_),
    .A3(_08868_),
    .B1(_08870_),
    .B2(_08871_),
    .X(_08872_));
 sky130_fd_sc_hd__mux2_1 _16403_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.temp[17] ),
    .A1(_08872_),
    .S(_06403_),
    .X(_08873_));
 sky130_fd_sc_hd__clkbuf_1 _16404_ (.A(_08873_),
    .X(_00947_));
 sky130_fd_sc_hd__nand3_1 _16405_ (.A(_07539_),
    .B(_07854_),
    .C(_08847_),
    .Y(_08874_));
 sky130_fd_sc_hd__a21oi_2 _16406_ (.A1(_08852_),
    .A2(_08686_),
    .B1(_06407_),
    .Y(_08875_));
 sky130_fd_sc_hd__a32o_1 _16407_ (.A1(_06408_),
    .A2(_08848_),
    .A3(_08874_),
    .B1(_08875_),
    .B2(_08853_),
    .X(_08876_));
 sky130_fd_sc_hd__mux2_1 _16408_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.temp[16] ),
    .A1(_08876_),
    .S(_06403_),
    .X(_08877_));
 sky130_fd_sc_hd__clkbuf_1 _16409_ (.A(_08877_),
    .X(_00946_));
 sky130_fd_sc_hd__a31o_1 _16410_ (.A1(_07593_),
    .A2(_07849_),
    .A3(_07851_),
    .B1(_07852_),
    .X(_08878_));
 sky130_fd_sc_hd__nor2_1 _16411_ (.A(_07538_),
    .B(_07853_),
    .Y(_08879_));
 sky130_fd_sc_hd__xnor2_2 _16412_ (.A(_08878_),
    .B(_08879_),
    .Y(_08880_));
 sky130_fd_sc_hd__o21ai_1 _16413_ (.A1(_08574_),
    .A2(_08689_),
    .B1(_08685_),
    .Y(_08881_));
 sky130_fd_sc_hd__o31a_1 _16414_ (.A1(_08574_),
    .A2(_08689_),
    .A3(_08685_),
    .B1(_08081_),
    .X(_08882_));
 sky130_fd_sc_hd__a22o_2 _16415_ (.A1(_06408_),
    .A2(_08880_),
    .B1(_08881_),
    .B2(_08882_),
    .X(_08883_));
 sky130_fd_sc_hd__mux2_1 _16416_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.temp[15] ),
    .A1(_08883_),
    .S(_06403_),
    .X(_08884_));
 sky130_fd_sc_hd__clkbuf_1 _16417_ (.A(_08884_),
    .X(_00945_));
 sky130_fd_sc_hd__inv_2 _16418_ (.A(\wfg_stim_sine_top.wfg_stim_sine.temp[14] ),
    .Y(_08885_));
 sky130_fd_sc_hd__nand2_2 _16419_ (.A(_07849_),
    .B(_07851_),
    .Y(_08886_));
 sky130_fd_sc_hd__or2_2 _16420_ (.A(_07592_),
    .B(_07852_),
    .X(_08887_));
 sky130_fd_sc_hd__xnor2_4 _16421_ (.A(_08886_),
    .B(_08887_),
    .Y(_08888_));
 sky130_fd_sc_hd__a21oi_1 _16422_ (.A1(_08590_),
    .A2(_08593_),
    .B1(_08595_),
    .Y(_08889_));
 sky130_fd_sc_hd__nor2_1 _16423_ (.A(_08889_),
    .B(_08684_),
    .Y(_08890_));
 sky130_fd_sc_hd__nor2_1 _16424_ (.A(_08683_),
    .B(_08890_),
    .Y(_08891_));
 sky130_fd_sc_hd__a21o_1 _16425_ (.A1(_08683_),
    .A2(_08890_),
    .B1(_06408_),
    .X(_08892_));
 sky130_fd_sc_hd__o221a_2 _16426_ (.A1(_08082_),
    .A2(_08888_),
    .B1(_08891_),
    .B2(_08892_),
    .C1(_06404_),
    .X(_08893_));
 sky130_fd_sc_hd__o21bai_1 _16427_ (.A1(_08885_),
    .A2(_06404_),
    .B1_N(_08893_),
    .Y(_00944_));
 sky130_fd_sc_hd__or2_1 _16428_ (.A(\wfg_stim_sine_top.wfg_stim_sine.cur_state[2] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.cur_state[1] ),
    .X(_08894_));
 sky130_fd_sc_hd__clkbuf_4 _16429_ (.A(_08894_),
    .X(_08895_));
 sky130_fd_sc_hd__clkbuf_4 _16430_ (.A(_08895_),
    .X(_08896_));
 sky130_fd_sc_hd__nor2_2 _16431_ (.A(\wfg_stim_sine_top.wfg_stim_sine.cur_state[2] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.cur_state[1] ),
    .Y(_08897_));
 sky130_fd_sc_hd__nand2_1 _16432_ (.A(\wfg_stim_sine_top.wfg_stim_sine.cur_state[0] ),
    .B(_08897_),
    .Y(_08898_));
 sky130_fd_sc_hd__clkbuf_4 _16433_ (.A(\wfg_stim_sine_top.wfg_stim_sine.iteration[1] ),
    .X(_08899_));
 sky130_fd_sc_hd__clkbuf_4 _16434_ (.A(_08899_),
    .X(_08900_));
 sky130_fd_sc_hd__clkbuf_4 _16435_ (.A(\wfg_stim_sine_top.wfg_stim_sine.iteration[0] ),
    .X(_08901_));
 sky130_fd_sc_hd__clkbuf_4 _16436_ (.A(_08901_),
    .X(_08902_));
 sky130_fd_sc_hd__nand2_2 _16437_ (.A(_08900_),
    .B(_08902_),
    .Y(_08903_));
 sky130_fd_sc_hd__clkbuf_4 _16438_ (.A(\wfg_stim_sine_top.wfg_stim_sine.iteration[2] ),
    .X(_08904_));
 sky130_fd_sc_hd__nand2_1 _16439_ (.A(\wfg_stim_sine_top.wfg_stim_sine.iteration[3] ),
    .B(_08904_),
    .Y(_08905_));
 sky130_fd_sc_hd__nor2_2 _16440_ (.A(_08903_),
    .B(_08905_),
    .Y(_08906_));
 sky130_fd_sc_hd__nor2_1 _16441_ (.A(_08898_),
    .B(_08906_),
    .Y(_08907_));
 sky130_fd_sc_hd__clkbuf_4 _16442_ (.A(_08904_),
    .X(_08908_));
 sky130_fd_sc_hd__buf_2 _16443_ (.A(_08908_),
    .X(_08909_));
 sky130_fd_sc_hd__clkbuf_4 _16444_ (.A(_08900_),
    .X(_08910_));
 sky130_fd_sc_hd__buf_2 _16445_ (.A(_08902_),
    .X(_08911_));
 sky130_fd_sc_hd__buf_4 _16446_ (.A(\wfg_stim_sine_top.wfg_stim_sine.iteration[3] ),
    .X(_08912_));
 sky130_fd_sc_hd__buf_2 _16447_ (.A(_08912_),
    .X(_08913_));
 sky130_fd_sc_hd__a41o_1 _16448_ (.A1(_08909_),
    .A2(_08910_),
    .A3(_08911_),
    .A4(_08897_),
    .B1(_08913_),
    .X(_08914_));
 sky130_fd_sc_hd__o21a_1 _16449_ (.A1(_08896_),
    .A2(_08907_),
    .B1(_08914_),
    .X(_00943_));
 sky130_fd_sc_hd__clkbuf_4 _16450_ (.A(_08898_),
    .X(_08915_));
 sky130_fd_sc_hd__buf_4 _16451_ (.A(_08915_),
    .X(_08916_));
 sky130_fd_sc_hd__xor2_1 _16452_ (.A(_08904_),
    .B(_08903_),
    .X(_08917_));
 sky130_fd_sc_hd__a2bb2o_1 _16453_ (.A1_N(_08916_),
    .A2_N(_08917_),
    .B1(_08909_),
    .B2(_08896_),
    .X(_00942_));
 sky130_fd_sc_hd__and2_2 _16454_ (.A(\wfg_stim_sine_top.wfg_stim_sine.cur_state[0] ),
    .B(_08897_),
    .X(_08918_));
 sky130_fd_sc_hd__clkbuf_8 _16455_ (.A(_08918_),
    .X(_08919_));
 sky130_fd_sc_hd__clkbuf_4 _16456_ (.A(\wfg_stim_sine_top.wfg_stim_sine.iteration[0] ),
    .X(_08920_));
 sky130_fd_sc_hd__or2_2 _16457_ (.A(_08899_),
    .B(_08920_),
    .X(_08921_));
 sky130_fd_sc_hd__buf_4 _16458_ (.A(_08895_),
    .X(_08922_));
 sky130_fd_sc_hd__a32o_1 _16459_ (.A1(_08903_),
    .A2(_08919_),
    .A3(_08921_),
    .B1(_08922_),
    .B2(_08910_),
    .X(_00941_));
 sky130_fd_sc_hd__mux2_1 _16460_ (.A0(_08919_),
    .A1(_08895_),
    .S(_08911_),
    .X(_08923_));
 sky130_fd_sc_hd__clkbuf_1 _16461_ (.A(_08923_),
    .X(_00940_));
 sky130_fd_sc_hd__or2_2 _16462_ (.A(\wfg_stim_sine_top.wfg_stim_sine.cur_state[0] ),
    .B(_08895_),
    .X(_08924_));
 sky130_fd_sc_hd__mux2_1 _16463_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.phase_in[15] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.quadrant[1] ),
    .S(_08924_),
    .X(_08925_));
 sky130_fd_sc_hd__clkbuf_1 _16464_ (.A(_08925_),
    .X(_00939_));
 sky130_fd_sc_hd__mux2_1 _16465_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.phase_in[14] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.quadrant[0] ),
    .S(_08924_),
    .X(_08926_));
 sky130_fd_sc_hd__clkbuf_1 _16466_ (.A(_08926_),
    .X(_00938_));
 sky130_fd_sc_hd__clkbuf_4 _16467_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[16] ),
    .X(_08927_));
 sky130_fd_sc_hd__clkbuf_4 _16468_ (.A(_08927_),
    .X(_08928_));
 sky130_fd_sc_hd__clkbuf_4 _16469_ (.A(_08928_),
    .X(_08929_));
 sky130_fd_sc_hd__clkbuf_4 _16470_ (.A(_08929_),
    .X(_08930_));
 sky130_fd_sc_hd__nor2_2 _16471_ (.A(_08930_),
    .B(_08906_),
    .Y(_08931_));
 sky130_fd_sc_hd__xnor2_1 _16472_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[15] ),
    .B(_08931_),
    .Y(_08932_));
 sky130_fd_sc_hd__nand2_1 _16473_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[14] ),
    .B(_08931_),
    .Y(_08933_));
 sky130_fd_sc_hd__or2_1 _16474_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[14] ),
    .B(_08931_),
    .X(_08934_));
 sky130_fd_sc_hd__nand2_1 _16475_ (.A(_08933_),
    .B(_08934_),
    .Y(_08935_));
 sky130_fd_sc_hd__or2_1 _16476_ (.A(\wfg_stim_sine_top.wfg_stim_sine.iteration[3] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.iteration[2] ),
    .X(_08936_));
 sky130_fd_sc_hd__buf_2 _16477_ (.A(_08936_),
    .X(_08937_));
 sky130_fd_sc_hd__nor2_1 _16478_ (.A(_08921_),
    .B(_08937_),
    .Y(_08938_));
 sky130_fd_sc_hd__nor3_1 _16479_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[13] ),
    .B(_08931_),
    .C(_08938_),
    .Y(_08939_));
 sky130_fd_sc_hd__nand2b_2 _16480_ (.A_N(_08899_),
    .B(_08901_),
    .Y(_08940_));
 sky130_fd_sc_hd__nor2_1 _16481_ (.A(_08937_),
    .B(_08940_),
    .Y(_08941_));
 sky130_fd_sc_hd__and2_1 _16482_ (.A(_08930_),
    .B(_08941_),
    .X(_08942_));
 sky130_fd_sc_hd__or2_1 _16483_ (.A(_08927_),
    .B(_08906_),
    .X(_08943_));
 sky130_fd_sc_hd__nor2_2 _16484_ (.A(_08900_),
    .B(_08936_),
    .Y(_08944_));
 sky130_fd_sc_hd__nor2_1 _16485_ (.A(_08943_),
    .B(_08944_),
    .Y(_08945_));
 sky130_fd_sc_hd__o21ai_1 _16486_ (.A1(_08942_),
    .A2(_08945_),
    .B1(\wfg_stim_sine_top.wfg_stim_sine.z[12] ),
    .Y(_08946_));
 sky130_fd_sc_hd__nor2_1 _16487_ (.A(_08906_),
    .B(_08938_),
    .Y(_08947_));
 sky130_fd_sc_hd__nor2_4 _16488_ (.A(\wfg_stim_sine_top.wfg_stim_sine.iteration[3] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.iteration[2] ),
    .Y(_08948_));
 sky130_fd_sc_hd__nand2_1 _16489_ (.A(_08900_),
    .B(_08948_),
    .Y(_08949_));
 sky130_fd_sc_hd__or2_1 _16490_ (.A(_08902_),
    .B(_08949_),
    .X(_08950_));
 sky130_fd_sc_hd__nand2_1 _16491_ (.A(_08929_),
    .B(_08950_),
    .Y(_08951_));
 sky130_fd_sc_hd__or2_1 _16492_ (.A(_08929_),
    .B(_08950_),
    .X(_08952_));
 sky130_fd_sc_hd__and3_1 _16493_ (.A(_08947_),
    .B(_08951_),
    .C(_08952_),
    .X(_08953_));
 sky130_fd_sc_hd__and2_1 _16494_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[11] ),
    .B(_08953_),
    .X(_08954_));
 sky130_fd_sc_hd__nor2_1 _16495_ (.A(_08943_),
    .B(_08938_),
    .Y(_08955_));
 sky130_fd_sc_hd__or2_1 _16496_ (.A(_08903_),
    .B(_08937_),
    .X(_08956_));
 sky130_fd_sc_hd__mux2_1 _16497_ (.A0(_08929_),
    .A1(_08955_),
    .S(_08956_),
    .X(_08957_));
 sky130_fd_sc_hd__nand2_1 _16498_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[10] ),
    .B(_08957_),
    .Y(_08958_));
 sky130_fd_sc_hd__inv_2 _16499_ (.A(\wfg_stim_sine_top.wfg_stim_sine.iteration[3] ),
    .Y(_08959_));
 sky130_fd_sc_hd__nand2_2 _16500_ (.A(_08959_),
    .B(_08904_),
    .Y(_08960_));
 sky130_fd_sc_hd__or3_1 _16501_ (.A(_08910_),
    .B(_08911_),
    .C(_08960_),
    .X(_08961_));
 sky130_fd_sc_hd__clkbuf_4 _16502_ (.A(_08959_),
    .X(_08962_));
 sky130_fd_sc_hd__nor2_1 _16503_ (.A(_08910_),
    .B(_08911_),
    .Y(_08963_));
 sky130_fd_sc_hd__a31o_1 _16504_ (.A1(_08962_),
    .A2(_08909_),
    .A3(_08963_),
    .B1(_08941_),
    .X(_08964_));
 sky130_fd_sc_hd__a22o_1 _16505_ (.A1(_08945_),
    .A2(_08961_),
    .B1(_08964_),
    .B2(_08929_),
    .X(_08965_));
 sky130_fd_sc_hd__nand2_1 _16506_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[9] ),
    .B(_08965_),
    .Y(_08966_));
 sky130_fd_sc_hd__clkbuf_4 _16507_ (.A(_08960_),
    .X(_08967_));
 sky130_fd_sc_hd__o21a_1 _16508_ (.A1(_08940_),
    .A2(_08967_),
    .B1(_08949_),
    .X(_08968_));
 sky130_fd_sc_hd__xnor2_1 _16509_ (.A(_08955_),
    .B(_08968_),
    .Y(_08969_));
 sky130_fd_sc_hd__and2_1 _16510_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[8] ),
    .B(_08969_),
    .X(_08970_));
 sky130_fd_sc_hd__or3b_1 _16511_ (.A(_08937_),
    .B(_08963_),
    .C_N(_08903_),
    .X(_08971_));
 sky130_fd_sc_hd__o21a_1 _16512_ (.A1(_08911_),
    .A2(_08967_),
    .B1(_08971_),
    .X(_08972_));
 sky130_fd_sc_hd__mux2_1 _16513_ (.A0(_08928_),
    .A1(_08955_),
    .S(_08972_),
    .X(_08973_));
 sky130_fd_sc_hd__and2_1 _16514_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[7] ),
    .B(_08973_),
    .X(_08974_));
 sky130_fd_sc_hd__and2_1 _16515_ (.A(_08959_),
    .B(\wfg_stim_sine_top.wfg_stim_sine.iteration[2] ),
    .X(_08975_));
 sky130_fd_sc_hd__clkbuf_4 _16516_ (.A(_08975_),
    .X(_08976_));
 sky130_fd_sc_hd__a21bo_1 _16517_ (.A1(_08911_),
    .A2(_08976_),
    .B1_N(_08971_),
    .X(_08977_));
 sky130_fd_sc_hd__mux2_1 _16518_ (.A0(_08955_),
    .A1(_08928_),
    .S(_08977_),
    .X(_08978_));
 sky130_fd_sc_hd__and2_1 _16519_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[6] ),
    .B(_08978_),
    .X(_08979_));
 sky130_fd_sc_hd__o211ai_2 _16520_ (.A1(_08903_),
    .A2(_08960_),
    .B1(_08950_),
    .C1(_08917_),
    .Y(_08980_));
 sky130_fd_sc_hd__inv_2 _16521_ (.A(\wfg_stim_sine_top.wfg_stim_sine.iteration[1] ),
    .Y(_08981_));
 sky130_fd_sc_hd__buf_4 _16522_ (.A(_08981_),
    .X(_08982_));
 sky130_fd_sc_hd__nor2_1 _16523_ (.A(_08982_),
    .B(_08911_),
    .Y(_08983_));
 sky130_fd_sc_hd__a22o_1 _16524_ (.A1(_08908_),
    .A2(_08963_),
    .B1(_08983_),
    .B2(_08905_),
    .X(_08984_));
 sky130_fd_sc_hd__nor2_1 _16525_ (.A(_08980_),
    .B(_08984_),
    .Y(_08985_));
 sky130_fd_sc_hd__o211ai_2 _16526_ (.A1(_08912_),
    .A2(_08982_),
    .B1(_08911_),
    .C1(_08905_),
    .Y(_08986_));
 sky130_fd_sc_hd__a21o_1 _16527_ (.A1(_08985_),
    .A2(_08986_),
    .B1(_08927_),
    .X(_08987_));
 sky130_fd_sc_hd__inv_2 _16528_ (.A(_08987_),
    .Y(_08988_));
 sky130_fd_sc_hd__or3_1 _16529_ (.A(_08959_),
    .B(_08908_),
    .C(_08921_),
    .X(_08989_));
 sky130_fd_sc_hd__o311a_1 _16530_ (.A1(_08982_),
    .A2(_08911_),
    .A3(_08967_),
    .B1(_08989_),
    .C1(_08971_),
    .X(_08990_));
 sky130_fd_sc_hd__mux2_1 _16531_ (.A0(_08928_),
    .A1(_08988_),
    .S(_08990_),
    .X(_08991_));
 sky130_fd_sc_hd__and2_1 _16532_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[5] ),
    .B(_08991_),
    .X(_08992_));
 sky130_fd_sc_hd__or3_1 _16533_ (.A(_08959_),
    .B(_08909_),
    .C(_08940_),
    .X(_08993_));
 sky130_fd_sc_hd__o211a_1 _16534_ (.A1(_08903_),
    .A2(_08967_),
    .B1(_08993_),
    .C1(_08949_),
    .X(_08994_));
 sky130_fd_sc_hd__nand2_1 _16535_ (.A(_08927_),
    .B(_08994_),
    .Y(_08995_));
 sky130_fd_sc_hd__or2_1 _16536_ (.A(_08927_),
    .B(_08994_),
    .X(_08996_));
 sky130_fd_sc_hd__and4_1 _16537_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[4] ),
    .B(_08947_),
    .C(_08995_),
    .D(_08996_),
    .X(_08997_));
 sky130_fd_sc_hd__o311a_1 _16538_ (.A1(_08909_),
    .A2(_08982_),
    .A3(_08911_),
    .B1(_08989_),
    .C1(_08961_),
    .X(_08998_));
 sky130_fd_sc_hd__xor2_1 _16539_ (.A(_08987_),
    .B(_08998_),
    .X(_08999_));
 sky130_fd_sc_hd__nand2_1 _16540_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[3] ),
    .B(_08999_),
    .Y(_09000_));
 sky130_fd_sc_hd__nor2_1 _16541_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[16] ),
    .B(_08985_),
    .Y(_09001_));
 sky130_fd_sc_hd__xnor2_1 _16542_ (.A(_08986_),
    .B(_09001_),
    .Y(_09002_));
 sky130_fd_sc_hd__and2_1 _16543_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[2] ),
    .B(_09002_),
    .X(_09003_));
 sky130_fd_sc_hd__inv_2 _16544_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[16] ),
    .Y(_09004_));
 sky130_fd_sc_hd__and2_1 _16545_ (.A(_09004_),
    .B(_08980_),
    .X(_09005_));
 sky130_fd_sc_hd__xor2_1 _16546_ (.A(_08984_),
    .B(_09005_),
    .X(_09006_));
 sky130_fd_sc_hd__and2_1 _16547_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[1] ),
    .B(_09006_),
    .X(_09007_));
 sky130_fd_sc_hd__and2_1 _16548_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[0] ),
    .B(_08980_),
    .X(_09008_));
 sky130_fd_sc_hd__nor2_1 _16549_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[1] ),
    .B(_09006_),
    .Y(_09009_));
 sky130_fd_sc_hd__nor2_1 _16550_ (.A(_09007_),
    .B(_09009_),
    .Y(_09010_));
 sky130_fd_sc_hd__and2_1 _16551_ (.A(_09008_),
    .B(_09010_),
    .X(_09011_));
 sky130_fd_sc_hd__nor2_1 _16552_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[2] ),
    .B(_09002_),
    .Y(_09012_));
 sky130_fd_sc_hd__or2_1 _16553_ (.A(_09003_),
    .B(_09012_),
    .X(_09013_));
 sky130_fd_sc_hd__o21ba_1 _16554_ (.A1(_09007_),
    .A2(_09011_),
    .B1_N(_09013_),
    .X(_09014_));
 sky130_fd_sc_hd__or2_1 _16555_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[3] ),
    .B(_08999_),
    .X(_09015_));
 sky130_fd_sc_hd__and2_1 _16556_ (.A(_09000_),
    .B(_09015_),
    .X(_09016_));
 sky130_fd_sc_hd__o21ai_1 _16557_ (.A1(_09003_),
    .A2(_09014_),
    .B1(_09016_),
    .Y(_09017_));
 sky130_fd_sc_hd__a31o_1 _16558_ (.A1(_08947_),
    .A2(_08995_),
    .A3(_08996_),
    .B1(\wfg_stim_sine_top.wfg_stim_sine.z[4] ),
    .X(_09018_));
 sky130_fd_sc_hd__or2b_1 _16559_ (.A(_08997_),
    .B_N(_09018_),
    .X(_09019_));
 sky130_fd_sc_hd__a21oi_1 _16560_ (.A1(_09000_),
    .A2(_09017_),
    .B1(_09019_),
    .Y(_09020_));
 sky130_fd_sc_hd__nor2_1 _16561_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[5] ),
    .B(_08991_),
    .Y(_09021_));
 sky130_fd_sc_hd__nor2_1 _16562_ (.A(_08992_),
    .B(_09021_),
    .Y(_09022_));
 sky130_fd_sc_hd__o21a_1 _16563_ (.A1(_08997_),
    .A2(_09020_),
    .B1(_09022_),
    .X(_09023_));
 sky130_fd_sc_hd__nor2_1 _16564_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[6] ),
    .B(_08978_),
    .Y(_09024_));
 sky130_fd_sc_hd__nor2_1 _16565_ (.A(_08979_),
    .B(_09024_),
    .Y(_09025_));
 sky130_fd_sc_hd__o21a_1 _16566_ (.A1(_08992_),
    .A2(_09023_),
    .B1(_09025_),
    .X(_09026_));
 sky130_fd_sc_hd__nor2_1 _16567_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[7] ),
    .B(_08973_),
    .Y(_09027_));
 sky130_fd_sc_hd__nor2_1 _16568_ (.A(_08974_),
    .B(_09027_),
    .Y(_09028_));
 sky130_fd_sc_hd__o21a_1 _16569_ (.A1(_08979_),
    .A2(_09026_),
    .B1(_09028_),
    .X(_09029_));
 sky130_fd_sc_hd__nor2_1 _16570_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[8] ),
    .B(_08969_),
    .Y(_09030_));
 sky130_fd_sc_hd__nor2_1 _16571_ (.A(_08970_),
    .B(_09030_),
    .Y(_09031_));
 sky130_fd_sc_hd__o21a_1 _16572_ (.A1(_08974_),
    .A2(_09029_),
    .B1(_09031_),
    .X(_09032_));
 sky130_fd_sc_hd__or2_1 _16573_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[9] ),
    .B(_08965_),
    .X(_09033_));
 sky130_fd_sc_hd__and2_1 _16574_ (.A(_08966_),
    .B(_09033_),
    .X(_09034_));
 sky130_fd_sc_hd__o21ai_1 _16575_ (.A1(_08970_),
    .A2(_09032_),
    .B1(_09034_),
    .Y(_09035_));
 sky130_fd_sc_hd__or2_1 _16576_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[10] ),
    .B(_08957_),
    .X(_09036_));
 sky130_fd_sc_hd__nand2_1 _16577_ (.A(_08958_),
    .B(_09036_),
    .Y(_09037_));
 sky130_fd_sc_hd__a21o_1 _16578_ (.A1(_08966_),
    .A2(_09035_),
    .B1(_09037_),
    .X(_09038_));
 sky130_fd_sc_hd__xnor2_1 _16579_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[11] ),
    .B(_08953_),
    .Y(_09039_));
 sky130_fd_sc_hd__a21oi_1 _16580_ (.A1(_08958_),
    .A2(_09038_),
    .B1(_09039_),
    .Y(_09040_));
 sky130_fd_sc_hd__or3_1 _16581_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[12] ),
    .B(_08942_),
    .C(_08945_),
    .X(_09041_));
 sky130_fd_sc_hd__o211ai_1 _16582_ (.A1(_08954_),
    .A2(_09040_),
    .B1(_08946_),
    .C1(_09041_),
    .Y(_09042_));
 sky130_fd_sc_hd__and2_1 _16583_ (.A(_08946_),
    .B(_09042_),
    .X(_09043_));
 sky130_fd_sc_hd__o21a_1 _16584_ (.A1(_08931_),
    .A2(_08938_),
    .B1(\wfg_stim_sine_top.wfg_stim_sine.z[13] ),
    .X(_09044_));
 sky130_fd_sc_hd__o21ba_1 _16585_ (.A1(_08939_),
    .A2(_09043_),
    .B1_N(_09044_),
    .X(_09045_));
 sky130_fd_sc_hd__or2_1 _16586_ (.A(_08935_),
    .B(_09045_),
    .X(_09046_));
 sky130_fd_sc_hd__or2_1 _16587_ (.A(_08932_),
    .B(_09046_),
    .X(_09047_));
 sky130_fd_sc_hd__nor2_1 _16588_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[15] ),
    .B(_08906_),
    .Y(_09048_));
 sky130_fd_sc_hd__o211a_1 _16589_ (.A1(_08930_),
    .A2(_09048_),
    .B1(_08933_),
    .C1(_08919_),
    .X(_09049_));
 sky130_fd_sc_hd__a22o_1 _16590_ (.A1(_08930_),
    .A2(_08896_),
    .B1(_09047_),
    .B2(_09049_),
    .X(_00937_));
 sky130_fd_sc_hd__buf_4 _16591_ (.A(_08918_),
    .X(_09050_));
 sky130_fd_sc_hd__nand3_1 _16592_ (.A(_08932_),
    .B(_08933_),
    .C(_09046_),
    .Y(_09051_));
 sky130_fd_sc_hd__a21o_1 _16593_ (.A1(_08933_),
    .A2(_09046_),
    .B1(_08932_),
    .X(_09052_));
 sky130_fd_sc_hd__a32o_1 _16594_ (.A1(_09050_),
    .A2(_09051_),
    .A3(_09052_),
    .B1(_08922_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.z[15] ),
    .X(_00936_));
 sky130_fd_sc_hd__nand2_1 _16595_ (.A(_08935_),
    .B(_09045_),
    .Y(_09053_));
 sky130_fd_sc_hd__buf_4 _16596_ (.A(_08895_),
    .X(_09054_));
 sky130_fd_sc_hd__a32o_1 _16597_ (.A1(_09050_),
    .A2(_09046_),
    .A3(_09053_),
    .B1(_09054_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.z[14] ),
    .X(_00935_));
 sky130_fd_sc_hd__clkbuf_4 _16598_ (.A(_08895_),
    .X(_09055_));
 sky130_fd_sc_hd__nor2_4 _16599_ (.A(\wfg_stim_sine_top.wfg_stim_sine.cur_state[0] ),
    .B(_08894_),
    .Y(_09056_));
 sky130_fd_sc_hd__clkbuf_4 _16600_ (.A(_09056_),
    .X(_09057_));
 sky130_fd_sc_hd__o21ai_1 _16601_ (.A1(_09044_),
    .A2(_08939_),
    .B1(_09043_),
    .Y(_09058_));
 sky130_fd_sc_hd__o311a_1 _16602_ (.A1(_09044_),
    .A2(_08939_),
    .A3(_09043_),
    .B1(_09058_),
    .C1(_08919_),
    .X(_09059_));
 sky130_fd_sc_hd__a221o_1 _16603_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.z[13] ),
    .A2(_09055_),
    .B1(_09057_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.phase_in[13] ),
    .C1(_09059_),
    .X(_00934_));
 sky130_fd_sc_hd__a211o_1 _16604_ (.A1(_08946_),
    .A2(_09041_),
    .B1(_08954_),
    .C1(_09040_),
    .X(_09060_));
 sky130_fd_sc_hd__and3_1 _16605_ (.A(_08918_),
    .B(_09042_),
    .C(_09060_),
    .X(_09061_));
 sky130_fd_sc_hd__a221o_1 _16606_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.z[12] ),
    .A2(_09055_),
    .B1(_09057_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.phase_in[12] ),
    .C1(_09061_),
    .X(_00933_));
 sky130_fd_sc_hd__and3_1 _16607_ (.A(_09039_),
    .B(_08958_),
    .C(_09038_),
    .X(_09062_));
 sky130_fd_sc_hd__or3_1 _16608_ (.A(_08915_),
    .B(_09040_),
    .C(_09062_),
    .X(_09063_));
 sky130_fd_sc_hd__a22oi_1 _16609_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.z[11] ),
    .A2(_08895_),
    .B1(_09056_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.phase_in[11] ),
    .Y(_09064_));
 sky130_fd_sc_hd__nand2_1 _16610_ (.A(_09063_),
    .B(_09064_),
    .Y(_00932_));
 sky130_fd_sc_hd__and3_1 _16611_ (.A(_09037_),
    .B(_08966_),
    .C(_09035_),
    .X(_09065_));
 sky130_fd_sc_hd__and3b_1 _16612_ (.A_N(_09065_),
    .B(_08918_),
    .C(_09038_),
    .X(_09066_));
 sky130_fd_sc_hd__a221o_1 _16613_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.z[10] ),
    .A2(_09055_),
    .B1(_09057_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.phase_in[10] ),
    .C1(_09066_),
    .X(_00931_));
 sky130_fd_sc_hd__or3_1 _16614_ (.A(_09034_),
    .B(_08970_),
    .C(_09032_),
    .X(_09067_));
 sky130_fd_sc_hd__and3_1 _16615_ (.A(_08918_),
    .B(_09035_),
    .C(_09067_),
    .X(_09068_));
 sky130_fd_sc_hd__a221o_1 _16616_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.z[9] ),
    .A2(_09055_),
    .B1(_09057_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.phase_in[9] ),
    .C1(_09068_),
    .X(_00930_));
 sky130_fd_sc_hd__nor2_1 _16617_ (.A(_08915_),
    .B(_09032_),
    .Y(_09069_));
 sky130_fd_sc_hd__o31a_1 _16618_ (.A1(_09031_),
    .A2(_08974_),
    .A3(_09029_),
    .B1(_09069_),
    .X(_09070_));
 sky130_fd_sc_hd__a221o_1 _16619_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.z[8] ),
    .A2(_09055_),
    .B1(_09057_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.phase_in[8] ),
    .C1(_09070_),
    .X(_00929_));
 sky130_fd_sc_hd__nor2_1 _16620_ (.A(_08915_),
    .B(_09029_),
    .Y(_09071_));
 sky130_fd_sc_hd__o31a_1 _16621_ (.A1(_09028_),
    .A2(_08979_),
    .A3(_09026_),
    .B1(_09071_),
    .X(_09072_));
 sky130_fd_sc_hd__a221o_1 _16622_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.z[7] ),
    .A2(_09055_),
    .B1(_09057_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.phase_in[7] ),
    .C1(_09072_),
    .X(_00928_));
 sky130_fd_sc_hd__nor2_1 _16623_ (.A(_08915_),
    .B(_09026_),
    .Y(_09073_));
 sky130_fd_sc_hd__o31a_1 _16624_ (.A1(_09025_),
    .A2(_08992_),
    .A3(_09023_),
    .B1(_09073_),
    .X(_09074_));
 sky130_fd_sc_hd__a221o_1 _16625_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.z[6] ),
    .A2(_09055_),
    .B1(_09057_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.phase_in[6] ),
    .C1(_09074_),
    .X(_00927_));
 sky130_fd_sc_hd__nor2_1 _16626_ (.A(_08898_),
    .B(_09023_),
    .Y(_09075_));
 sky130_fd_sc_hd__o31a_1 _16627_ (.A1(_09022_),
    .A2(_08997_),
    .A3(_09020_),
    .B1(_09075_),
    .X(_09076_));
 sky130_fd_sc_hd__a221o_1 _16628_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.z[5] ),
    .A2(_09055_),
    .B1(_09057_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.phase_in[5] ),
    .C1(_09076_),
    .X(_00926_));
 sky130_fd_sc_hd__and3_1 _16629_ (.A(_09019_),
    .B(_09000_),
    .C(_09017_),
    .X(_09077_));
 sky130_fd_sc_hd__or3_1 _16630_ (.A(_08915_),
    .B(_09020_),
    .C(_09077_),
    .X(_09078_));
 sky130_fd_sc_hd__a22oi_1 _16631_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.z[4] ),
    .A2(_08895_),
    .B1(_09056_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.phase_in[4] ),
    .Y(_09079_));
 sky130_fd_sc_hd__nand2_1 _16632_ (.A(_09078_),
    .B(_09079_),
    .Y(_00925_));
 sky130_fd_sc_hd__or3_1 _16633_ (.A(_09016_),
    .B(_09003_),
    .C(_09014_),
    .X(_09080_));
 sky130_fd_sc_hd__and3_1 _16634_ (.A(_08918_),
    .B(_09017_),
    .C(_09080_),
    .X(_09081_));
 sky130_fd_sc_hd__a221o_1 _16635_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.z[3] ),
    .A2(_09055_),
    .B1(_09057_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.phase_in[3] ),
    .C1(_09081_),
    .X(_00924_));
 sky130_fd_sc_hd__or3b_1 _16636_ (.A(_09007_),
    .B(_09011_),
    .C_N(_09013_),
    .X(_09082_));
 sky130_fd_sc_hd__and3b_1 _16637_ (.A_N(_09014_),
    .B(_09082_),
    .C(_08918_),
    .X(_09083_));
 sky130_fd_sc_hd__a221o_1 _16638_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.z[2] ),
    .A2(_09055_),
    .B1(_09057_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.phase_in[2] ),
    .C1(_09083_),
    .X(_00923_));
 sky130_fd_sc_hd__nor2_1 _16639_ (.A(_08915_),
    .B(_09011_),
    .Y(_09084_));
 sky130_fd_sc_hd__o21a_1 _16640_ (.A1(_09008_),
    .A2(_09010_),
    .B1(_09084_),
    .X(_09085_));
 sky130_fd_sc_hd__a221o_1 _16641_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.z[1] ),
    .A2(_08895_),
    .B1(_09056_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.phase_in[1] ),
    .C1(_09085_),
    .X(_00922_));
 sky130_fd_sc_hd__buf_4 _16642_ (.A(_08897_),
    .X(_09086_));
 sky130_fd_sc_hd__nor2_1 _16643_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[0] ),
    .B(_08980_),
    .Y(_09087_));
 sky130_fd_sc_hd__o21ai_1 _16644_ (.A1(_09008_),
    .A2(_09087_),
    .B1(_08919_),
    .Y(_09088_));
 sky130_fd_sc_hd__o221a_1 _16645_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.z[0] ),
    .A2(_09086_),
    .B1(_08924_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.phase_in[0] ),
    .C1(_09088_),
    .X(_00921_));
 sky130_fd_sc_hd__mux2_1 _16646_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[15] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.x[16] ),
    .S(_08920_),
    .X(_09089_));
 sky130_fd_sc_hd__mux2_1 _16647_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[16] ),
    .A1(_09089_),
    .S(_08982_),
    .X(_09090_));
 sky130_fd_sc_hd__or2b_1 _16648_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[16] ),
    .B_N(_08904_),
    .X(_09091_));
 sky130_fd_sc_hd__o21a_1 _16649_ (.A1(_08909_),
    .A2(_09090_),
    .B1(_09091_),
    .X(_09092_));
 sky130_fd_sc_hd__or2_1 _16650_ (.A(_08962_),
    .B(\wfg_stim_sine_top.wfg_stim_sine.x[16] ),
    .X(_09093_));
 sky130_fd_sc_hd__clkbuf_2 _16651_ (.A(_09093_),
    .X(_09094_));
 sky130_fd_sc_hd__o21ai_1 _16652_ (.A1(_08913_),
    .A2(_09092_),
    .B1(_09094_),
    .Y(_09095_));
 sky130_fd_sc_hd__mux2_1 _16653_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[14] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.x[15] ),
    .S(_08901_),
    .X(_09096_));
 sky130_fd_sc_hd__mux2_1 _16654_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[16] ),
    .A1(_09096_),
    .S(_08981_),
    .X(_09097_));
 sky130_fd_sc_hd__o21a_1 _16655_ (.A1(_08909_),
    .A2(_09097_),
    .B1(_09091_),
    .X(_09098_));
 sky130_fd_sc_hd__o21ai_1 _16656_ (.A1(_08913_),
    .A2(_09098_),
    .B1(_09094_),
    .Y(_09099_));
 sky130_fd_sc_hd__mux2_1 _16657_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[13] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.x[14] ),
    .S(_08920_),
    .X(_09100_));
 sky130_fd_sc_hd__mux2_1 _16658_ (.A0(_09089_),
    .A1(_09100_),
    .S(_08981_),
    .X(_09101_));
 sky130_fd_sc_hd__o21ai_1 _16659_ (.A1(_08908_),
    .A2(_09101_),
    .B1(_09091_),
    .Y(_09102_));
 sky130_fd_sc_hd__a21boi_1 _16660_ (.A1(_08962_),
    .A2(_09102_),
    .B1_N(_09094_),
    .Y(_09103_));
 sky130_fd_sc_hd__inv_2 _16661_ (.A(_09103_),
    .Y(_09104_));
 sky130_fd_sc_hd__mux2_1 _16662_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[11] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.x[12] ),
    .S(_08920_),
    .X(_09105_));
 sky130_fd_sc_hd__mux2_1 _16663_ (.A0(_09105_),
    .A1(_09100_),
    .S(_08910_),
    .X(_09106_));
 sky130_fd_sc_hd__mux2_1 _16664_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[9] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.x[10] ),
    .S(_08920_),
    .X(_09107_));
 sky130_fd_sc_hd__mux2_1 _16665_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[7] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.x[8] ),
    .S(_08902_),
    .X(_09108_));
 sky130_fd_sc_hd__mux2_1 _16666_ (.A0(_09107_),
    .A1(_09108_),
    .S(_08982_),
    .X(_09109_));
 sky130_fd_sc_hd__or2_1 _16667_ (.A(_08937_),
    .B(_09109_),
    .X(_09110_));
 sky130_fd_sc_hd__o221a_1 _16668_ (.A1(_08959_),
    .A2(_09092_),
    .B1(_09106_),
    .B2(_08967_),
    .C1(_09110_),
    .X(_09111_));
 sky130_fd_sc_hd__mux2_1 _16669_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[8] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.x[9] ),
    .S(_08920_),
    .X(_09112_));
 sky130_fd_sc_hd__mux2_1 _16670_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[10] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.x[11] ),
    .S(_08901_),
    .X(_09113_));
 sky130_fd_sc_hd__mux2_1 _16671_ (.A0(_09112_),
    .A1(_09113_),
    .S(_08899_),
    .X(_09114_));
 sky130_fd_sc_hd__mux2_1 _16672_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[12] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.x[13] ),
    .S(_08920_),
    .X(_09115_));
 sky130_fd_sc_hd__mux2_1 _16673_ (.A0(_09115_),
    .A1(_09096_),
    .S(_08899_),
    .X(_09116_));
 sky130_fd_sc_hd__mux2_1 _16674_ (.A0(_09114_),
    .A1(_09116_),
    .S(_08904_),
    .X(_09117_));
 sky130_fd_sc_hd__mux2_1 _16675_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[2] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.x[3] ),
    .S(_08920_),
    .X(_09118_));
 sky130_fd_sc_hd__or3_1 _16676_ (.A(_08899_),
    .B(_08902_),
    .C(\wfg_stim_sine_top.wfg_stim_sine.x[0] ),
    .X(_09119_));
 sky130_fd_sc_hd__o221a_1 _16677_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.x[1] ),
    .A2(_08940_),
    .B1(_09118_),
    .B2(_08981_),
    .C1(_09119_),
    .X(_09120_));
 sky130_fd_sc_hd__mux2_1 _16678_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[4] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.x[5] ),
    .S(_08920_),
    .X(_09121_));
 sky130_fd_sc_hd__mux2_1 _16679_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[6] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.x[7] ),
    .S(_08920_),
    .X(_09122_));
 sky130_fd_sc_hd__mux2_1 _16680_ (.A0(_09121_),
    .A1(_09122_),
    .S(_08900_),
    .X(_09123_));
 sky130_fd_sc_hd__a22o_1 _16681_ (.A1(_08948_),
    .A2(_09120_),
    .B1(_09123_),
    .B2(_08976_),
    .X(_09124_));
 sky130_fd_sc_hd__a21oi_2 _16682_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.iteration[3] ),
    .A2(_09117_),
    .B1(_09124_),
    .Y(_09125_));
 sky130_fd_sc_hd__mux2_1 _16683_ (.A0(_09107_),
    .A1(_09105_),
    .S(_08900_),
    .X(_09126_));
 sky130_fd_sc_hd__mux2_1 _16684_ (.A0(_09126_),
    .A1(_09101_),
    .S(_08904_),
    .X(_09127_));
 sky130_fd_sc_hd__mux2_1 _16685_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[5] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.x[6] ),
    .S(_08902_),
    .X(_09128_));
 sky130_fd_sc_hd__mux2_1 _16686_ (.A0(_09128_),
    .A1(_09108_),
    .S(_08900_),
    .X(_09129_));
 sky130_fd_sc_hd__mux2_1 _16687_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[3] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.x[4] ),
    .S(_08902_),
    .X(_09130_));
 sky130_fd_sc_hd__o221a_1 _16688_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.x[1] ),
    .A2(_08921_),
    .B1(_08940_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.x[2] ),
    .C1(_08948_),
    .X(_09131_));
 sky130_fd_sc_hd__o21a_1 _16689_ (.A1(_08982_),
    .A2(_09130_),
    .B1(_09131_),
    .X(_09132_));
 sky130_fd_sc_hd__a221oi_2 _16690_ (.A1(_08912_),
    .A2(_09127_),
    .B1(_09129_),
    .B2(_08976_),
    .C1(_09132_),
    .Y(_09133_));
 sky130_fd_sc_hd__and2_1 _16691_ (.A(_09125_),
    .B(_09133_),
    .X(_09134_));
 sky130_fd_sc_hd__mux2_1 _16692_ (.A0(_09113_),
    .A1(_09115_),
    .S(_08910_),
    .X(_09135_));
 sky130_fd_sc_hd__or2b_1 _16693_ (.A(_09097_),
    .B_N(_08904_),
    .X(_09136_));
 sky130_fd_sc_hd__o21ai_2 _16694_ (.A1(_08908_),
    .A2(_09135_),
    .B1(_09136_),
    .Y(_09137_));
 sky130_fd_sc_hd__mux2_1 _16695_ (.A0(_09112_),
    .A1(_09122_),
    .S(_08982_),
    .X(_09138_));
 sky130_fd_sc_hd__and3_1 _16696_ (.A(_08910_),
    .B(_08948_),
    .C(_09121_),
    .X(_09139_));
 sky130_fd_sc_hd__a221o_1 _16697_ (.A1(_08944_),
    .A2(_09118_),
    .B1(_09138_),
    .B2(_08976_),
    .C1(_09139_),
    .X(_09140_));
 sky130_fd_sc_hd__o21ba_1 _16698_ (.A1(_08959_),
    .A2(_09137_),
    .B1_N(_09140_),
    .X(_09141_));
 sky130_fd_sc_hd__and2_1 _16699_ (.A(_09134_),
    .B(_09141_),
    .X(_09142_));
 sky130_fd_sc_hd__mux2_1 _16700_ (.A0(_09106_),
    .A1(_09090_),
    .S(_08908_),
    .X(_09143_));
 sky130_fd_sc_hd__and3_1 _16701_ (.A(_08910_),
    .B(_08948_),
    .C(_09128_),
    .X(_09144_));
 sky130_fd_sc_hd__a221o_1 _16702_ (.A1(_08944_),
    .A2(_09130_),
    .B1(_09109_),
    .B2(_08976_),
    .C1(_09144_),
    .X(_09145_));
 sky130_fd_sc_hd__a21oi_2 _16703_ (.A1(_08912_),
    .A2(_09143_),
    .B1(_09145_),
    .Y(_09146_));
 sky130_fd_sc_hd__o21a_1 _16704_ (.A1(_08908_),
    .A2(_09116_),
    .B1(_09091_),
    .X(_09147_));
 sky130_fd_sc_hd__or2_1 _16705_ (.A(_08936_),
    .B(_09123_),
    .X(_09148_));
 sky130_fd_sc_hd__o221a_1 _16706_ (.A1(_08960_),
    .A2(_09114_),
    .B1(_09147_),
    .B2(_08959_),
    .C1(_09148_),
    .X(_09149_));
 sky130_fd_sc_hd__inv_2 _16707_ (.A(_09149_),
    .Y(_09150_));
 sky130_fd_sc_hd__o22a_1 _16708_ (.A1(_08960_),
    .A2(_09126_),
    .B1(_09129_),
    .B2(_08936_),
    .X(_09151_));
 sky130_fd_sc_hd__a21bo_1 _16709_ (.A1(_08912_),
    .A2(_09102_),
    .B1_N(_09151_),
    .X(_09152_));
 sky130_fd_sc_hd__and4_1 _16710_ (.A(_09142_),
    .B(_09146_),
    .C(_09150_),
    .D(_09152_),
    .X(_09153_));
 sky130_fd_sc_hd__o22a_1 _16711_ (.A1(_08967_),
    .A2(_09135_),
    .B1(_09138_),
    .B2(_08937_),
    .X(_09154_));
 sky130_fd_sc_hd__o21ai_2 _16712_ (.A1(_08962_),
    .A2(_09098_),
    .B1(_09154_),
    .Y(_09155_));
 sky130_fd_sc_hd__and3b_1 _16713_ (.A_N(_09111_),
    .B(_09153_),
    .C(_09155_),
    .X(_09156_));
 sky130_fd_sc_hd__o21ai_2 _16714_ (.A1(_08912_),
    .A2(_09117_),
    .B1(_09094_),
    .Y(_09157_));
 sky130_fd_sc_hd__o21ai_1 _16715_ (.A1(_08913_),
    .A2(_09127_),
    .B1(_09094_),
    .Y(_09158_));
 sky130_fd_sc_hd__a21bo_1 _16716_ (.A1(_08962_),
    .A2(_09137_),
    .B1_N(_09094_),
    .X(_09159_));
 sky130_fd_sc_hd__and4_1 _16717_ (.A(_09156_),
    .B(_09157_),
    .C(_09158_),
    .D(_09159_),
    .X(_09160_));
 sky130_fd_sc_hd__o21ai_1 _16718_ (.A1(_08913_),
    .A2(_09143_),
    .B1(_09094_),
    .Y(_09161_));
 sky130_fd_sc_hd__o21ai_1 _16719_ (.A1(_08913_),
    .A2(_09147_),
    .B1(_09094_),
    .Y(_09162_));
 sky130_fd_sc_hd__a31o_1 _16720_ (.A1(_09160_),
    .A2(_09161_),
    .A3(_09162_),
    .B1(_08930_),
    .X(_09163_));
 sky130_fd_sc_hd__o21a_1 _16721_ (.A1(_08930_),
    .A2(_09104_),
    .B1(_09163_),
    .X(_09164_));
 sky130_fd_sc_hd__o21a_1 _16722_ (.A1(_08930_),
    .A2(_09099_),
    .B1(_09164_),
    .X(_09165_));
 sky130_fd_sc_hd__xnor2_1 _16723_ (.A(_09095_),
    .B(_09165_),
    .Y(_09166_));
 sky130_fd_sc_hd__nand2_1 _16724_ (.A(\wfg_stim_sine_top.wfg_stim_sine.y[15] ),
    .B(_09166_),
    .Y(_09167_));
 sky130_fd_sc_hd__xnor2_1 _16725_ (.A(_09099_),
    .B(_09164_),
    .Y(_09168_));
 sky130_fd_sc_hd__nand2_1 _16726_ (.A(\wfg_stim_sine_top.wfg_stim_sine.y[14] ),
    .B(_09168_),
    .Y(_09169_));
 sky130_fd_sc_hd__or2_1 _16727_ (.A(\wfg_stim_sine_top.wfg_stim_sine.y[14] ),
    .B(_09168_),
    .X(_09170_));
 sky130_fd_sc_hd__and2_1 _16728_ (.A(_09169_),
    .B(_09170_),
    .X(_09171_));
 sky130_fd_sc_hd__xnor2_1 _16729_ (.A(_09104_),
    .B(_09163_),
    .Y(_09172_));
 sky130_fd_sc_hd__and2_1 _16730_ (.A(\wfg_stim_sine_top.wfg_stim_sine.y[13] ),
    .B(_09172_),
    .X(_09173_));
 sky130_fd_sc_hd__nor2_1 _16731_ (.A(\wfg_stim_sine_top.wfg_stim_sine.y[13] ),
    .B(_09172_),
    .Y(_09174_));
 sky130_fd_sc_hd__nor2_1 _16732_ (.A(_09173_),
    .B(_09174_),
    .Y(_09175_));
 sky130_fd_sc_hd__a21o_1 _16733_ (.A1(_09160_),
    .A2(_09161_),
    .B1(_08929_),
    .X(_09176_));
 sky130_fd_sc_hd__xnor2_1 _16734_ (.A(_09162_),
    .B(_09176_),
    .Y(_09177_));
 sky130_fd_sc_hd__nor2_1 _16735_ (.A(_08929_),
    .B(_09160_),
    .Y(_09178_));
 sky130_fd_sc_hd__xnor2_1 _16736_ (.A(_09161_),
    .B(_09178_),
    .Y(_09179_));
 sky130_fd_sc_hd__and2b_1 _16737_ (.A_N(_09179_),
    .B(\wfg_stim_sine_top.wfg_stim_sine.y[11] ),
    .X(_09180_));
 sky130_fd_sc_hd__a31o_1 _16738_ (.A1(_09156_),
    .A2(_09157_),
    .A3(_09158_),
    .B1(_08929_),
    .X(_09181_));
 sky130_fd_sc_hd__xor2_1 _16739_ (.A(_09159_),
    .B(_09181_),
    .X(_09182_));
 sky130_fd_sc_hd__and2b_1 _16740_ (.A_N(_09182_),
    .B(\wfg_stim_sine_top.wfg_stim_sine.y[10] ),
    .X(_09183_));
 sky130_fd_sc_hd__a21o_1 _16741_ (.A1(_09156_),
    .A2(_09157_),
    .B1(_08928_),
    .X(_09184_));
 sky130_fd_sc_hd__xor2_1 _16742_ (.A(_09158_),
    .B(_09184_),
    .X(_09185_));
 sky130_fd_sc_hd__and2b_1 _16743_ (.A_N(_09185_),
    .B(\wfg_stim_sine_top.wfg_stim_sine.y[9] ),
    .X(_09186_));
 sky130_fd_sc_hd__or2_1 _16744_ (.A(_08928_),
    .B(_09156_),
    .X(_09187_));
 sky130_fd_sc_hd__xor2_1 _16745_ (.A(_09157_),
    .B(_09187_),
    .X(_09188_));
 sky130_fd_sc_hd__and2b_1 _16746_ (.A_N(_09188_),
    .B(\wfg_stim_sine_top.wfg_stim_sine.y[8] ),
    .X(_09189_));
 sky130_fd_sc_hd__a21oi_1 _16747_ (.A1(_09153_),
    .A2(_09155_),
    .B1(_08928_),
    .Y(_09190_));
 sky130_fd_sc_hd__xnor2_1 _16748_ (.A(_09111_),
    .B(_09190_),
    .Y(_09191_));
 sky130_fd_sc_hd__nand2_1 _16749_ (.A(\wfg_stim_sine_top.wfg_stim_sine.y[7] ),
    .B(_09191_),
    .Y(_09192_));
 sky130_fd_sc_hd__or2_1 _16750_ (.A(_08927_),
    .B(_09153_),
    .X(_09193_));
 sky130_fd_sc_hd__xnor2_1 _16751_ (.A(_09155_),
    .B(_09193_),
    .Y(_09194_));
 sky130_fd_sc_hd__nand2_1 _16752_ (.A(\wfg_stim_sine_top.wfg_stim_sine.y[6] ),
    .B(_09194_),
    .Y(_09195_));
 sky130_fd_sc_hd__a31o_1 _16753_ (.A1(_09142_),
    .A2(_09146_),
    .A3(_09150_),
    .B1(_08927_),
    .X(_09196_));
 sky130_fd_sc_hd__xnor2_1 _16754_ (.A(_09152_),
    .B(_09196_),
    .Y(_09197_));
 sky130_fd_sc_hd__and2_1 _16755_ (.A(\wfg_stim_sine_top.wfg_stim_sine.y[5] ),
    .B(_09197_),
    .X(_09198_));
 sky130_fd_sc_hd__a21oi_1 _16756_ (.A1(_09142_),
    .A2(_09146_),
    .B1(_08927_),
    .Y(_09199_));
 sky130_fd_sc_hd__xnor2_1 _16757_ (.A(_09149_),
    .B(_09199_),
    .Y(_09200_));
 sky130_fd_sc_hd__and2_1 _16758_ (.A(\wfg_stim_sine_top.wfg_stim_sine.y[4] ),
    .B(_09200_),
    .X(_09201_));
 sky130_fd_sc_hd__inv_2 _16759_ (.A(\wfg_stim_sine_top.wfg_stim_sine.y[3] ),
    .Y(_09202_));
 sky130_fd_sc_hd__nor2_1 _16760_ (.A(_08927_),
    .B(_09142_),
    .Y(_09203_));
 sky130_fd_sc_hd__xnor2_1 _16761_ (.A(_09146_),
    .B(_09203_),
    .Y(_09204_));
 sky130_fd_sc_hd__nor2_1 _16762_ (.A(_09202_),
    .B(_09204_),
    .Y(_09205_));
 sky130_fd_sc_hd__inv_2 _16763_ (.A(\wfg_stim_sine_top.wfg_stim_sine.y[2] ),
    .Y(_09206_));
 sky130_fd_sc_hd__or2_1 _16764_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[16] ),
    .B(_09134_),
    .X(_09207_));
 sky130_fd_sc_hd__xor2_1 _16765_ (.A(_09141_),
    .B(_09207_),
    .X(_09208_));
 sky130_fd_sc_hd__nor2_1 _16766_ (.A(_09206_),
    .B(_09208_),
    .Y(_09209_));
 sky130_fd_sc_hd__or2_1 _16767_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[16] ),
    .B(_09125_),
    .X(_09210_));
 sky130_fd_sc_hd__xnor2_1 _16768_ (.A(_09133_),
    .B(_09210_),
    .Y(_09211_));
 sky130_fd_sc_hd__nand2_1 _16769_ (.A(\wfg_stim_sine_top.wfg_stim_sine.y[1] ),
    .B(_09211_),
    .Y(_09212_));
 sky130_fd_sc_hd__nor2_1 _16770_ (.A(\wfg_stim_sine_top.wfg_stim_sine.y[0] ),
    .B(_09125_),
    .Y(_09213_));
 sky130_fd_sc_hd__xnor2_1 _16771_ (.A(\wfg_stim_sine_top.wfg_stim_sine.y[1] ),
    .B(_09211_),
    .Y(_09214_));
 sky130_fd_sc_hd__or2_1 _16772_ (.A(_09213_),
    .B(_09214_),
    .X(_09215_));
 sky130_fd_sc_hd__xnor2_1 _16773_ (.A(_09206_),
    .B(_09208_),
    .Y(_09216_));
 sky130_fd_sc_hd__a21oi_1 _16774_ (.A1(_09212_),
    .A2(_09215_),
    .B1(_09216_),
    .Y(_09217_));
 sky130_fd_sc_hd__xnor2_1 _16775_ (.A(_09202_),
    .B(_09204_),
    .Y(_09218_));
 sky130_fd_sc_hd__o21ba_1 _16776_ (.A1(_09209_),
    .A2(_09217_),
    .B1_N(_09218_),
    .X(_09219_));
 sky130_fd_sc_hd__xor2_1 _16777_ (.A(\wfg_stim_sine_top.wfg_stim_sine.y[4] ),
    .B(_09200_),
    .X(_09220_));
 sky130_fd_sc_hd__o21a_1 _16778_ (.A1(_09205_),
    .A2(_09219_),
    .B1(_09220_),
    .X(_09221_));
 sky130_fd_sc_hd__nor2_1 _16779_ (.A(\wfg_stim_sine_top.wfg_stim_sine.y[5] ),
    .B(_09197_),
    .Y(_09222_));
 sky130_fd_sc_hd__nor2_1 _16780_ (.A(_09198_),
    .B(_09222_),
    .Y(_09223_));
 sky130_fd_sc_hd__o21a_1 _16781_ (.A1(_09201_),
    .A2(_09221_),
    .B1(_09223_),
    .X(_09224_));
 sky130_fd_sc_hd__or2_1 _16782_ (.A(\wfg_stim_sine_top.wfg_stim_sine.y[6] ),
    .B(_09194_),
    .X(_09225_));
 sky130_fd_sc_hd__and2_1 _16783_ (.A(_09195_),
    .B(_09225_),
    .X(_09226_));
 sky130_fd_sc_hd__o21ai_1 _16784_ (.A1(_09198_),
    .A2(_09224_),
    .B1(_09226_),
    .Y(_09227_));
 sky130_fd_sc_hd__or2_1 _16785_ (.A(\wfg_stim_sine_top.wfg_stim_sine.y[7] ),
    .B(_09191_),
    .X(_09228_));
 sky130_fd_sc_hd__and2_1 _16786_ (.A(_09192_),
    .B(_09228_),
    .X(_09229_));
 sky130_fd_sc_hd__a21bo_1 _16787_ (.A1(_09195_),
    .A2(_09227_),
    .B1_N(_09229_),
    .X(_09230_));
 sky130_fd_sc_hd__and2b_1 _16788_ (.A_N(\wfg_stim_sine_top.wfg_stim_sine.y[8] ),
    .B(_09188_),
    .X(_09231_));
 sky130_fd_sc_hd__nor2_1 _16789_ (.A(_09189_),
    .B(_09231_),
    .Y(_09232_));
 sky130_fd_sc_hd__a21boi_1 _16790_ (.A1(_09192_),
    .A2(_09230_),
    .B1_N(_09232_),
    .Y(_09233_));
 sky130_fd_sc_hd__and2b_1 _16791_ (.A_N(\wfg_stim_sine_top.wfg_stim_sine.y[9] ),
    .B(_09185_),
    .X(_09234_));
 sky130_fd_sc_hd__nor2_1 _16792_ (.A(_09186_),
    .B(_09234_),
    .Y(_09235_));
 sky130_fd_sc_hd__o21a_1 _16793_ (.A1(_09189_),
    .A2(_09233_),
    .B1(_09235_),
    .X(_09236_));
 sky130_fd_sc_hd__and2b_1 _16794_ (.A_N(\wfg_stim_sine_top.wfg_stim_sine.y[10] ),
    .B(_09182_),
    .X(_09237_));
 sky130_fd_sc_hd__nor2_1 _16795_ (.A(_09183_),
    .B(_09237_),
    .Y(_09238_));
 sky130_fd_sc_hd__o21a_1 _16796_ (.A1(_09186_),
    .A2(_09236_),
    .B1(_09238_),
    .X(_09239_));
 sky130_fd_sc_hd__and2b_1 _16797_ (.A_N(\wfg_stim_sine_top.wfg_stim_sine.y[11] ),
    .B(_09179_),
    .X(_09240_));
 sky130_fd_sc_hd__nor2_1 _16798_ (.A(_09180_),
    .B(_09240_),
    .Y(_09241_));
 sky130_fd_sc_hd__o21a_1 _16799_ (.A1(_09183_),
    .A2(_09239_),
    .B1(_09241_),
    .X(_09242_));
 sky130_fd_sc_hd__xor2_1 _16800_ (.A(\wfg_stim_sine_top.wfg_stim_sine.y[12] ),
    .B(_09177_),
    .X(_09243_));
 sky130_fd_sc_hd__o21ai_1 _16801_ (.A1(_09180_),
    .A2(_09242_),
    .B1(_09243_),
    .Y(_09244_));
 sky130_fd_sc_hd__a21bo_1 _16802_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[12] ),
    .A2(_09177_),
    .B1_N(_09244_),
    .X(_09245_));
 sky130_fd_sc_hd__a21o_1 _16803_ (.A1(_09175_),
    .A2(_09245_),
    .B1(_09173_),
    .X(_09246_));
 sky130_fd_sc_hd__nand2_1 _16804_ (.A(_09171_),
    .B(_09246_),
    .Y(_09247_));
 sky130_fd_sc_hd__or2_1 _16805_ (.A(\wfg_stim_sine_top.wfg_stim_sine.y[15] ),
    .B(_09166_),
    .X(_09248_));
 sky130_fd_sc_hd__nand2_1 _16806_ (.A(_09167_),
    .B(_09248_),
    .Y(_09249_));
 sky130_fd_sc_hd__a21o_1 _16807_ (.A1(_09169_),
    .A2(_09247_),
    .B1(_09249_),
    .X(_09250_));
 sky130_fd_sc_hd__xor2_1 _16808_ (.A(\wfg_stim_sine_top.wfg_stim_sine.y[16] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.x[16] ),
    .X(_09251_));
 sky130_fd_sc_hd__o21a_1 _16809_ (.A1(_08930_),
    .A2(_09095_),
    .B1(_09165_),
    .X(_09252_));
 sky130_fd_sc_hd__xnor2_1 _16810_ (.A(_09251_),
    .B(_09252_),
    .Y(_09253_));
 sky130_fd_sc_hd__a21oi_1 _16811_ (.A1(_09167_),
    .A2(_09250_),
    .B1(_09253_),
    .Y(_09254_));
 sky130_fd_sc_hd__a31o_1 _16812_ (.A1(_09167_),
    .A2(_09250_),
    .A3(_09253_),
    .B1(_08915_),
    .X(_09255_));
 sky130_fd_sc_hd__a2bb2o_1 _16813_ (.A1_N(_09254_),
    .A2_N(_09255_),
    .B1(\wfg_stim_sine_top.wfg_stim_sine.y[16] ),
    .B2(_08896_),
    .X(_00920_));
 sky130_fd_sc_hd__nand3_1 _16814_ (.A(_09249_),
    .B(_09169_),
    .C(_09247_),
    .Y(_09256_));
 sky130_fd_sc_hd__a32o_1 _16815_ (.A1(_09050_),
    .A2(_09250_),
    .A3(_09256_),
    .B1(_09054_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.y[15] ),
    .X(_00919_));
 sky130_fd_sc_hd__xor2_1 _16816_ (.A(_09171_),
    .B(_09246_),
    .X(_09257_));
 sky130_fd_sc_hd__a22o_1 _16817_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[14] ),
    .A2(_08896_),
    .B1(_09050_),
    .B2(_09257_),
    .X(_00918_));
 sky130_fd_sc_hd__xor2_1 _16818_ (.A(_09175_),
    .B(_09245_),
    .X(_09258_));
 sky130_fd_sc_hd__a22o_1 _16819_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[13] ),
    .A2(_08896_),
    .B1(_09050_),
    .B2(_09258_),
    .X(_00917_));
 sky130_fd_sc_hd__or3_1 _16820_ (.A(_09243_),
    .B(_09180_),
    .C(_09242_),
    .X(_09259_));
 sky130_fd_sc_hd__a32o_1 _16821_ (.A1(_09050_),
    .A2(_09244_),
    .A3(_09259_),
    .B1(_09054_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.y[12] ),
    .X(_00916_));
 sky130_fd_sc_hd__or3_1 _16822_ (.A(_09241_),
    .B(_09183_),
    .C(_09239_),
    .X(_09260_));
 sky130_fd_sc_hd__buf_4 _16823_ (.A(_08915_),
    .X(_09261_));
 sky130_fd_sc_hd__nor2_1 _16824_ (.A(_09261_),
    .B(_09242_),
    .Y(_09262_));
 sky130_fd_sc_hd__a22o_1 _16825_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[11] ),
    .A2(_08896_),
    .B1(_09260_),
    .B2(_09262_),
    .X(_00915_));
 sky130_fd_sc_hd__or3_1 _16826_ (.A(_09238_),
    .B(_09186_),
    .C(_09236_),
    .X(_09263_));
 sky130_fd_sc_hd__nor2_1 _16827_ (.A(_09261_),
    .B(_09239_),
    .Y(_09264_));
 sky130_fd_sc_hd__a22o_1 _16828_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[10] ),
    .A2(_08896_),
    .B1(_09263_),
    .B2(_09264_),
    .X(_00914_));
 sky130_fd_sc_hd__or3_1 _16829_ (.A(_09235_),
    .B(_09189_),
    .C(_09233_),
    .X(_09265_));
 sky130_fd_sc_hd__nor2_1 _16830_ (.A(_09261_),
    .B(_09236_),
    .Y(_09266_));
 sky130_fd_sc_hd__a22o_1 _16831_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[9] ),
    .A2(_08896_),
    .B1(_09265_),
    .B2(_09266_),
    .X(_00913_));
 sky130_fd_sc_hd__nand3b_1 _16832_ (.A_N(_09232_),
    .B(_09192_),
    .C(_09230_),
    .Y(_09267_));
 sky130_fd_sc_hd__nor2_1 _16833_ (.A(_09261_),
    .B(_09233_),
    .Y(_09268_));
 sky130_fd_sc_hd__a22o_1 _16834_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[8] ),
    .A2(_08922_),
    .B1(_09267_),
    .B2(_09268_),
    .X(_00912_));
 sky130_fd_sc_hd__nand3b_1 _16835_ (.A_N(_09229_),
    .B(_09195_),
    .C(_09227_),
    .Y(_09269_));
 sky130_fd_sc_hd__a32o_1 _16836_ (.A1(_09050_),
    .A2(_09230_),
    .A3(_09269_),
    .B1(_09054_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.y[7] ),
    .X(_00911_));
 sky130_fd_sc_hd__or3_1 _16837_ (.A(_09226_),
    .B(_09198_),
    .C(_09224_),
    .X(_09270_));
 sky130_fd_sc_hd__a32o_1 _16838_ (.A1(_09050_),
    .A2(_09227_),
    .A3(_09270_),
    .B1(_09054_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.y[6] ),
    .X(_00910_));
 sky130_fd_sc_hd__or3_1 _16839_ (.A(_09223_),
    .B(_09201_),
    .C(_09221_),
    .X(_09271_));
 sky130_fd_sc_hd__nor2_1 _16840_ (.A(_09261_),
    .B(_09224_),
    .Y(_09272_));
 sky130_fd_sc_hd__a22o_1 _16841_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[5] ),
    .A2(_08922_),
    .B1(_09271_),
    .B2(_09272_),
    .X(_00909_));
 sky130_fd_sc_hd__or3_1 _16842_ (.A(_09220_),
    .B(_09205_),
    .C(_09219_),
    .X(_09273_));
 sky130_fd_sc_hd__nor2_1 _16843_ (.A(_09261_),
    .B(_09221_),
    .Y(_09274_));
 sky130_fd_sc_hd__a22o_1 _16844_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[4] ),
    .A2(_08922_),
    .B1(_09273_),
    .B2(_09274_),
    .X(_00908_));
 sky130_fd_sc_hd__nor2_1 _16845_ (.A(_09209_),
    .B(_09217_),
    .Y(_09275_));
 sky130_fd_sc_hd__nand2_1 _16846_ (.A(_09218_),
    .B(_09275_),
    .Y(_09276_));
 sky130_fd_sc_hd__nor2_1 _16847_ (.A(_09261_),
    .B(_09219_),
    .Y(_09277_));
 sky130_fd_sc_hd__a22o_1 _16848_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[3] ),
    .A2(_08922_),
    .B1(_09276_),
    .B2(_09277_),
    .X(_00907_));
 sky130_fd_sc_hd__and3_1 _16849_ (.A(_09212_),
    .B(_09215_),
    .C(_09216_),
    .X(_09278_));
 sky130_fd_sc_hd__o32ai_1 _16850_ (.A1(_09261_),
    .A2(_09217_),
    .A3(_09278_),
    .B1(_09086_),
    .B2(_09206_),
    .Y(_00906_));
 sky130_fd_sc_hd__nand2_1 _16851_ (.A(_09213_),
    .B(_09214_),
    .Y(_09279_));
 sky130_fd_sc_hd__a32o_1 _16852_ (.A1(_08919_),
    .A2(_09215_),
    .A3(_09279_),
    .B1(_09054_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.y[1] ),
    .X(_00905_));
 sky130_fd_sc_hd__nor2_1 _16853_ (.A(_08895_),
    .B(_09125_),
    .Y(_09280_));
 sky130_fd_sc_hd__a21oi_1 _16854_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[0] ),
    .A2(_09280_),
    .B1(_09056_),
    .Y(_09281_));
 sky130_fd_sc_hd__o21a_1 _16855_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[0] ),
    .A2(_09280_),
    .B1(_09281_),
    .X(_00904_));
 sky130_fd_sc_hd__clkinv_2 _16856_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[15] ),
    .Y(_09282_));
 sky130_fd_sc_hd__mux2_1 _16857_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.y[15] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[16] ),
    .S(_08901_),
    .X(_09283_));
 sky130_fd_sc_hd__mux2_1 _16858_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.y[16] ),
    .A1(_09283_),
    .S(_08982_),
    .X(_09284_));
 sky130_fd_sc_hd__or2b_1 _16859_ (.A(\wfg_stim_sine_top.wfg_stim_sine.y[16] ),
    .B_N(_08908_),
    .X(_09285_));
 sky130_fd_sc_hd__o21a_1 _16860_ (.A1(_08909_),
    .A2(_09284_),
    .B1(_09285_),
    .X(_09286_));
 sky130_fd_sc_hd__or2_1 _16861_ (.A(_08962_),
    .B(\wfg_stim_sine_top.wfg_stim_sine.y[16] ),
    .X(_09287_));
 sky130_fd_sc_hd__clkbuf_2 _16862_ (.A(_09287_),
    .X(_09288_));
 sky130_fd_sc_hd__o21a_1 _16863_ (.A1(_08913_),
    .A2(_09286_),
    .B1(_09288_),
    .X(_09289_));
 sky130_fd_sc_hd__mux2_1 _16864_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.y[11] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[12] ),
    .S(_08901_),
    .X(_09290_));
 sky130_fd_sc_hd__mux2_1 _16865_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.y[13] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[14] ),
    .S(\wfg_stim_sine_top.wfg_stim_sine.iteration[0] ),
    .X(_09291_));
 sky130_fd_sc_hd__mux2_1 _16866_ (.A0(_09290_),
    .A1(_09291_),
    .S(_08910_),
    .X(_09292_));
 sky130_fd_sc_hd__mux2_1 _16867_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.y[9] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[10] ),
    .S(_08901_),
    .X(_09293_));
 sky130_fd_sc_hd__mux2_1 _16868_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.y[7] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[8] ),
    .S(_08901_),
    .X(_09294_));
 sky130_fd_sc_hd__mux2_1 _16869_ (.A0(_09293_),
    .A1(_09294_),
    .S(_08982_),
    .X(_09295_));
 sky130_fd_sc_hd__or2_1 _16870_ (.A(_08937_),
    .B(_09295_),
    .X(_09296_));
 sky130_fd_sc_hd__o221a_1 _16871_ (.A1(_08962_),
    .A2(_09286_),
    .B1(_09292_),
    .B2(_08967_),
    .C1(_09296_),
    .X(_09297_));
 sky130_fd_sc_hd__mux2_1 _16872_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.y[8] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[9] ),
    .S(\wfg_stim_sine_top.wfg_stim_sine.iteration[0] ),
    .X(_09298_));
 sky130_fd_sc_hd__mux2_1 _16873_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.y[10] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[11] ),
    .S(\wfg_stim_sine_top.wfg_stim_sine.iteration[0] ),
    .X(_09299_));
 sky130_fd_sc_hd__mux2_1 _16874_ (.A0(_09298_),
    .A1(_09299_),
    .S(_08899_),
    .X(_09300_));
 sky130_fd_sc_hd__mux2_1 _16875_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.y[12] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[13] ),
    .S(\wfg_stim_sine_top.wfg_stim_sine.iteration[0] ),
    .X(_09301_));
 sky130_fd_sc_hd__mux2_1 _16876_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.y[14] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[15] ),
    .S(\wfg_stim_sine_top.wfg_stim_sine.iteration[0] ),
    .X(_09302_));
 sky130_fd_sc_hd__mux2_1 _16877_ (.A0(_09301_),
    .A1(_09302_),
    .S(_08899_),
    .X(_09303_));
 sky130_fd_sc_hd__mux2_2 _16878_ (.A0(_09300_),
    .A1(_09303_),
    .S(\wfg_stim_sine_top.wfg_stim_sine.iteration[2] ),
    .X(_09304_));
 sky130_fd_sc_hd__mux2_1 _16879_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.y[4] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[5] ),
    .S(_08902_),
    .X(_09305_));
 sky130_fd_sc_hd__mux2_1 _16880_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.y[6] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[7] ),
    .S(_08902_),
    .X(_09306_));
 sky130_fd_sc_hd__mux2_1 _16881_ (.A0(_09305_),
    .A1(_09306_),
    .S(_08900_),
    .X(_09307_));
 sky130_fd_sc_hd__mux2_1 _16882_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.y[2] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[3] ),
    .S(_08902_),
    .X(_09308_));
 sky130_fd_sc_hd__o221a_1 _16883_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[0] ),
    .A2(_08921_),
    .B1(_08940_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.y[1] ),
    .C1(_08948_),
    .X(_09309_));
 sky130_fd_sc_hd__o21a_1 _16884_ (.A1(_08981_),
    .A2(_09308_),
    .B1(_09309_),
    .X(_09310_));
 sky130_fd_sc_hd__a221oi_4 _16885_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.iteration[3] ),
    .A2(_09304_),
    .B1(_09307_),
    .B2(_08976_),
    .C1(_09310_),
    .Y(_09311_));
 sky130_fd_sc_hd__mux2_1 _16886_ (.A0(_09293_),
    .A1(_09290_),
    .S(_08899_),
    .X(_09312_));
 sky130_fd_sc_hd__mux2_1 _16887_ (.A0(_09283_),
    .A1(_09291_),
    .S(_08981_),
    .X(_09313_));
 sky130_fd_sc_hd__mux2_1 _16888_ (.A0(_09312_),
    .A1(_09313_),
    .S(\wfg_stim_sine_top.wfg_stim_sine.iteration[2] ),
    .X(_09314_));
 sky130_fd_sc_hd__mux2_1 _16889_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.y[3] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[4] ),
    .S(_08901_),
    .X(_09315_));
 sky130_fd_sc_hd__or2_1 _16890_ (.A(_08981_),
    .B(_09315_),
    .X(_09316_));
 sky130_fd_sc_hd__o22a_1 _16891_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[1] ),
    .A2(_08921_),
    .B1(_08940_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.y[2] ),
    .X(_09317_));
 sky130_fd_sc_hd__mux2_1 _16892_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.y[5] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[6] ),
    .S(_08901_),
    .X(_09318_));
 sky130_fd_sc_hd__mux2_1 _16893_ (.A0(_09318_),
    .A1(_09294_),
    .S(_08899_),
    .X(_09319_));
 sky130_fd_sc_hd__a32o_1 _16894_ (.A1(_08948_),
    .A2(_09316_),
    .A3(_09317_),
    .B1(_09319_),
    .B2(_08976_),
    .X(_09320_));
 sky130_fd_sc_hd__a21oi_1 _16895_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.iteration[3] ),
    .A2(_09314_),
    .B1(_09320_),
    .Y(_09321_));
 sky130_fd_sc_hd__and2_1 _16896_ (.A(_09311_),
    .B(_09321_),
    .X(_09322_));
 sky130_fd_sc_hd__mux2_1 _16897_ (.A0(_09299_),
    .A1(_09301_),
    .S(_08900_),
    .X(_09323_));
 sky130_fd_sc_hd__mux2_1 _16898_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.y[16] ),
    .A1(_09302_),
    .S(_08981_),
    .X(_09324_));
 sky130_fd_sc_hd__or2b_1 _16899_ (.A(_09324_),
    .B_N(_08904_),
    .X(_09325_));
 sky130_fd_sc_hd__o21ai_1 _16900_ (.A1(_08904_),
    .A2(_09323_),
    .B1(_09325_),
    .Y(_09326_));
 sky130_fd_sc_hd__mux2_1 _16901_ (.A0(_09298_),
    .A1(_09306_),
    .S(_08981_),
    .X(_09327_));
 sky130_fd_sc_hd__and3_1 _16902_ (.A(_08900_),
    .B(_08948_),
    .C(_09305_),
    .X(_09328_));
 sky130_fd_sc_hd__a221o_1 _16903_ (.A1(_08944_),
    .A2(_09308_),
    .B1(_09327_),
    .B2(_08976_),
    .C1(_09328_),
    .X(_09329_));
 sky130_fd_sc_hd__o21ba_1 _16904_ (.A1(_08959_),
    .A2(_09326_),
    .B1_N(_09329_),
    .X(_09330_));
 sky130_fd_sc_hd__mux2_1 _16905_ (.A0(_09292_),
    .A1(_09284_),
    .S(_08908_),
    .X(_09331_));
 sky130_fd_sc_hd__and3_1 _16906_ (.A(_08910_),
    .B(_08948_),
    .C(_09318_),
    .X(_09332_));
 sky130_fd_sc_hd__a221o_1 _16907_ (.A1(_08944_),
    .A2(_09315_),
    .B1(_09295_),
    .B2(_08976_),
    .C1(_09332_),
    .X(_09333_));
 sky130_fd_sc_hd__a21oi_1 _16908_ (.A1(_08912_),
    .A2(_09331_),
    .B1(_09333_),
    .Y(_09334_));
 sky130_fd_sc_hd__nand3_1 _16909_ (.A(_09322_),
    .B(_09330_),
    .C(_09334_),
    .Y(_09335_));
 sky130_fd_sc_hd__o21a_1 _16910_ (.A1(_08908_),
    .A2(_09303_),
    .B1(_09285_),
    .X(_09336_));
 sky130_fd_sc_hd__or2_1 _16911_ (.A(_08937_),
    .B(_09307_),
    .X(_09337_));
 sky130_fd_sc_hd__o221a_1 _16912_ (.A1(_08967_),
    .A2(_09300_),
    .B1(_09336_),
    .B2(_08959_),
    .C1(_09337_),
    .X(_09338_));
 sky130_fd_sc_hd__o21ai_1 _16913_ (.A1(_08909_),
    .A2(_09313_),
    .B1(_09285_),
    .Y(_09339_));
 sky130_fd_sc_hd__nand2_1 _16914_ (.A(_08912_),
    .B(_09339_),
    .Y(_09340_));
 sky130_fd_sc_hd__o221a_1 _16915_ (.A1(_08967_),
    .A2(_09312_),
    .B1(_09319_),
    .B2(_08937_),
    .C1(_09340_),
    .X(_09341_));
 sky130_fd_sc_hd__nor3_1 _16916_ (.A(_09335_),
    .B(_09338_),
    .C(_09341_),
    .Y(_09342_));
 sky130_fd_sc_hd__o21a_1 _16917_ (.A1(_08909_),
    .A2(_09324_),
    .B1(_09285_),
    .X(_09343_));
 sky130_fd_sc_hd__o22a_1 _16918_ (.A1(_08967_),
    .A2(_09323_),
    .B1(_09327_),
    .B2(_08937_),
    .X(_09344_));
 sky130_fd_sc_hd__o21ai_1 _16919_ (.A1(_08962_),
    .A2(_09343_),
    .B1(_09344_),
    .Y(_09345_));
 sky130_fd_sc_hd__and3b_1 _16920_ (.A_N(_09297_),
    .B(_09342_),
    .C(_09345_),
    .X(_09346_));
 sky130_fd_sc_hd__o21ai_1 _16921_ (.A1(_08912_),
    .A2(_09304_),
    .B1(_09288_),
    .Y(_09347_));
 sky130_fd_sc_hd__and2_1 _16922_ (.A(_09346_),
    .B(_09347_),
    .X(_09348_));
 sky130_fd_sc_hd__o21ai_1 _16923_ (.A1(_08912_),
    .A2(_09314_),
    .B1(_09288_),
    .Y(_09349_));
 sky130_fd_sc_hd__a21bo_1 _16924_ (.A1(_08962_),
    .A2(_09326_),
    .B1_N(_09288_),
    .X(_09350_));
 sky130_fd_sc_hd__and3_1 _16925_ (.A(_09348_),
    .B(_09349_),
    .C(_09350_),
    .X(_09351_));
 sky130_fd_sc_hd__o21ai_1 _16926_ (.A1(_08913_),
    .A2(_09331_),
    .B1(_09288_),
    .Y(_09352_));
 sky130_fd_sc_hd__nand2_1 _16927_ (.A(_09351_),
    .B(_09352_),
    .Y(_09353_));
 sky130_fd_sc_hd__o21a_1 _16928_ (.A1(_08913_),
    .A2(_09336_),
    .B1(_09288_),
    .X(_09354_));
 sky130_fd_sc_hd__a21boi_1 _16929_ (.A1(_08962_),
    .A2(_09339_),
    .B1_N(_09288_),
    .Y(_09355_));
 sky130_fd_sc_hd__nor3_1 _16930_ (.A(_09353_),
    .B(_09354_),
    .C(_09355_),
    .Y(_09356_));
 sky130_fd_sc_hd__o21ai_1 _16931_ (.A1(_08913_),
    .A2(_09343_),
    .B1(_09288_),
    .Y(_09357_));
 sky130_fd_sc_hd__a21o_1 _16932_ (.A1(_09356_),
    .A2(_09357_),
    .B1(_08930_),
    .X(_09358_));
 sky130_fd_sc_hd__xor2_1 _16933_ (.A(_09289_),
    .B(_09358_),
    .X(_09359_));
 sky130_fd_sc_hd__or2_1 _16934_ (.A(_09282_),
    .B(_09359_),
    .X(_09360_));
 sky130_fd_sc_hd__or2_1 _16935_ (.A(_08930_),
    .B(_09356_),
    .X(_09361_));
 sky130_fd_sc_hd__xor2_1 _16936_ (.A(_09357_),
    .B(_09361_),
    .X(_09362_));
 sky130_fd_sc_hd__and2_1 _16937_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[14] ),
    .B(_09362_),
    .X(_09363_));
 sky130_fd_sc_hd__o21a_1 _16938_ (.A1(_09353_),
    .A2(_09354_),
    .B1(_09004_),
    .X(_09364_));
 sky130_fd_sc_hd__xor2_1 _16939_ (.A(_09355_),
    .B(_09364_),
    .X(_09365_));
 sky130_fd_sc_hd__nand2_1 _16940_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[13] ),
    .B(_09365_),
    .Y(_09366_));
 sky130_fd_sc_hd__nand2_1 _16941_ (.A(_09004_),
    .B(_09353_),
    .Y(_09367_));
 sky130_fd_sc_hd__xnor2_1 _16942_ (.A(_09354_),
    .B(_09367_),
    .Y(_09368_));
 sky130_fd_sc_hd__nand2_1 _16943_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[12] ),
    .B(_09368_),
    .Y(_09369_));
 sky130_fd_sc_hd__or2_1 _16944_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[12] ),
    .B(_09368_),
    .X(_09370_));
 sky130_fd_sc_hd__nand2_1 _16945_ (.A(_09369_),
    .B(_09370_),
    .Y(_09371_));
 sky130_fd_sc_hd__nor2_1 _16946_ (.A(_08929_),
    .B(_09351_),
    .Y(_09372_));
 sky130_fd_sc_hd__xnor2_1 _16947_ (.A(_09352_),
    .B(_09372_),
    .Y(_09373_));
 sky130_fd_sc_hd__a31o_1 _16948_ (.A1(_09346_),
    .A2(_09347_),
    .A3(_09349_),
    .B1(_08929_),
    .X(_09374_));
 sky130_fd_sc_hd__xor2_1 _16949_ (.A(_09350_),
    .B(_09374_),
    .X(_09375_));
 sky130_fd_sc_hd__and2_1 _16950_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[10] ),
    .B(_09375_),
    .X(_09376_));
 sky130_fd_sc_hd__nor2_1 _16951_ (.A(_08928_),
    .B(_09348_),
    .Y(_09377_));
 sky130_fd_sc_hd__xnor2_1 _16952_ (.A(_09349_),
    .B(_09377_),
    .Y(_09378_));
 sky130_fd_sc_hd__nand2_1 _16953_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[9] ),
    .B(_09378_),
    .Y(_09379_));
 sky130_fd_sc_hd__nor2_1 _16954_ (.A(_08928_),
    .B(_09346_),
    .Y(_09380_));
 sky130_fd_sc_hd__xnor2_1 _16955_ (.A(_09347_),
    .B(_09380_),
    .Y(_09381_));
 sky130_fd_sc_hd__nand2_1 _16956_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[8] ),
    .B(_09381_),
    .Y(_09382_));
 sky130_fd_sc_hd__a21o_1 _16957_ (.A1(_09342_),
    .A2(_09345_),
    .B1(_08928_),
    .X(_09383_));
 sky130_fd_sc_hd__xnor2_1 _16958_ (.A(_09297_),
    .B(_09383_),
    .Y(_09384_));
 sky130_fd_sc_hd__nand2_1 _16959_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[7] ),
    .B(_09384_),
    .Y(_09385_));
 sky130_fd_sc_hd__nor2_1 _16960_ (.A(_08927_),
    .B(_09342_),
    .Y(_09386_));
 sky130_fd_sc_hd__xnor2_1 _16961_ (.A(_09345_),
    .B(_09386_),
    .Y(_09387_));
 sky130_fd_sc_hd__nand2_1 _16962_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[6] ),
    .B(_09387_),
    .Y(_09388_));
 sky130_fd_sc_hd__o21a_1 _16963_ (.A1(_09335_),
    .A2(_09338_),
    .B1(_09004_),
    .X(_09389_));
 sky130_fd_sc_hd__xor2_1 _16964_ (.A(_09341_),
    .B(_09389_),
    .X(_09390_));
 sky130_fd_sc_hd__nand2_1 _16965_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[5] ),
    .B(_09390_),
    .Y(_09391_));
 sky130_fd_sc_hd__nand2_1 _16966_ (.A(_09004_),
    .B(_09335_),
    .Y(_09392_));
 sky130_fd_sc_hd__xnor2_1 _16967_ (.A(_09338_),
    .B(_09392_),
    .Y(_09393_));
 sky130_fd_sc_hd__nand2_1 _16968_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[4] ),
    .B(_09393_),
    .Y(_09394_));
 sky130_fd_sc_hd__a21oi_1 _16969_ (.A1(_09322_),
    .A2(_09330_),
    .B1(\wfg_stim_sine_top.wfg_stim_sine.z[16] ),
    .Y(_09395_));
 sky130_fd_sc_hd__xnor2_1 _16970_ (.A(_09334_),
    .B(_09395_),
    .Y(_09396_));
 sky130_fd_sc_hd__nand2_1 _16971_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[3] ),
    .B(_09396_),
    .Y(_09397_));
 sky130_fd_sc_hd__or2_1 _16972_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[16] ),
    .B(_09322_),
    .X(_09398_));
 sky130_fd_sc_hd__xor2_1 _16973_ (.A(_09330_),
    .B(_09398_),
    .X(_09399_));
 sky130_fd_sc_hd__nand2_1 _16974_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[2] ),
    .B(_09399_),
    .Y(_09400_));
 sky130_fd_sc_hd__nor2_1 _16975_ (.A(\wfg_stim_sine_top.wfg_stim_sine.z[16] ),
    .B(_09311_),
    .Y(_09401_));
 sky130_fd_sc_hd__xnor2_1 _16976_ (.A(_09321_),
    .B(_09401_),
    .Y(_09402_));
 sky130_fd_sc_hd__nand2_1 _16977_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[1] ),
    .B(_09402_),
    .Y(_09403_));
 sky130_fd_sc_hd__xor2_1 _16978_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[1] ),
    .B(_09402_),
    .X(_09404_));
 sky130_fd_sc_hd__and2b_1 _16979_ (.A_N(_09311_),
    .B(\wfg_stim_sine_top.wfg_stim_sine.x[0] ),
    .X(_09405_));
 sky130_fd_sc_hd__nand2_1 _16980_ (.A(_09404_),
    .B(_09405_),
    .Y(_09406_));
 sky130_fd_sc_hd__xor2_1 _16981_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[2] ),
    .B(_09399_),
    .X(_09407_));
 sky130_fd_sc_hd__a21bo_1 _16982_ (.A1(_09403_),
    .A2(_09406_),
    .B1_N(_09407_),
    .X(_09408_));
 sky130_fd_sc_hd__or2_1 _16983_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[3] ),
    .B(_09396_),
    .X(_09409_));
 sky130_fd_sc_hd__and2_1 _16984_ (.A(_09397_),
    .B(_09409_),
    .X(_09410_));
 sky130_fd_sc_hd__a21bo_1 _16985_ (.A1(_09400_),
    .A2(_09408_),
    .B1_N(_09410_),
    .X(_09411_));
 sky130_fd_sc_hd__or2_1 _16986_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[4] ),
    .B(_09393_),
    .X(_09412_));
 sky130_fd_sc_hd__nand2_1 _16987_ (.A(_09394_),
    .B(_09412_),
    .Y(_09413_));
 sky130_fd_sc_hd__a21o_1 _16988_ (.A1(_09397_),
    .A2(_09411_),
    .B1(_09413_),
    .X(_09414_));
 sky130_fd_sc_hd__or2_1 _16989_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[5] ),
    .B(_09390_),
    .X(_09415_));
 sky130_fd_sc_hd__nand2_1 _16990_ (.A(_09391_),
    .B(_09415_),
    .Y(_09416_));
 sky130_fd_sc_hd__a21o_1 _16991_ (.A1(_09394_),
    .A2(_09414_),
    .B1(_09416_),
    .X(_09417_));
 sky130_fd_sc_hd__or2_1 _16992_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[6] ),
    .B(_09387_),
    .X(_09418_));
 sky130_fd_sc_hd__nand2_1 _16993_ (.A(_09388_),
    .B(_09418_),
    .Y(_09419_));
 sky130_fd_sc_hd__a21o_1 _16994_ (.A1(_09391_),
    .A2(_09417_),
    .B1(_09419_),
    .X(_09420_));
 sky130_fd_sc_hd__or2_1 _16995_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[7] ),
    .B(_09384_),
    .X(_09421_));
 sky130_fd_sc_hd__nand2_1 _16996_ (.A(_09385_),
    .B(_09421_),
    .Y(_09422_));
 sky130_fd_sc_hd__a21o_1 _16997_ (.A1(_09388_),
    .A2(_09420_),
    .B1(_09422_),
    .X(_09423_));
 sky130_fd_sc_hd__or2_1 _16998_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[8] ),
    .B(_09381_),
    .X(_09424_));
 sky130_fd_sc_hd__nand2_1 _16999_ (.A(_09382_),
    .B(_09424_),
    .Y(_09425_));
 sky130_fd_sc_hd__a21o_1 _17000_ (.A1(_09385_),
    .A2(_09423_),
    .B1(_09425_),
    .X(_09426_));
 sky130_fd_sc_hd__or2_1 _17001_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[9] ),
    .B(_09378_),
    .X(_09427_));
 sky130_fd_sc_hd__nand2_1 _17002_ (.A(_09379_),
    .B(_09427_),
    .Y(_09428_));
 sky130_fd_sc_hd__a21o_1 _17003_ (.A1(_09382_),
    .A2(_09426_),
    .B1(_09428_),
    .X(_09429_));
 sky130_fd_sc_hd__nor2_1 _17004_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[10] ),
    .B(_09375_),
    .Y(_09430_));
 sky130_fd_sc_hd__or2_1 _17005_ (.A(_09376_),
    .B(_09430_),
    .X(_09431_));
 sky130_fd_sc_hd__a21oi_1 _17006_ (.A1(_09379_),
    .A2(_09429_),
    .B1(_09431_),
    .Y(_09432_));
 sky130_fd_sc_hd__xnor2_1 _17007_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[11] ),
    .B(_09373_),
    .Y(_09433_));
 sky130_fd_sc_hd__o21ba_1 _17008_ (.A1(_09376_),
    .A2(_09432_),
    .B1_N(_09433_),
    .X(_09434_));
 sky130_fd_sc_hd__a21o_1 _17009_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.x[11] ),
    .A2(_09373_),
    .B1(_09434_),
    .X(_09435_));
 sky130_fd_sc_hd__or2b_1 _17010_ (.A(_09371_),
    .B_N(_09435_),
    .X(_09436_));
 sky130_fd_sc_hd__or2_1 _17011_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[13] ),
    .B(_09365_),
    .X(_09437_));
 sky130_fd_sc_hd__nand2_1 _17012_ (.A(_09366_),
    .B(_09437_),
    .Y(_09438_));
 sky130_fd_sc_hd__a21o_1 _17013_ (.A1(_09369_),
    .A2(_09436_),
    .B1(_09438_),
    .X(_09439_));
 sky130_fd_sc_hd__nor2_1 _17014_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[14] ),
    .B(_09362_),
    .Y(_09440_));
 sky130_fd_sc_hd__or2_1 _17015_ (.A(_09363_),
    .B(_09440_),
    .X(_09441_));
 sky130_fd_sc_hd__a21oi_1 _17016_ (.A1(_09366_),
    .A2(_09439_),
    .B1(_09441_),
    .Y(_09442_));
 sky130_fd_sc_hd__nand2_1 _17017_ (.A(_09282_),
    .B(_09359_),
    .Y(_09443_));
 sky130_fd_sc_hd__and2_1 _17018_ (.A(_09360_),
    .B(_09443_),
    .X(_09444_));
 sky130_fd_sc_hd__o21ai_1 _17019_ (.A1(_09363_),
    .A2(_09442_),
    .B1(_09444_),
    .Y(_09445_));
 sky130_fd_sc_hd__a21boi_1 _17020_ (.A1(_09004_),
    .A2(_09289_),
    .B1_N(_09358_),
    .Y(_09446_));
 sky130_fd_sc_hd__xor2_1 _17021_ (.A(_09251_),
    .B(_09446_),
    .X(_09447_));
 sky130_fd_sc_hd__a21oi_1 _17022_ (.A1(_09360_),
    .A2(_09445_),
    .B1(_09447_),
    .Y(_09448_));
 sky130_fd_sc_hd__a31o_1 _17023_ (.A1(_09360_),
    .A2(_09445_),
    .A3(_09447_),
    .B1(_08915_),
    .X(_09449_));
 sky130_fd_sc_hd__a2bb2o_1 _17024_ (.A1_N(_09448_),
    .A2_N(_09449_),
    .B1(\wfg_stim_sine_top.wfg_stim_sine.x[16] ),
    .B2(_08896_),
    .X(_00903_));
 sky130_fd_sc_hd__or3_1 _17025_ (.A(_09444_),
    .B(_09363_),
    .C(_09442_),
    .X(_09450_));
 sky130_fd_sc_hd__a21oi_1 _17026_ (.A1(_09445_),
    .A2(_09450_),
    .B1(_09261_),
    .Y(_09451_));
 sky130_fd_sc_hd__a21oi_1 _17027_ (.A1(_09282_),
    .A2(_08922_),
    .B1(_09451_),
    .Y(_00902_));
 sky130_fd_sc_hd__and3_1 _17028_ (.A(_09441_),
    .B(_09366_),
    .C(_09439_),
    .X(_09452_));
 sky130_fd_sc_hd__nor2_1 _17029_ (.A(_09442_),
    .B(_09452_),
    .Y(_09453_));
 sky130_fd_sc_hd__a22o_1 _17030_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.x[14] ),
    .A2(_08922_),
    .B1(_09050_),
    .B2(_09453_),
    .X(_00901_));
 sky130_fd_sc_hd__nand3_1 _17031_ (.A(_09438_),
    .B(_09369_),
    .C(_09436_),
    .Y(_09454_));
 sky130_fd_sc_hd__a32o_1 _17032_ (.A1(_08919_),
    .A2(_09439_),
    .A3(_09454_),
    .B1(_09054_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.x[13] ),
    .X(_00900_));
 sky130_fd_sc_hd__xnor2_1 _17033_ (.A(_09371_),
    .B(_09435_),
    .Y(_09455_));
 sky130_fd_sc_hd__o22a_1 _17034_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.x[12] ),
    .A2(_09086_),
    .B1(_08916_),
    .B2(_09455_),
    .X(_00899_));
 sky130_fd_sc_hd__or2_1 _17035_ (.A(_09376_),
    .B(_09432_),
    .X(_09456_));
 sky130_fd_sc_hd__xnor2_1 _17036_ (.A(_09433_),
    .B(_09456_),
    .Y(_09457_));
 sky130_fd_sc_hd__o22a_1 _17037_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.x[11] ),
    .A2(_09086_),
    .B1(_08916_),
    .B2(_09457_),
    .X(_00898_));
 sky130_fd_sc_hd__and3_1 _17038_ (.A(_09431_),
    .B(_09379_),
    .C(_09429_),
    .X(_09458_));
 sky130_fd_sc_hd__nor2_1 _17039_ (.A(_09432_),
    .B(_09458_),
    .Y(_09459_));
 sky130_fd_sc_hd__a22o_1 _17040_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.x[10] ),
    .A2(_08922_),
    .B1(_09050_),
    .B2(_09459_),
    .X(_00897_));
 sky130_fd_sc_hd__nand3_1 _17041_ (.A(_09428_),
    .B(_09382_),
    .C(_09426_),
    .Y(_09460_));
 sky130_fd_sc_hd__and2_1 _17042_ (.A(_09429_),
    .B(_09460_),
    .X(_09461_));
 sky130_fd_sc_hd__o22a_1 _17043_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.x[9] ),
    .A2(_09086_),
    .B1(_08916_),
    .B2(_09461_),
    .X(_00896_));
 sky130_fd_sc_hd__nand3_1 _17044_ (.A(_09425_),
    .B(_09385_),
    .C(_09423_),
    .Y(_09462_));
 sky130_fd_sc_hd__and2_1 _17045_ (.A(_09426_),
    .B(_09462_),
    .X(_09463_));
 sky130_fd_sc_hd__o22a_1 _17046_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.x[8] ),
    .A2(_09086_),
    .B1(_08916_),
    .B2(_09463_),
    .X(_00895_));
 sky130_fd_sc_hd__nand3_1 _17047_ (.A(_09422_),
    .B(_09388_),
    .C(_09420_),
    .Y(_09464_));
 sky130_fd_sc_hd__a32o_1 _17048_ (.A1(_08919_),
    .A2(_09423_),
    .A3(_09464_),
    .B1(_09054_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.x[7] ),
    .X(_00894_));
 sky130_fd_sc_hd__nand3_1 _17049_ (.A(_09419_),
    .B(_09391_),
    .C(_09417_),
    .Y(_09465_));
 sky130_fd_sc_hd__and2_1 _17050_ (.A(_09420_),
    .B(_09465_),
    .X(_09466_));
 sky130_fd_sc_hd__o22a_1 _17051_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.x[6] ),
    .A2(_09086_),
    .B1(_08916_),
    .B2(_09466_),
    .X(_00893_));
 sky130_fd_sc_hd__nand3_1 _17052_ (.A(_09416_),
    .B(_09394_),
    .C(_09414_),
    .Y(_09467_));
 sky130_fd_sc_hd__and2_1 _17053_ (.A(_09417_),
    .B(_09467_),
    .X(_09468_));
 sky130_fd_sc_hd__o22a_1 _17054_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.x[5] ),
    .A2(_09086_),
    .B1(_08916_),
    .B2(_09468_),
    .X(_00892_));
 sky130_fd_sc_hd__nand3_1 _17055_ (.A(_09413_),
    .B(_09397_),
    .C(_09411_),
    .Y(_09469_));
 sky130_fd_sc_hd__and2_1 _17056_ (.A(_09414_),
    .B(_09469_),
    .X(_09470_));
 sky130_fd_sc_hd__o22a_1 _17057_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.x[4] ),
    .A2(_09086_),
    .B1(_08916_),
    .B2(_09470_),
    .X(_00891_));
 sky130_fd_sc_hd__nand3b_1 _17058_ (.A_N(_09410_),
    .B(_09400_),
    .C(_09408_),
    .Y(_09471_));
 sky130_fd_sc_hd__a32o_1 _17059_ (.A1(_08919_),
    .A2(_09411_),
    .A3(_09471_),
    .B1(_09054_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.x[3] ),
    .X(_00890_));
 sky130_fd_sc_hd__nand2_1 _17060_ (.A(_09403_),
    .B(_09406_),
    .Y(_09472_));
 sky130_fd_sc_hd__xor2_1 _17061_ (.A(_09472_),
    .B(_09407_),
    .X(_09473_));
 sky130_fd_sc_hd__o22a_1 _17062_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.x[2] ),
    .A2(_09086_),
    .B1(_08916_),
    .B2(_09473_),
    .X(_00889_));
 sky130_fd_sc_hd__or2_1 _17063_ (.A(_09404_),
    .B(_09405_),
    .X(_09474_));
 sky130_fd_sc_hd__a32o_1 _17064_ (.A1(_08919_),
    .A2(_09406_),
    .A3(_09474_),
    .B1(_09054_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.x[1] ),
    .X(_00888_));
 sky130_fd_sc_hd__or2b_1 _17065_ (.A(\wfg_stim_sine_top.wfg_stim_sine.x[0] ),
    .B_N(_09311_),
    .X(_09475_));
 sky130_fd_sc_hd__nor2_1 _17066_ (.A(_09261_),
    .B(_09405_),
    .Y(_09476_));
 sky130_fd_sc_hd__a22o_1 _17067_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.x[0] ),
    .A2(_08922_),
    .B1(_09475_),
    .B2(_09476_),
    .X(_00887_));
 sky130_fd_sc_hd__or2_1 _17068_ (.A(\wfg_stim_sine_top.offset_val_q[17] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[31] ),
    .X(_09477_));
 sky130_fd_sc_hd__and2_1 _17069_ (.A(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[17] ),
    .B(_09477_),
    .X(_09478_));
 sky130_fd_sc_hd__nand2_1 _17070_ (.A(\wfg_stim_sine_top.offset_val_q[17] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[31] ),
    .Y(_09479_));
 sky130_fd_sc_hd__nand2_1 _17071_ (.A(_00023_),
    .B(_09479_),
    .Y(_09480_));
 sky130_fd_sc_hd__o22a_1 _17072_ (.A1(\wfg_interconnect_top.stimulus_0[17] ),
    .A2(_00023_),
    .B1(_09478_),
    .B2(_09480_),
    .X(_00886_));
 sky130_fd_sc_hd__buf_2 _17073_ (.A(_06356_),
    .X(_09481_));
 sky130_fd_sc_hd__inv_2 _17074_ (.A(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[17] ),
    .Y(_09482_));
 sky130_fd_sc_hd__nor2_2 _17075_ (.A(_09482_),
    .B(_09477_),
    .Y(_09483_));
 sky130_fd_sc_hd__clkbuf_2 _17076_ (.A(_09483_),
    .X(_09484_));
 sky130_fd_sc_hd__or2_1 _17077_ (.A(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[16] ),
    .B(_09484_),
    .X(_09485_));
 sky130_fd_sc_hd__o21a_2 _17078_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[17] ),
    .A2(_09479_),
    .B1(_00023_),
    .X(_09486_));
 sky130_fd_sc_hd__a22o_1 _17079_ (.A1(\wfg_interconnect_top.stimulus_0[16] ),
    .A2(_09481_),
    .B1(_09485_),
    .B2(_09486_),
    .X(_00885_));
 sky130_fd_sc_hd__buf_2 _17080_ (.A(_09486_),
    .X(_09487_));
 sky130_fd_sc_hd__or2_1 _17081_ (.A(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[15] ),
    .B(_09484_),
    .X(_09488_));
 sky130_fd_sc_hd__a22o_1 _17082_ (.A1(\wfg_interconnect_top.stimulus_0[15] ),
    .A2(_09481_),
    .B1(_09487_),
    .B2(_09488_),
    .X(_00884_));
 sky130_fd_sc_hd__or2_1 _17083_ (.A(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[14] ),
    .B(_09484_),
    .X(_09489_));
 sky130_fd_sc_hd__a22o_1 _17084_ (.A1(\wfg_interconnect_top.stimulus_0[14] ),
    .A2(_09481_),
    .B1(_09487_),
    .B2(_09489_),
    .X(_00883_));
 sky130_fd_sc_hd__or2_1 _17085_ (.A(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[13] ),
    .B(_09484_),
    .X(_09490_));
 sky130_fd_sc_hd__a22o_1 _17086_ (.A1(\wfg_interconnect_top.stimulus_0[13] ),
    .A2(_09481_),
    .B1(_09487_),
    .B2(_09490_),
    .X(_00882_));
 sky130_fd_sc_hd__or2_1 _17087_ (.A(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[12] ),
    .B(_09484_),
    .X(_09491_));
 sky130_fd_sc_hd__a22o_1 _17088_ (.A1(\wfg_interconnect_top.stimulus_0[12] ),
    .A2(_09481_),
    .B1(_09487_),
    .B2(_09491_),
    .X(_00881_));
 sky130_fd_sc_hd__or2_1 _17089_ (.A(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[11] ),
    .B(_09484_),
    .X(_09492_));
 sky130_fd_sc_hd__a22o_1 _17090_ (.A1(\wfg_interconnect_top.stimulus_0[11] ),
    .A2(_09481_),
    .B1(_09487_),
    .B2(_09492_),
    .X(_00880_));
 sky130_fd_sc_hd__or2_1 _17091_ (.A(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[10] ),
    .B(_09484_),
    .X(_09493_));
 sky130_fd_sc_hd__a22o_1 _17092_ (.A1(\wfg_interconnect_top.stimulus_0[10] ),
    .A2(_09481_),
    .B1(_09487_),
    .B2(_09493_),
    .X(_00879_));
 sky130_fd_sc_hd__or2_1 _17093_ (.A(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[9] ),
    .B(_09484_),
    .X(_09494_));
 sky130_fd_sc_hd__a22o_1 _17094_ (.A1(\wfg_interconnect_top.stimulus_0[9] ),
    .A2(_09481_),
    .B1(_09487_),
    .B2(_09494_),
    .X(_00878_));
 sky130_fd_sc_hd__or2_1 _17095_ (.A(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[8] ),
    .B(_09484_),
    .X(_09495_));
 sky130_fd_sc_hd__a22o_1 _17096_ (.A1(\wfg_interconnect_top.stimulus_0[8] ),
    .A2(_09481_),
    .B1(_09487_),
    .B2(_09495_),
    .X(_00877_));
 sky130_fd_sc_hd__or2_1 _17097_ (.A(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[7] ),
    .B(_09484_),
    .X(_09496_));
 sky130_fd_sc_hd__a22o_1 _17098_ (.A1(\wfg_interconnect_top.stimulus_0[7] ),
    .A2(_09481_),
    .B1(_09487_),
    .B2(_09496_),
    .X(_00876_));
 sky130_fd_sc_hd__or2_1 _17099_ (.A(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[6] ),
    .B(_09483_),
    .X(_09497_));
 sky130_fd_sc_hd__a22o_1 _17100_ (.A1(\wfg_interconnect_top.stimulus_0[6] ),
    .A2(_06356_),
    .B1(_09487_),
    .B2(_09497_),
    .X(_00875_));
 sky130_fd_sc_hd__or2_1 _17101_ (.A(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[5] ),
    .B(_09483_),
    .X(_09498_));
 sky130_fd_sc_hd__a22o_1 _17102_ (.A1(\wfg_interconnect_top.stimulus_0[5] ),
    .A2(_06356_),
    .B1(_09486_),
    .B2(_09498_),
    .X(_00874_));
 sky130_fd_sc_hd__or2_1 _17103_ (.A(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[4] ),
    .B(_09483_),
    .X(_09499_));
 sky130_fd_sc_hd__a22o_1 _17104_ (.A1(\wfg_interconnect_top.stimulus_0[4] ),
    .A2(_06356_),
    .B1(_09486_),
    .B2(_09499_),
    .X(_00873_));
 sky130_fd_sc_hd__or2_1 _17105_ (.A(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[3] ),
    .B(_09483_),
    .X(_09500_));
 sky130_fd_sc_hd__a22o_1 _17106_ (.A1(\wfg_interconnect_top.stimulus_0[3] ),
    .A2(_06356_),
    .B1(_09486_),
    .B2(_09500_),
    .X(_00872_));
 sky130_fd_sc_hd__or2_1 _17107_ (.A(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[2] ),
    .B(_09483_),
    .X(_09501_));
 sky130_fd_sc_hd__a22o_1 _17108_ (.A1(\wfg_interconnect_top.stimulus_0[2] ),
    .A2(_06356_),
    .B1(_09486_),
    .B2(_09501_),
    .X(_00871_));
 sky130_fd_sc_hd__or2_1 _17109_ (.A(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[1] ),
    .B(_09483_),
    .X(_09502_));
 sky130_fd_sc_hd__a22o_1 _17110_ (.A1(\wfg_interconnect_top.stimulus_0[1] ),
    .A2(_06356_),
    .B1(_09486_),
    .B2(_09502_),
    .X(_00870_));
 sky130_fd_sc_hd__or2_1 _17111_ (.A(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[0] ),
    .B(_09483_),
    .X(_09503_));
 sky130_fd_sc_hd__a22o_1 _17112_ (.A1(\wfg_interconnect_top.stimulus_0[0] ),
    .A2(_06356_),
    .B1(_09486_),
    .B2(_09503_),
    .X(_00869_));
 sky130_fd_sc_hd__nand2_2 _17113_ (.A(\wfg_stim_sine_top.wfg_stim_sine.quadrant[1] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.quadrant[0] ),
    .Y(_09504_));
 sky130_fd_sc_hd__mux2_1 _17114_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[0] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[0] ),
    .S(_09504_),
    .X(_09505_));
 sky130_fd_sc_hd__mux2_1 _17115_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[1] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[1] ),
    .S(_09504_),
    .X(_09506_));
 sky130_fd_sc_hd__or2_1 _17116_ (.A(_09505_),
    .B(_09506_),
    .X(_09507_));
 sky130_fd_sc_hd__mux2_1 _17117_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[2] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[2] ),
    .S(_09504_),
    .X(_09508_));
 sky130_fd_sc_hd__or2_1 _17118_ (.A(_09507_),
    .B(_09508_),
    .X(_09509_));
 sky130_fd_sc_hd__mux2_1 _17119_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[3] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[3] ),
    .S(_09504_),
    .X(_09510_));
 sky130_fd_sc_hd__or2_1 _17120_ (.A(_09509_),
    .B(_09510_),
    .X(_09511_));
 sky130_fd_sc_hd__mux2_1 _17121_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[4] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[4] ),
    .S(_09504_),
    .X(_09512_));
 sky130_fd_sc_hd__or2_1 _17122_ (.A(_09511_),
    .B(_09512_),
    .X(_09513_));
 sky130_fd_sc_hd__mux2_1 _17123_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[5] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[5] ),
    .S(_09504_),
    .X(_09514_));
 sky130_fd_sc_hd__or2_1 _17124_ (.A(_09513_),
    .B(_09514_),
    .X(_09515_));
 sky130_fd_sc_hd__clkbuf_4 _17125_ (.A(_09504_),
    .X(_09516_));
 sky130_fd_sc_hd__mux2_1 _17126_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[6] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[6] ),
    .S(_09516_),
    .X(_09517_));
 sky130_fd_sc_hd__nor2_1 _17127_ (.A(_09515_),
    .B(_09517_),
    .Y(_09518_));
 sky130_fd_sc_hd__mux2_1 _17128_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[7] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[7] ),
    .S(_09516_),
    .X(_09519_));
 sky130_fd_sc_hd__inv_2 _17129_ (.A(_09519_),
    .Y(_09520_));
 sky130_fd_sc_hd__nand2_1 _17130_ (.A(_09518_),
    .B(_09520_),
    .Y(_09521_));
 sky130_fd_sc_hd__mux2_1 _17131_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[8] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[8] ),
    .S(_09516_),
    .X(_09522_));
 sky130_fd_sc_hd__nor2_1 _17132_ (.A(_09521_),
    .B(_09522_),
    .Y(_09523_));
 sky130_fd_sc_hd__mux2_1 _17133_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[9] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[9] ),
    .S(_09516_),
    .X(_09524_));
 sky130_fd_sc_hd__inv_2 _17134_ (.A(_09524_),
    .Y(_09525_));
 sky130_fd_sc_hd__nand2_1 _17135_ (.A(_09523_),
    .B(_09525_),
    .Y(_09526_));
 sky130_fd_sc_hd__mux2_1 _17136_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[10] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[10] ),
    .S(_09516_),
    .X(_09527_));
 sky130_fd_sc_hd__nor2_1 _17137_ (.A(_09526_),
    .B(_09527_),
    .Y(_09528_));
 sky130_fd_sc_hd__mux2_1 _17138_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[11] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[11] ),
    .S(_09516_),
    .X(_09529_));
 sky130_fd_sc_hd__inv_2 _17139_ (.A(_09529_),
    .Y(_09530_));
 sky130_fd_sc_hd__nand2_1 _17140_ (.A(_09528_),
    .B(_09530_),
    .Y(_09531_));
 sky130_fd_sc_hd__mux2_1 _17141_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[12] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[12] ),
    .S(_09516_),
    .X(_09532_));
 sky130_fd_sc_hd__nor2_1 _17142_ (.A(_09531_),
    .B(_09532_),
    .Y(_09533_));
 sky130_fd_sc_hd__mux2_1 _17143_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[13] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[13] ),
    .S(_09516_),
    .X(_09534_));
 sky130_fd_sc_hd__inv_2 _17144_ (.A(_09534_),
    .Y(_09535_));
 sky130_fd_sc_hd__nand2_1 _17145_ (.A(_09533_),
    .B(_09535_),
    .Y(_09536_));
 sky130_fd_sc_hd__mux2_1 _17146_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[14] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[14] ),
    .S(_09516_),
    .X(_09537_));
 sky130_fd_sc_hd__nor2_1 _17147_ (.A(_09536_),
    .B(_09537_),
    .Y(_09538_));
 sky130_fd_sc_hd__mux2_1 _17148_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.x[15] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.y[15] ),
    .S(_09516_),
    .X(_09539_));
 sky130_fd_sc_hd__inv_2 _17149_ (.A(_09539_),
    .Y(_09540_));
 sky130_fd_sc_hd__inv_2 _17150_ (.A(\wfg_stim_sine_top.wfg_stim_sine.quadrant[1] ),
    .Y(_09541_));
 sky130_fd_sc_hd__a21oi_4 _17151_ (.A1(_09538_),
    .A2(_09540_),
    .B1(_09541_),
    .Y(_09542_));
 sky130_fd_sc_hd__mux2_2 _17152_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.y[16] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.x[16] ),
    .S(\wfg_stim_sine_top.wfg_stim_sine.quadrant[0] ),
    .X(_09543_));
 sky130_fd_sc_hd__xor2_4 _17153_ (.A(_09542_),
    .B(_09543_),
    .X(_09544_));
 sky130_fd_sc_hd__nor3b_4 _17154_ (.A(\wfg_stim_sine_top.wfg_stim_sine.cur_state[2] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.cur_state[0] ),
    .C_N(\wfg_stim_sine_top.wfg_stim_sine.cur_state[1] ),
    .Y(_09545_));
 sky130_fd_sc_hd__mux2_1 _17155_ (.A0(_08085_),
    .A1(_09544_),
    .S(_09545_),
    .X(_09546_));
 sky130_fd_sc_hd__clkbuf_1 _17156_ (.A(_09546_),
    .X(_00868_));
 sky130_fd_sc_hd__or3b_1 _17157_ (.A(\wfg_stim_sine_top.wfg_stim_sine.cur_state[2] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.cur_state[0] ),
    .C_N(\wfg_stim_sine_top.wfg_stim_sine.cur_state[1] ),
    .X(_09547_));
 sky130_fd_sc_hd__buf_2 _17158_ (.A(_09547_),
    .X(_09548_));
 sky130_fd_sc_hd__buf_2 _17159_ (.A(_09548_),
    .X(_09549_));
 sky130_fd_sc_hd__o21a_1 _17160_ (.A1(_09538_),
    .A2(_09540_),
    .B1(_09542_),
    .X(_09550_));
 sky130_fd_sc_hd__a21oi_1 _17161_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.quadrant[0] ),
    .A2(_09282_),
    .B1(\wfg_stim_sine_top.wfg_stim_sine.quadrant[1] ),
    .Y(_09551_));
 sky130_fd_sc_hd__or2_2 _17162_ (.A(\wfg_stim_sine_top.wfg_stim_sine.quadrant[1] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.quadrant[0] ),
    .X(_09552_));
 sky130_fd_sc_hd__buf_2 _17163_ (.A(_09552_),
    .X(_09553_));
 sky130_fd_sc_hd__buf_2 _17164_ (.A(_09545_),
    .X(_09554_));
 sky130_fd_sc_hd__o221a_2 _17165_ (.A1(_09550_),
    .A2(_09551_),
    .B1(_09553_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.y[15] ),
    .C1(_09554_),
    .X(_09555_));
 sky130_fd_sc_hd__a21o_1 _17166_ (.A1(_06672_),
    .A2(_09549_),
    .B1(_09555_),
    .X(_00867_));
 sky130_fd_sc_hd__buf_2 _17167_ (.A(_09541_),
    .X(_09556_));
 sky130_fd_sc_hd__nor2_1 _17168_ (.A(_09541_),
    .B(_09538_),
    .Y(_09557_));
 sky130_fd_sc_hd__nand2_1 _17169_ (.A(_09536_),
    .B(_09537_),
    .Y(_09558_));
 sky130_fd_sc_hd__nor2_1 _17170_ (.A(\wfg_stim_sine_top.wfg_stim_sine.quadrant[1] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.quadrant[0] ),
    .Y(_09559_));
 sky130_fd_sc_hd__a221o_2 _17171_ (.A1(_09556_),
    .A2(\wfg_stim_sine_top.wfg_stim_sine.x[14] ),
    .B1(_09557_),
    .B2(_09558_),
    .C1(_09559_),
    .X(_09560_));
 sky130_fd_sc_hd__o21a_2 _17172_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[14] ),
    .A2(_09553_),
    .B1(_09554_),
    .X(_09561_));
 sky130_fd_sc_hd__a22o_1 _17173_ (.A1(_06510_),
    .A2(_09549_),
    .B1(_09560_),
    .B2(_09561_),
    .X(_00866_));
 sky130_fd_sc_hd__or2_1 _17174_ (.A(_09533_),
    .B(_09535_),
    .X(_09562_));
 sky130_fd_sc_hd__a21o_1 _17175_ (.A1(_09536_),
    .A2(_09562_),
    .B1(_09556_),
    .X(_09563_));
 sky130_fd_sc_hd__nand2_1 _17176_ (.A(_09541_),
    .B(\wfg_stim_sine_top.wfg_stim_sine.quadrant[0] ),
    .Y(_09564_));
 sky130_fd_sc_hd__buf_2 _17177_ (.A(_09564_),
    .X(_09565_));
 sky130_fd_sc_hd__o221a_2 _17178_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[13] ),
    .A2(_09553_),
    .B1(_09565_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.x[13] ),
    .C1(_09554_),
    .X(_09566_));
 sky130_fd_sc_hd__a22o_1 _17179_ (.A1(_06513_),
    .A2(_09549_),
    .B1(_09563_),
    .B2(_09566_),
    .X(_00865_));
 sky130_fd_sc_hd__and2_1 _17180_ (.A(_09531_),
    .B(_09532_),
    .X(_09567_));
 sky130_fd_sc_hd__o21ai_2 _17181_ (.A1(_09533_),
    .A2(_09567_),
    .B1(\wfg_stim_sine_top.wfg_stim_sine.quadrant[1] ),
    .Y(_09568_));
 sky130_fd_sc_hd__o221a_2 _17182_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[12] ),
    .A2(_09553_),
    .B1(_09565_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.x[12] ),
    .C1(_09554_),
    .X(_09569_));
 sky130_fd_sc_hd__a22o_1 _17183_ (.A1(_06423_),
    .A2(_09549_),
    .B1(_09568_),
    .B2(_09569_),
    .X(_00864_));
 sky130_fd_sc_hd__or2_1 _17184_ (.A(_09528_),
    .B(_09530_),
    .X(_09570_));
 sky130_fd_sc_hd__a21o_1 _17185_ (.A1(_09531_),
    .A2(_09570_),
    .B1(_09556_),
    .X(_09571_));
 sky130_fd_sc_hd__o221a_2 _17186_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[11] ),
    .A2(_09553_),
    .B1(_09565_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.x[11] ),
    .C1(_09554_),
    .X(_09572_));
 sky130_fd_sc_hd__a22o_1 _17187_ (.A1(_06432_),
    .A2(_09549_),
    .B1(_09571_),
    .B2(_09572_),
    .X(_00863_));
 sky130_fd_sc_hd__and2_1 _17188_ (.A(_09526_),
    .B(_09527_),
    .X(_09573_));
 sky130_fd_sc_hd__o21ai_2 _17189_ (.A1(_09528_),
    .A2(_09573_),
    .B1(\wfg_stim_sine_top.wfg_stim_sine.quadrant[1] ),
    .Y(_09574_));
 sky130_fd_sc_hd__o221a_2 _17190_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[10] ),
    .A2(_09553_),
    .B1(_09565_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.x[10] ),
    .C1(_09554_),
    .X(_09575_));
 sky130_fd_sc_hd__a22o_1 _17191_ (.A1(_06770_),
    .A2(_09549_),
    .B1(_09574_),
    .B2(_09575_),
    .X(_00862_));
 sky130_fd_sc_hd__or2_1 _17192_ (.A(_09523_),
    .B(_09525_),
    .X(_09576_));
 sky130_fd_sc_hd__a21o_1 _17193_ (.A1(_09526_),
    .A2(_09576_),
    .B1(_09556_),
    .X(_09577_));
 sky130_fd_sc_hd__o221a_2 _17194_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[9] ),
    .A2(_09553_),
    .B1(_09565_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.x[9] ),
    .C1(_09554_),
    .X(_09578_));
 sky130_fd_sc_hd__a22o_1 _17195_ (.A1(_06430_),
    .A2(_09549_),
    .B1(_09577_),
    .B2(_09578_),
    .X(_00861_));
 sky130_fd_sc_hd__and2_1 _17196_ (.A(_09521_),
    .B(_09522_),
    .X(_09579_));
 sky130_fd_sc_hd__o21ai_2 _17197_ (.A1(_09523_),
    .A2(_09579_),
    .B1(\wfg_stim_sine_top.wfg_stim_sine.quadrant[1] ),
    .Y(_09580_));
 sky130_fd_sc_hd__o221a_2 _17198_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[8] ),
    .A2(_09553_),
    .B1(_09565_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.x[8] ),
    .C1(_09554_),
    .X(_09581_));
 sky130_fd_sc_hd__a22o_1 _17199_ (.A1(_06748_),
    .A2(_09549_),
    .B1(_09580_),
    .B2(_09581_),
    .X(_00860_));
 sky130_fd_sc_hd__or2_1 _17200_ (.A(_09518_),
    .B(_09520_),
    .X(_09582_));
 sky130_fd_sc_hd__a21o_1 _17201_ (.A1(_09521_),
    .A2(_09582_),
    .B1(_09556_),
    .X(_09583_));
 sky130_fd_sc_hd__o221a_2 _17202_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[7] ),
    .A2(_09553_),
    .B1(_09565_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.x[7] ),
    .C1(_09554_),
    .X(_09584_));
 sky130_fd_sc_hd__a22o_1 _17203_ (.A1(_06754_),
    .A2(_09549_),
    .B1(_09583_),
    .B2(_09584_),
    .X(_00859_));
 sky130_fd_sc_hd__and2_1 _17204_ (.A(_09515_),
    .B(_09517_),
    .X(_09585_));
 sky130_fd_sc_hd__o21ai_2 _17205_ (.A1(_09518_),
    .A2(_09585_),
    .B1(\wfg_stim_sine_top.wfg_stim_sine.quadrant[1] ),
    .Y(_09586_));
 sky130_fd_sc_hd__o221a_2 _17206_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[6] ),
    .A2(_09553_),
    .B1(_09565_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.x[6] ),
    .C1(_09554_),
    .X(_09587_));
 sky130_fd_sc_hd__a22o_1 _17207_ (.A1(_06742_),
    .A2(_09549_),
    .B1(_09586_),
    .B2(_09587_),
    .X(_00858_));
 sky130_fd_sc_hd__nand2_1 _17208_ (.A(_09513_),
    .B(_09514_),
    .Y(_09588_));
 sky130_fd_sc_hd__a21o_1 _17209_ (.A1(_09515_),
    .A2(_09588_),
    .B1(_09556_),
    .X(_09589_));
 sky130_fd_sc_hd__o221a_2 _17210_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[5] ),
    .A2(_09552_),
    .B1(_09565_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.x[5] ),
    .C1(_09545_),
    .X(_09590_));
 sky130_fd_sc_hd__a22o_1 _17211_ (.A1(_06752_),
    .A2(_09548_),
    .B1(_09589_),
    .B2(_09590_),
    .X(_00857_));
 sky130_fd_sc_hd__nand2_1 _17212_ (.A(_09511_),
    .B(_09512_),
    .Y(_09591_));
 sky130_fd_sc_hd__a21o_1 _17213_ (.A1(_09513_),
    .A2(_09591_),
    .B1(_09556_),
    .X(_09592_));
 sky130_fd_sc_hd__o221a_2 _17214_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[4] ),
    .A2(_09552_),
    .B1(_09565_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.x[4] ),
    .C1(_09545_),
    .X(_09593_));
 sky130_fd_sc_hd__a22o_1 _17215_ (.A1(_07007_),
    .A2(_09548_),
    .B1(_09592_),
    .B2(_09593_),
    .X(_00856_));
 sky130_fd_sc_hd__nand2_1 _17216_ (.A(_09509_),
    .B(_09510_),
    .Y(_09594_));
 sky130_fd_sc_hd__a21o_1 _17217_ (.A1(_09511_),
    .A2(_09594_),
    .B1(_09556_),
    .X(_09595_));
 sky130_fd_sc_hd__o221a_1 _17218_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[3] ),
    .A2(_09552_),
    .B1(_09564_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.x[3] ),
    .C1(_09545_),
    .X(_09596_));
 sky130_fd_sc_hd__a22o_1 _17219_ (.A1(_06996_),
    .A2(_09548_),
    .B1(_09595_),
    .B2(_09596_),
    .X(_00855_));
 sky130_fd_sc_hd__nand2_1 _17220_ (.A(_09507_),
    .B(_09508_),
    .Y(_09597_));
 sky130_fd_sc_hd__a21o_1 _17221_ (.A1(_09509_),
    .A2(_09597_),
    .B1(_09556_),
    .X(_09598_));
 sky130_fd_sc_hd__o221a_2 _17222_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[2] ),
    .A2(_09552_),
    .B1(_09564_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.x[2] ),
    .C1(_09545_),
    .X(_09599_));
 sky130_fd_sc_hd__a22o_1 _17223_ (.A1(_06972_),
    .A2(_09548_),
    .B1(_09598_),
    .B2(_09599_),
    .X(_00854_));
 sky130_fd_sc_hd__nand2_1 _17224_ (.A(_09505_),
    .B(_09506_),
    .Y(_09600_));
 sky130_fd_sc_hd__a21o_1 _17225_ (.A1(_09507_),
    .A2(_09600_),
    .B1(_09556_),
    .X(_09601_));
 sky130_fd_sc_hd__o221a_1 _17226_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.y[1] ),
    .A2(_09552_),
    .B1(_09564_),
    .B2(\wfg_stim_sine_top.wfg_stim_sine.x[1] ),
    .C1(_09545_),
    .X(_09602_));
 sky130_fd_sc_hd__a22o_1 _17227_ (.A1(_07493_),
    .A2(_09548_),
    .B1(_09601_),
    .B2(_09602_),
    .X(_00853_));
 sky130_fd_sc_hd__mux2_2 _17228_ (.A0(\wfg_stim_sine_top.wfg_stim_sine.y[0] ),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.x[0] ),
    .S(\wfg_stim_sine_top.wfg_stim_sine.quadrant[0] ),
    .X(_09603_));
 sky130_fd_sc_hd__mux2_1 _17229_ (.A0(_07689_),
    .A1(_09603_),
    .S(_09545_),
    .X(_09604_));
 sky130_fd_sc_hd__clkbuf_1 _17230_ (.A(_09604_),
    .X(_00852_));
 sky130_fd_sc_hd__nor2_2 _17231_ (.A(_06356_),
    .B(_06360_),
    .Y(_09605_));
 sky130_fd_sc_hd__or3b_1 _17232_ (.A(\wfg_stim_sine_top.wfg_stim_sine.cur_state[1] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.cur_state[0] ),
    .C_N(\wfg_stim_sine_top.wfg_stim_sine.cur_state[2] ),
    .X(_09606_));
 sky130_fd_sc_hd__buf_4 _17233_ (.A(_09606_),
    .X(_09607_));
 sky130_fd_sc_hd__buf_4 _17234_ (.A(_09607_),
    .X(_09608_));
 sky130_fd_sc_hd__or3b_1 _17235_ (.A(_08773_),
    .B(_09605_),
    .C_N(_09608_),
    .X(_09609_));
 sky130_fd_sc_hd__clkbuf_1 _17236_ (.A(_09609_),
    .X(_00850_));
 sky130_fd_sc_hd__inv_2 _17237_ (.A(\wfg_stim_sine_top.ctrl_en_q ),
    .Y(_09610_));
 sky130_fd_sc_hd__a211o_1 _17238_ (.A1(_09610_),
    .A2(_09056_),
    .B1(_09605_),
    .C1(_08907_),
    .X(_09611_));
 sky130_fd_sc_hd__a21oi_1 _17239_ (.A1(_08916_),
    .A2(_09548_),
    .B1(_09611_),
    .Y(_00849_));
 sky130_fd_sc_hd__a21oi_1 _17240_ (.A1(\wfg_stim_sine_top.wfg_stim_sine.cur_state[2] ),
    .A2(\wfg_stim_sine_top.wfg_stim_sine.cur_state[1] ),
    .B1(\wfg_stim_sine_top.wfg_stim_sine.cur_state[0] ),
    .Y(_09612_));
 sky130_fd_sc_hd__o22a_1 _17241_ (.A1(\wfg_stim_sine_top.ctrl_en_q ),
    .A2(_08924_),
    .B1(_09611_),
    .B2(_09612_),
    .X(_00848_));
 sky130_fd_sc_hd__nand2_1 _17242_ (.A(_09479_),
    .B(_09477_),
    .Y(_09613_));
 sky130_fd_sc_hd__nor2_1 _17243_ (.A(\wfg_stim_sine_top.offset_val_q[16] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[30] ),
    .Y(_09614_));
 sky130_fd_sc_hd__nor2_1 _17244_ (.A(\wfg_stim_sine_top.offset_val_q[14] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[28] ),
    .Y(_09615_));
 sky130_fd_sc_hd__nor2_1 _17245_ (.A(\wfg_stim_sine_top.offset_val_q[12] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[26] ),
    .Y(_09616_));
 sky130_fd_sc_hd__nor2_1 _17246_ (.A(\wfg_stim_sine_top.offset_val_q[10] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[24] ),
    .Y(_09617_));
 sky130_fd_sc_hd__nor2_1 _17247_ (.A(\wfg_stim_sine_top.offset_val_q[8] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[22] ),
    .Y(_09618_));
 sky130_fd_sc_hd__nor2_1 _17248_ (.A(\wfg_stim_sine_top.offset_val_q[7] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[21] ),
    .Y(_09619_));
 sky130_fd_sc_hd__nor2_1 _17249_ (.A(\wfg_stim_sine_top.offset_val_q[6] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[20] ),
    .Y(_09620_));
 sky130_fd_sc_hd__nor2_1 _17250_ (.A(\wfg_stim_sine_top.offset_val_q[5] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[19] ),
    .Y(_09621_));
 sky130_fd_sc_hd__or2_1 _17251_ (.A(\wfg_stim_sine_top.offset_val_q[4] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[18] ),
    .X(_09622_));
 sky130_fd_sc_hd__nor2_1 _17252_ (.A(\wfg_stim_sine_top.offset_val_q[2] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[16] ),
    .Y(_09623_));
 sky130_fd_sc_hd__nor2_1 _17253_ (.A(\wfg_stim_sine_top.offset_val_q[1] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[15] ),
    .Y(_09624_));
 sky130_fd_sc_hd__nand2_1 _17254_ (.A(\wfg_stim_sine_top.offset_val_q[0] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[14] ),
    .Y(_09625_));
 sky130_fd_sc_hd__and2_1 _17255_ (.A(\wfg_stim_sine_top.offset_val_q[1] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[15] ),
    .X(_09626_));
 sky130_fd_sc_hd__o21ba_1 _17256_ (.A1(_09624_),
    .A2(_09625_),
    .B1_N(_09626_),
    .X(_09627_));
 sky130_fd_sc_hd__nand2_1 _17257_ (.A(\wfg_stim_sine_top.offset_val_q[2] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[16] ),
    .Y(_09628_));
 sky130_fd_sc_hd__o21ai_1 _17258_ (.A1(_09623_),
    .A2(_09627_),
    .B1(_09628_),
    .Y(_09629_));
 sky130_fd_sc_hd__a21o_1 _17259_ (.A1(\wfg_stim_sine_top.offset_val_q[3] ),
    .A2(\wfg_stim_sine_top.wfg_stim_sine.temp[17] ),
    .B1(_09629_),
    .X(_09630_));
 sky130_fd_sc_hd__o21a_1 _17260_ (.A1(\wfg_stim_sine_top.offset_val_q[3] ),
    .A2(\wfg_stim_sine_top.wfg_stim_sine.temp[17] ),
    .B1(_09630_),
    .X(_09631_));
 sky130_fd_sc_hd__and2_1 _17261_ (.A(\wfg_stim_sine_top.offset_val_q[4] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[18] ),
    .X(_09632_));
 sky130_fd_sc_hd__a21oi_1 _17262_ (.A1(_09622_),
    .A2(_09631_),
    .B1(_09632_),
    .Y(_09633_));
 sky130_fd_sc_hd__and2_1 _17263_ (.A(\wfg_stim_sine_top.offset_val_q[5] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[19] ),
    .X(_09634_));
 sky130_fd_sc_hd__o21ba_1 _17264_ (.A1(_09621_),
    .A2(_09633_),
    .B1_N(_09634_),
    .X(_09635_));
 sky130_fd_sc_hd__nand2_1 _17265_ (.A(\wfg_stim_sine_top.offset_val_q[6] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[20] ),
    .Y(_09636_));
 sky130_fd_sc_hd__o21a_1 _17266_ (.A1(_09620_),
    .A2(_09635_),
    .B1(_09636_),
    .X(_09637_));
 sky130_fd_sc_hd__nand2_1 _17267_ (.A(\wfg_stim_sine_top.offset_val_q[7] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[21] ),
    .Y(_09638_));
 sky130_fd_sc_hd__o21a_1 _17268_ (.A1(_09619_),
    .A2(_09637_),
    .B1(_09638_),
    .X(_09639_));
 sky130_fd_sc_hd__nand2_1 _17269_ (.A(\wfg_stim_sine_top.offset_val_q[8] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[22] ),
    .Y(_09640_));
 sky130_fd_sc_hd__o21ai_1 _17270_ (.A1(_09618_),
    .A2(_09639_),
    .B1(_09640_),
    .Y(_09641_));
 sky130_fd_sc_hd__a21o_1 _17271_ (.A1(\wfg_stim_sine_top.offset_val_q[9] ),
    .A2(\wfg_stim_sine_top.wfg_stim_sine.temp[23] ),
    .B1(_09641_),
    .X(_09642_));
 sky130_fd_sc_hd__o21ai_1 _17272_ (.A1(\wfg_stim_sine_top.offset_val_q[9] ),
    .A2(\wfg_stim_sine_top.wfg_stim_sine.temp[23] ),
    .B1(_09642_),
    .Y(_09643_));
 sky130_fd_sc_hd__nand2_1 _17273_ (.A(\wfg_stim_sine_top.offset_val_q[10] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[24] ),
    .Y(_09644_));
 sky130_fd_sc_hd__o21ai_1 _17274_ (.A1(_09617_),
    .A2(_09643_),
    .B1(_09644_),
    .Y(_09645_));
 sky130_fd_sc_hd__a21o_1 _17275_ (.A1(\wfg_stim_sine_top.offset_val_q[11] ),
    .A2(\wfg_stim_sine_top.wfg_stim_sine.temp[25] ),
    .B1(_09645_),
    .X(_09646_));
 sky130_fd_sc_hd__o21ai_1 _17276_ (.A1(\wfg_stim_sine_top.offset_val_q[11] ),
    .A2(\wfg_stim_sine_top.wfg_stim_sine.temp[25] ),
    .B1(_09646_),
    .Y(_09647_));
 sky130_fd_sc_hd__nand2_1 _17277_ (.A(\wfg_stim_sine_top.offset_val_q[12] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[26] ),
    .Y(_09648_));
 sky130_fd_sc_hd__o21ai_1 _17278_ (.A1(_09616_),
    .A2(_09647_),
    .B1(_09648_),
    .Y(_09649_));
 sky130_fd_sc_hd__a21o_1 _17279_ (.A1(\wfg_stim_sine_top.offset_val_q[13] ),
    .A2(\wfg_stim_sine_top.wfg_stim_sine.temp[27] ),
    .B1(_09649_),
    .X(_09650_));
 sky130_fd_sc_hd__o21ai_1 _17280_ (.A1(\wfg_stim_sine_top.offset_val_q[13] ),
    .A2(\wfg_stim_sine_top.wfg_stim_sine.temp[27] ),
    .B1(_09650_),
    .Y(_09651_));
 sky130_fd_sc_hd__nand2_1 _17281_ (.A(\wfg_stim_sine_top.offset_val_q[14] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[28] ),
    .Y(_09652_));
 sky130_fd_sc_hd__o21ai_1 _17282_ (.A1(_09615_),
    .A2(_09651_),
    .B1(_09652_),
    .Y(_09653_));
 sky130_fd_sc_hd__a21o_1 _17283_ (.A1(\wfg_stim_sine_top.offset_val_q[15] ),
    .A2(\wfg_stim_sine_top.wfg_stim_sine.temp[29] ),
    .B1(_09653_),
    .X(_09654_));
 sky130_fd_sc_hd__o21ai_1 _17284_ (.A1(\wfg_stim_sine_top.offset_val_q[15] ),
    .A2(\wfg_stim_sine_top.wfg_stim_sine.temp[29] ),
    .B1(_09654_),
    .Y(_09655_));
 sky130_fd_sc_hd__and2_1 _17285_ (.A(\wfg_stim_sine_top.offset_val_q[16] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[30] ),
    .X(_09656_));
 sky130_fd_sc_hd__o21bai_1 _17286_ (.A1(_09614_),
    .A2(_09655_),
    .B1_N(_09656_),
    .Y(_09657_));
 sky130_fd_sc_hd__xnor2_1 _17287_ (.A(_09613_),
    .B(_09657_),
    .Y(_09658_));
 sky130_fd_sc_hd__mux2_1 _17288_ (.A0(_09658_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[17] ),
    .S(_09608_),
    .X(_09659_));
 sky130_fd_sc_hd__clkbuf_1 _17289_ (.A(_09659_),
    .X(_00847_));
 sky130_fd_sc_hd__nor2_1 _17290_ (.A(_09656_),
    .B(_09614_),
    .Y(_09660_));
 sky130_fd_sc_hd__xnor2_1 _17291_ (.A(_09660_),
    .B(_09655_),
    .Y(_09661_));
 sky130_fd_sc_hd__mux2_1 _17292_ (.A0(_09661_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[16] ),
    .S(_09608_),
    .X(_09662_));
 sky130_fd_sc_hd__clkbuf_1 _17293_ (.A(_09662_),
    .X(_00846_));
 sky130_fd_sc_hd__xnor2_1 _17294_ (.A(\wfg_stim_sine_top.offset_val_q[15] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[29] ),
    .Y(_09663_));
 sky130_fd_sc_hd__xnor2_1 _17295_ (.A(_09653_),
    .B(_09663_),
    .Y(_09664_));
 sky130_fd_sc_hd__mux2_1 _17296_ (.A0(_09664_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[15] ),
    .S(_09608_),
    .X(_09665_));
 sky130_fd_sc_hd__clkbuf_1 _17297_ (.A(_09665_),
    .X(_00845_));
 sky130_fd_sc_hd__and2b_1 _17298_ (.A_N(_09615_),
    .B(_09652_),
    .X(_09666_));
 sky130_fd_sc_hd__xnor2_1 _17299_ (.A(_09651_),
    .B(_09666_),
    .Y(_09667_));
 sky130_fd_sc_hd__mux2_1 _17300_ (.A0(_09667_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[14] ),
    .S(_09608_),
    .X(_09668_));
 sky130_fd_sc_hd__clkbuf_1 _17301_ (.A(_09668_),
    .X(_00844_));
 sky130_fd_sc_hd__xnor2_1 _17302_ (.A(\wfg_stim_sine_top.offset_val_q[13] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[27] ),
    .Y(_09669_));
 sky130_fd_sc_hd__xnor2_1 _17303_ (.A(_09649_),
    .B(_09669_),
    .Y(_09670_));
 sky130_fd_sc_hd__mux2_1 _17304_ (.A0(_09670_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[13] ),
    .S(_09608_),
    .X(_09671_));
 sky130_fd_sc_hd__clkbuf_1 _17305_ (.A(_09671_),
    .X(_00843_));
 sky130_fd_sc_hd__and2b_1 _17306_ (.A_N(_09616_),
    .B(_09648_),
    .X(_09672_));
 sky130_fd_sc_hd__xnor2_1 _17307_ (.A(_09647_),
    .B(_09672_),
    .Y(_09673_));
 sky130_fd_sc_hd__mux2_1 _17308_ (.A0(_09673_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[12] ),
    .S(_09608_),
    .X(_09674_));
 sky130_fd_sc_hd__clkbuf_1 _17309_ (.A(_09674_),
    .X(_00842_));
 sky130_fd_sc_hd__xnor2_1 _17310_ (.A(\wfg_stim_sine_top.offset_val_q[11] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[25] ),
    .Y(_09675_));
 sky130_fd_sc_hd__xnor2_1 _17311_ (.A(_09645_),
    .B(_09675_),
    .Y(_09676_));
 sky130_fd_sc_hd__mux2_1 _17312_ (.A0(_09676_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[11] ),
    .S(_09608_),
    .X(_09677_));
 sky130_fd_sc_hd__clkbuf_1 _17313_ (.A(_09677_),
    .X(_00841_));
 sky130_fd_sc_hd__and2b_1 _17314_ (.A_N(_09617_),
    .B(_09644_),
    .X(_09678_));
 sky130_fd_sc_hd__xnor2_1 _17315_ (.A(_09643_),
    .B(_09678_),
    .Y(_09679_));
 sky130_fd_sc_hd__mux2_1 _17316_ (.A0(_09679_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[10] ),
    .S(_09608_),
    .X(_09680_));
 sky130_fd_sc_hd__clkbuf_1 _17317_ (.A(_09680_),
    .X(_00840_));
 sky130_fd_sc_hd__xnor2_1 _17318_ (.A(\wfg_stim_sine_top.offset_val_q[9] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[23] ),
    .Y(_09681_));
 sky130_fd_sc_hd__xnor2_1 _17319_ (.A(_09641_),
    .B(_09681_),
    .Y(_09682_));
 sky130_fd_sc_hd__mux2_1 _17320_ (.A0(_09682_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[9] ),
    .S(_09608_),
    .X(_09683_));
 sky130_fd_sc_hd__clkbuf_1 _17321_ (.A(_09683_),
    .X(_00839_));
 sky130_fd_sc_hd__and2b_1 _17322_ (.A_N(_09618_),
    .B(_09640_),
    .X(_09684_));
 sky130_fd_sc_hd__xnor2_1 _17323_ (.A(_09639_),
    .B(_09684_),
    .Y(_09685_));
 sky130_fd_sc_hd__mux2_1 _17324_ (.A0(_09685_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[8] ),
    .S(_09607_),
    .X(_09686_));
 sky130_fd_sc_hd__clkbuf_1 _17325_ (.A(_09686_),
    .X(_00838_));
 sky130_fd_sc_hd__and2b_1 _17326_ (.A_N(_09619_),
    .B(_09638_),
    .X(_09687_));
 sky130_fd_sc_hd__xnor2_1 _17327_ (.A(_09637_),
    .B(_09687_),
    .Y(_09688_));
 sky130_fd_sc_hd__mux2_1 _17328_ (.A0(_09688_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[7] ),
    .S(_09607_),
    .X(_09689_));
 sky130_fd_sc_hd__clkbuf_1 _17329_ (.A(_09689_),
    .X(_00837_));
 sky130_fd_sc_hd__and2b_1 _17330_ (.A_N(_09620_),
    .B(_09636_),
    .X(_09690_));
 sky130_fd_sc_hd__xnor2_1 _17331_ (.A(_09635_),
    .B(_09690_),
    .Y(_09691_));
 sky130_fd_sc_hd__mux2_1 _17332_ (.A0(_09691_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[6] ),
    .S(_09607_),
    .X(_09692_));
 sky130_fd_sc_hd__clkbuf_1 _17333_ (.A(_09692_),
    .X(_00836_));
 sky130_fd_sc_hd__nor2_1 _17334_ (.A(_09634_),
    .B(_09621_),
    .Y(_09693_));
 sky130_fd_sc_hd__xnor2_1 _17335_ (.A(_09693_),
    .B(_09633_),
    .Y(_09694_));
 sky130_fd_sc_hd__mux2_1 _17336_ (.A0(_09694_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[5] ),
    .S(_09607_),
    .X(_09695_));
 sky130_fd_sc_hd__clkbuf_1 _17337_ (.A(_09695_),
    .X(_00835_));
 sky130_fd_sc_hd__or2b_1 _17338_ (.A(_09632_),
    .B_N(_09622_),
    .X(_09696_));
 sky130_fd_sc_hd__xnor2_1 _17339_ (.A(_09696_),
    .B(_09631_),
    .Y(_09697_));
 sky130_fd_sc_hd__mux2_1 _17340_ (.A0(_09697_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[4] ),
    .S(_09607_),
    .X(_09698_));
 sky130_fd_sc_hd__clkbuf_1 _17341_ (.A(_09698_),
    .X(_00834_));
 sky130_fd_sc_hd__xnor2_1 _17342_ (.A(\wfg_stim_sine_top.offset_val_q[3] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[17] ),
    .Y(_09699_));
 sky130_fd_sc_hd__xnor2_1 _17343_ (.A(_09629_),
    .B(_09699_),
    .Y(_09700_));
 sky130_fd_sc_hd__mux2_1 _17344_ (.A0(_09700_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[3] ),
    .S(_09607_),
    .X(_09701_));
 sky130_fd_sc_hd__clkbuf_1 _17345_ (.A(_09701_),
    .X(_00833_));
 sky130_fd_sc_hd__or2b_1 _17346_ (.A(_09623_),
    .B_N(_09628_),
    .X(_09702_));
 sky130_fd_sc_hd__xor2_1 _17347_ (.A(_09627_),
    .B(_09702_),
    .X(_09703_));
 sky130_fd_sc_hd__mux2_1 _17348_ (.A0(_09703_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[2] ),
    .S(_09607_),
    .X(_09704_));
 sky130_fd_sc_hd__clkbuf_1 _17349_ (.A(_09704_),
    .X(_00832_));
 sky130_fd_sc_hd__nor2_1 _17350_ (.A(_09626_),
    .B(_09624_),
    .Y(_09705_));
 sky130_fd_sc_hd__xnor2_1 _17351_ (.A(_09705_),
    .B(_09625_),
    .Y(_09706_));
 sky130_fd_sc_hd__mux2_1 _17352_ (.A0(_09706_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[1] ),
    .S(_09607_),
    .X(_09707_));
 sky130_fd_sc_hd__clkbuf_1 _17353_ (.A(_09707_),
    .X(_00831_));
 sky130_fd_sc_hd__or2_1 _17354_ (.A(\wfg_stim_sine_top.offset_val_q[0] ),
    .B(\wfg_stim_sine_top.wfg_stim_sine.temp[14] ),
    .X(_09708_));
 sky130_fd_sc_hd__and2_1 _17355_ (.A(_09625_),
    .B(_09708_),
    .X(_09709_));
 sky130_fd_sc_hd__mux2_1 _17356_ (.A0(_09709_),
    .A1(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[0] ),
    .S(_09607_),
    .X(_09710_));
 sky130_fd_sc_hd__clkbuf_1 _17357_ (.A(_09710_),
    .X(_00830_));
 sky130_fd_sc_hd__nor2b_2 _17358_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_dly ),
    .B_N(\wfg_subcore_top.wfg_subcore.temp_subcycle ),
    .Y(_09711_));
 sky130_fd_sc_hd__clkinv_2 _17359_ (.A(\wfg_subcore_top.active_o ),
    .Y(_09712_));
 sky130_fd_sc_hd__nor2_2 _17360_ (.A(_09712_),
    .B(_02709_),
    .Y(_09713_));
 sky130_fd_sc_hd__and3_1 _17361_ (.A(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[2] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[1] ),
    .C(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[0] ),
    .X(_09714_));
 sky130_fd_sc_hd__and3_1 _17362_ (.A(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[4] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[3] ),
    .C(_09714_),
    .X(_09715_));
 sky130_fd_sc_hd__and3_1 _17363_ (.A(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[6] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[5] ),
    .C(_09715_),
    .X(_09716_));
 sky130_fd_sc_hd__and3_1 _17364_ (.A(_09711_),
    .B(_09713_),
    .C(_09716_),
    .X(_09717_));
 sky130_fd_sc_hd__a21boi_1 _17365_ (.A1(_09711_),
    .A2(_09716_),
    .B1_N(_09713_),
    .Y(_09718_));
 sky130_fd_sc_hd__mux2_1 _17366_ (.A0(_09717_),
    .A1(_09718_),
    .S(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[7] ),
    .X(_09719_));
 sky130_fd_sc_hd__clkbuf_1 _17367_ (.A(_09719_),
    .X(_00772_));
 sky130_fd_sc_hd__a31o_1 _17368_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[5] ),
    .A2(_09715_),
    .A3(_09711_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[6] ),
    .X(_09720_));
 sky130_fd_sc_hd__and2_1 _17369_ (.A(_09718_),
    .B(_09720_),
    .X(_09721_));
 sky130_fd_sc_hd__clkbuf_1 _17370_ (.A(_09721_),
    .X(_00771_));
 sky130_fd_sc_hd__nand2_1 _17371_ (.A(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[5] ),
    .B(_09715_),
    .Y(_09722_));
 sky130_fd_sc_hd__or2b_1 _17372_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_dly ),
    .B_N(\wfg_subcore_top.wfg_subcore.temp_subcycle ),
    .X(_09723_));
 sky130_fd_sc_hd__and2_1 _17373_ (.A(_09715_),
    .B(_09711_),
    .X(_09724_));
 sky130_fd_sc_hd__o221a_1 _17374_ (.A1(_09722_),
    .A2(_09723_),
    .B1(_09724_),
    .B2(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[5] ),
    .C1(_09713_),
    .X(_00770_));
 sky130_fd_sc_hd__a31o_1 _17375_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[3] ),
    .A2(_09714_),
    .A3(_09711_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[4] ),
    .X(_09725_));
 sky130_fd_sc_hd__and3b_1 _17376_ (.A_N(_09724_),
    .B(_09725_),
    .C(_09713_),
    .X(_09726_));
 sky130_fd_sc_hd__clkbuf_1 _17377_ (.A(_09726_),
    .X(_00769_));
 sky130_fd_sc_hd__and2_1 _17378_ (.A(_09714_),
    .B(_09711_),
    .X(_09727_));
 sky130_fd_sc_hd__a21boi_1 _17379_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[3] ),
    .A2(_09727_),
    .B1_N(_09713_),
    .Y(_09728_));
 sky130_fd_sc_hd__o21a_1 _17380_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[3] ),
    .A2(_09727_),
    .B1(_09728_),
    .X(_00768_));
 sky130_fd_sc_hd__a31o_1 _17381_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[1] ),
    .A2(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[0] ),
    .A3(_09711_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[2] ),
    .X(_09729_));
 sky130_fd_sc_hd__and3b_1 _17382_ (.A_N(_09727_),
    .B(_09729_),
    .C(_09713_),
    .X(_09730_));
 sky130_fd_sc_hd__clkbuf_1 _17383_ (.A(_09730_),
    .X(_00767_));
 sky130_fd_sc_hd__nand2_1 _17384_ (.A(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[1] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[0] ),
    .Y(_09731_));
 sky130_fd_sc_hd__a21o_1 _17385_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[0] ),
    .A2(_09711_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[1] ),
    .X(_09732_));
 sky130_fd_sc_hd__o211a_1 _17386_ (.A1(_09731_),
    .A2(_09723_),
    .B1(_09713_),
    .C1(_09732_),
    .X(_00766_));
 sky130_fd_sc_hd__a211o_1 _17387_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[0] ),
    .A2(_09711_),
    .B1(_02709_),
    .C1(_09712_),
    .X(_09733_));
 sky130_fd_sc_hd__o21ba_1 _17388_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[0] ),
    .A2(_09711_),
    .B1_N(_09733_),
    .X(_00765_));
 sky130_fd_sc_hd__or3_1 _17389_ (.A(\wfg_subcore_top.wfg_subcore.sync_count[2] ),
    .B(\wfg_subcore_top.wfg_subcore.sync_count[1] ),
    .C(\wfg_subcore_top.wfg_subcore.sync_count[0] ),
    .X(_09734_));
 sky130_fd_sc_hd__or2_1 _17390_ (.A(\wfg_subcore_top.wfg_subcore.sync_count[3] ),
    .B(_09734_),
    .X(_09735_));
 sky130_fd_sc_hd__or3_1 _17391_ (.A(\wfg_subcore_top.wfg_subcore.sync_count[5] ),
    .B(\wfg_subcore_top.wfg_subcore.sync_count[4] ),
    .C(_09735_),
    .X(_09736_));
 sky130_fd_sc_hd__or2_1 _17392_ (.A(\wfg_subcore_top.wfg_subcore.sync_count[6] ),
    .B(_09736_),
    .X(_09737_));
 sky130_fd_sc_hd__or2_1 _17393_ (.A(\wfg_subcore_top.wfg_subcore.sync_count[7] ),
    .B(_09737_),
    .X(_09738_));
 sky130_fd_sc_hd__buf_2 _17394_ (.A(_09738_),
    .X(_09739_));
 sky130_fd_sc_hd__or3_1 _17395_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_count[2] ),
    .B(\wfg_subcore_top.wfg_subcore.subcycle_count[1] ),
    .C(\wfg_subcore_top.wfg_subcore.subcycle_count[0] ),
    .X(_09740_));
 sky130_fd_sc_hd__or2_2 _17396_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_count[3] ),
    .B(_09740_),
    .X(_09741_));
 sky130_fd_sc_hd__or3_1 _17397_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_count[5] ),
    .B(\wfg_subcore_top.wfg_subcore.subcycle_count[4] ),
    .C(_09741_),
    .X(_09742_));
 sky130_fd_sc_hd__or2_1 _17398_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_count[6] ),
    .B(_09742_),
    .X(_09743_));
 sky130_fd_sc_hd__or3_1 _17399_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_count[8] ),
    .B(\wfg_subcore_top.wfg_subcore.subcycle_count[7] ),
    .C(_09743_),
    .X(_09744_));
 sky130_fd_sc_hd__or2_1 _17400_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_count[9] ),
    .B(_09744_),
    .X(_09745_));
 sky130_fd_sc_hd__or3_1 _17401_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_count[11] ),
    .B(\wfg_subcore_top.wfg_subcore.subcycle_count[10] ),
    .C(_09745_),
    .X(_09746_));
 sky130_fd_sc_hd__or2_1 _17402_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_count[12] ),
    .B(_09746_),
    .X(_09747_));
 sky130_fd_sc_hd__or2_1 _17403_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_count[13] ),
    .B(_09747_),
    .X(_09748_));
 sky130_fd_sc_hd__or2_1 _17404_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_count[14] ),
    .B(_09748_),
    .X(_09749_));
 sky130_fd_sc_hd__or2_1 _17405_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_count[15] ),
    .B(_09749_),
    .X(_09750_));
 sky130_fd_sc_hd__buf_2 _17406_ (.A(_09750_),
    .X(_09751_));
 sky130_fd_sc_hd__nor2_1 _17407_ (.A(_09739_),
    .B(_09751_),
    .Y(_09752_));
 sky130_fd_sc_hd__o21ai_1 _17408_ (.A1(\wfg_subcore_top.wfg_subcore.temp_sync ),
    .A2(_09752_),
    .B1(\wfg_subcore_top.active_o ),
    .Y(_09753_));
 sky130_fd_sc_hd__a21oi_1 _17409_ (.A1(\wfg_subcore_top.wfg_subcore.temp_sync ),
    .A2(_09752_),
    .B1(_09753_),
    .Y(_00762_));
 sky130_fd_sc_hd__nor2_4 _17410_ (.A(_09712_),
    .B(_09751_),
    .Y(_09754_));
 sky130_fd_sc_hd__and2_1 _17411_ (.A(\wfg_subcore_top.active_o ),
    .B(_09751_),
    .X(_09755_));
 sky130_fd_sc_hd__buf_2 _17412_ (.A(_09755_),
    .X(_09756_));
 sky130_fd_sc_hd__mux2_1 _17413_ (.A0(_09754_),
    .A1(_09756_),
    .S(\wfg_subcore_top.wfg_subcore.temp_subcycle ),
    .X(_09757_));
 sky130_fd_sc_hd__clkbuf_1 _17414_ (.A(_09757_),
    .X(_00761_));
 sky130_fd_sc_hd__inv_2 _17415_ (.A(\wfg_subcore_top.cfg_sync_q[7] ),
    .Y(_09758_));
 sky130_fd_sc_hd__nand2_1 _17416_ (.A(\wfg_subcore_top.wfg_subcore.sync_count[7] ),
    .B(_09737_),
    .Y(_09759_));
 sky130_fd_sc_hd__o21ai_1 _17417_ (.A1(_09758_),
    .A2(_09739_),
    .B1(_09759_),
    .Y(_09760_));
 sky130_fd_sc_hd__a22o_1 _17418_ (.A1(\wfg_subcore_top.wfg_subcore.sync_count[7] ),
    .A2(_09756_),
    .B1(_09754_),
    .B2(_09760_),
    .X(_00760_));
 sky130_fd_sc_hd__nand2_1 _17419_ (.A(\wfg_subcore_top.wfg_subcore.sync_count[6] ),
    .B(_09736_),
    .Y(_09761_));
 sky130_fd_sc_hd__o2bb2a_1 _17420_ (.A1_N(_09737_),
    .A2_N(_09761_),
    .B1(_09739_),
    .B2(\wfg_subcore_top.cfg_sync_q[6] ),
    .X(_09762_));
 sky130_fd_sc_hd__a22o_1 _17421_ (.A1(\wfg_subcore_top.wfg_subcore.sync_count[6] ),
    .A2(_09756_),
    .B1(_09754_),
    .B2(_09762_),
    .X(_00759_));
 sky130_fd_sc_hd__o21ai_1 _17422_ (.A1(\wfg_subcore_top.wfg_subcore.sync_count[4] ),
    .A2(_09735_),
    .B1(\wfg_subcore_top.wfg_subcore.sync_count[5] ),
    .Y(_09763_));
 sky130_fd_sc_hd__o2bb2a_1 _17423_ (.A1_N(_09736_),
    .A2_N(_09763_),
    .B1(_09739_),
    .B2(\wfg_subcore_top.cfg_sync_q[5] ),
    .X(_09764_));
 sky130_fd_sc_hd__a22o_1 _17424_ (.A1(\wfg_subcore_top.wfg_subcore.sync_count[5] ),
    .A2(_09756_),
    .B1(_09754_),
    .B2(_09764_),
    .X(_00758_));
 sky130_fd_sc_hd__or2_1 _17425_ (.A(\wfg_subcore_top.cfg_sync_q[4] ),
    .B(_09739_),
    .X(_09765_));
 sky130_fd_sc_hd__xnor2_1 _17426_ (.A(\wfg_subcore_top.wfg_subcore.sync_count[4] ),
    .B(_09735_),
    .Y(_09766_));
 sky130_fd_sc_hd__a32o_1 _17427_ (.A1(_09754_),
    .A2(_09765_),
    .A3(_09766_),
    .B1(_09756_),
    .B2(\wfg_subcore_top.wfg_subcore.sync_count[4] ),
    .X(_00757_));
 sky130_fd_sc_hd__nand2_1 _17428_ (.A(\wfg_subcore_top.wfg_subcore.sync_count[3] ),
    .B(_09734_),
    .Y(_09767_));
 sky130_fd_sc_hd__o2bb2a_1 _17429_ (.A1_N(_09735_),
    .A2_N(_09767_),
    .B1(_09739_),
    .B2(\wfg_subcore_top.cfg_sync_q[3] ),
    .X(_09768_));
 sky130_fd_sc_hd__a22o_1 _17430_ (.A1(\wfg_subcore_top.wfg_subcore.sync_count[3] ),
    .A2(_09756_),
    .B1(_09754_),
    .B2(_09768_),
    .X(_00756_));
 sky130_fd_sc_hd__o21ai_1 _17431_ (.A1(\wfg_subcore_top.wfg_subcore.sync_count[1] ),
    .A2(\wfg_subcore_top.wfg_subcore.sync_count[0] ),
    .B1(\wfg_subcore_top.wfg_subcore.sync_count[2] ),
    .Y(_09769_));
 sky130_fd_sc_hd__o2bb2a_1 _17432_ (.A1_N(_09734_),
    .A2_N(_09769_),
    .B1(_09739_),
    .B2(\wfg_subcore_top.cfg_sync_q[2] ),
    .X(_09770_));
 sky130_fd_sc_hd__a22o_1 _17433_ (.A1(\wfg_subcore_top.wfg_subcore.sync_count[2] ),
    .A2(_09756_),
    .B1(_09754_),
    .B2(_09770_),
    .X(_00755_));
 sky130_fd_sc_hd__and2_1 _17434_ (.A(\wfg_subcore_top.wfg_subcore.sync_count[1] ),
    .B(\wfg_subcore_top.wfg_subcore.sync_count[0] ),
    .X(_09771_));
 sky130_fd_sc_hd__nor2_1 _17435_ (.A(\wfg_subcore_top.wfg_subcore.sync_count[1] ),
    .B(\wfg_subcore_top.wfg_subcore.sync_count[0] ),
    .Y(_09772_));
 sky130_fd_sc_hd__o22a_1 _17436_ (.A1(\wfg_subcore_top.cfg_sync_q[1] ),
    .A2(_09739_),
    .B1(_09771_),
    .B2(_09772_),
    .X(_09773_));
 sky130_fd_sc_hd__a22o_1 _17437_ (.A1(\wfg_subcore_top.wfg_subcore.sync_count[1] ),
    .A2(_09756_),
    .B1(_09754_),
    .B2(_09773_),
    .X(_00754_));
 sky130_fd_sc_hd__o21ba_1 _17438_ (.A1(\wfg_subcore_top.cfg_sync_q[0] ),
    .A2(_09739_),
    .B1_N(\wfg_subcore_top.wfg_subcore.sync_count[0] ),
    .X(_09774_));
 sky130_fd_sc_hd__a22o_1 _17439_ (.A1(\wfg_subcore_top.wfg_subcore.sync_count[0] ),
    .A2(_09756_),
    .B1(_09754_),
    .B2(_09774_),
    .X(_00753_));
 sky130_fd_sc_hd__inv_2 _17440_ (.A(\wfg_drive_pat_top.cfg_end_q[13] ),
    .Y(_09775_));
 sky130_fd_sc_hd__mux2_1 _17441_ (.A0(\wfg_core_top.wfg_core.subcycle_pls_cnt[5] ),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[5] ),
    .S(\wfg_drive_pat_top.cfg_core_sel_q ),
    .X(_09776_));
 sky130_fd_sc_hd__mux2_1 _17442_ (.A0(\wfg_core_top.wfg_core.subcycle_pls_cnt[7] ),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[7] ),
    .S(\wfg_drive_pat_top.cfg_core_sel_q ),
    .X(_09777_));
 sky130_fd_sc_hd__inv_2 _17443_ (.A(\wfg_drive_pat_top.cfg_end_q[15] ),
    .Y(_09778_));
 sky130_fd_sc_hd__mux2_1 _17444_ (.A0(\wfg_core_top.wfg_core.subcycle_pls_cnt[2] ),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[2] ),
    .S(\wfg_drive_pat_top.cfg_core_sel_q ),
    .X(_09779_));
 sky130_fd_sc_hd__xor2_1 _17445_ (.A(\wfg_drive_pat_top.cfg_end_q[10] ),
    .B(_09779_),
    .X(_09780_));
 sky130_fd_sc_hd__a221o_1 _17446_ (.A1(_09775_),
    .A2(_09776_),
    .B1(_09777_),
    .B2(_09778_),
    .C1(_09780_),
    .X(_09781_));
 sky130_fd_sc_hd__buf_4 _17447_ (.A(\wfg_drive_pat_top.cfg_core_sel_q ),
    .X(_09782_));
 sky130_fd_sc_hd__or2b_1 _17448_ (.A(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[1] ),
    .B_N(\wfg_drive_pat_top.cfg_core_sel_q ),
    .X(_09783_));
 sky130_fd_sc_hd__o21ai_2 _17449_ (.A1(_09782_),
    .A2(\wfg_core_top.wfg_core.subcycle_pls_cnt[1] ),
    .B1(_09783_),
    .Y(_09784_));
 sky130_fd_sc_hd__xnor2_1 _17450_ (.A(\wfg_drive_pat_top.cfg_end_q[9] ),
    .B(_09784_),
    .Y(_09785_));
 sky130_fd_sc_hd__inv_2 _17451_ (.A(_09776_),
    .Y(_09786_));
 sky130_fd_sc_hd__or2b_1 _17452_ (.A(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[3] ),
    .B_N(_09782_),
    .X(_09787_));
 sky130_fd_sc_hd__o21ai_2 _17453_ (.A1(_09782_),
    .A2(\wfg_core_top.wfg_core.subcycle_pls_cnt[3] ),
    .B1(_09787_),
    .Y(_09788_));
 sky130_fd_sc_hd__a22o_1 _17454_ (.A1(\wfg_drive_pat_top.cfg_end_q[13] ),
    .A2(_09786_),
    .B1(_09788_),
    .B2(\wfg_drive_pat_top.cfg_end_q[11] ),
    .X(_09789_));
 sky130_fd_sc_hd__or3_1 _17455_ (.A(_09781_),
    .B(_09785_),
    .C(_09789_),
    .X(_09790_));
 sky130_fd_sc_hd__clkbuf_4 _17456_ (.A(_09790_),
    .X(_09791_));
 sky130_fd_sc_hd__mux2_1 _17457_ (.A0(\wfg_core_top.wfg_core.subcycle_pls_cnt[0] ),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[0] ),
    .S(_09782_),
    .X(_09792_));
 sky130_fd_sc_hd__inv_2 _17458_ (.A(\wfg_drive_pat_top.cfg_end_q[8] ),
    .Y(_09793_));
 sky130_fd_sc_hd__or2b_1 _17459_ (.A(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[4] ),
    .B_N(_09782_),
    .X(_09794_));
 sky130_fd_sc_hd__o21ai_2 _17460_ (.A1(_09782_),
    .A2(\wfg_core_top.wfg_core.subcycle_pls_cnt[4] ),
    .B1(_09794_),
    .Y(_09795_));
 sky130_fd_sc_hd__a22oi_1 _17461_ (.A1(_09793_),
    .A2(_09792_),
    .B1(_09795_),
    .B2(\wfg_drive_pat_top.cfg_end_q[12] ),
    .Y(_09796_));
 sky130_fd_sc_hd__o221a_1 _17462_ (.A1(\wfg_drive_pat_top.cfg_end_q[11] ),
    .A2(_09788_),
    .B1(_09792_),
    .B2(_09793_),
    .C1(_09796_),
    .X(_09797_));
 sky130_fd_sc_hd__mux2_1 _17463_ (.A0(\wfg_core_top.wfg_core.subcycle_pls_cnt[6] ),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[6] ),
    .S(_09782_),
    .X(_09798_));
 sky130_fd_sc_hd__xnor2_1 _17464_ (.A(\wfg_drive_pat_top.cfg_end_q[14] ),
    .B(_09798_),
    .Y(_09799_));
 sky130_fd_sc_hd__o221a_1 _17465_ (.A1(_09778_),
    .A2(_09777_),
    .B1(_09795_),
    .B2(\wfg_drive_pat_top.cfg_end_q[12] ),
    .C1(_09799_),
    .X(_09800_));
 sky130_fd_sc_hd__nand2_4 _17466_ (.A(_09797_),
    .B(_09800_),
    .Y(_09801_));
 sky130_fd_sc_hd__nor2_1 _17467_ (.A(_09791_),
    .B(_09801_),
    .Y(_09802_));
 sky130_fd_sc_hd__buf_4 _17468_ (.A(_09802_),
    .X(_09803_));
 sky130_fd_sc_hd__clkbuf_4 _17469_ (.A(_09803_),
    .X(_09804_));
 sky130_fd_sc_hd__clkbuf_4 _17470_ (.A(_09804_),
    .X(_09805_));
 sky130_fd_sc_hd__nand2_1 _17471_ (.A(\wfg_drive_pat_top.patsel1_high_q[9] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[9].drv.axis_data_ff ),
    .Y(_09806_));
 sky130_fd_sc_hd__clkbuf_4 _17472_ (.A(_09801_),
    .X(_09807_));
 sky130_fd_sc_hd__clkbuf_4 _17473_ (.A(_09791_),
    .X(_09808_));
 sky130_fd_sc_hd__a211o_1 _17474_ (.A1(\wfg_drive_pat_top.patsel0_low_q[9] ),
    .A2(_09806_),
    .B1(_09807_),
    .C1(_09808_),
    .X(_09809_));
 sky130_fd_sc_hd__o211a_1 _17475_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[9].drv.axis_data_ff ),
    .A2(_09805_),
    .B1(_09809_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[9].drv.ctrl_en_q_i ),
    .X(_09810_));
 sky130_fd_sc_hd__inv_2 _17476_ (.A(\wfg_drive_pat_top.cfg_begin_q[7] ),
    .Y(_09811_));
 sky130_fd_sc_hd__a2bb2o_1 _17477_ (.A1_N(_09788_),
    .A2_N(\wfg_drive_pat_top.cfg_begin_q[3] ),
    .B1(_09811_),
    .B2(_09777_),
    .X(_09812_));
 sky130_fd_sc_hd__a2bb2o_1 _17478_ (.A1_N(\wfg_drive_pat_top.cfg_begin_q[5] ),
    .A2_N(_09786_),
    .B1(_09788_),
    .B2(\wfg_drive_pat_top.cfg_begin_q[3] ),
    .X(_09813_));
 sky130_fd_sc_hd__inv_2 _17479_ (.A(\wfg_drive_pat_top.cfg_begin_q[0] ),
    .Y(_09814_));
 sky130_fd_sc_hd__inv_2 _17480_ (.A(\wfg_drive_pat_top.cfg_begin_q[6] ),
    .Y(_09815_));
 sky130_fd_sc_hd__a22o_1 _17481_ (.A1(_09814_),
    .A2(_09792_),
    .B1(_09798_),
    .B2(_09815_),
    .X(_09816_));
 sky130_fd_sc_hd__a221o_1 _17482_ (.A1(\wfg_drive_pat_top.cfg_begin_q[5] ),
    .A2(_09786_),
    .B1(_09795_),
    .B2(\wfg_drive_pat_top.cfg_begin_q[4] ),
    .C1(_09816_),
    .X(_09817_));
 sky130_fd_sc_hd__nor3_2 _17483_ (.A(_09812_),
    .B(_09813_),
    .C(_09817_),
    .Y(_09818_));
 sky130_fd_sc_hd__or2_1 _17484_ (.A(\wfg_drive_pat_top.cfg_begin_q[1] ),
    .B(_09784_),
    .X(_09819_));
 sky130_fd_sc_hd__nand2_1 _17485_ (.A(\wfg_drive_pat_top.cfg_begin_q[1] ),
    .B(_09784_),
    .Y(_09820_));
 sky130_fd_sc_hd__xnor2_1 _17486_ (.A(\wfg_drive_pat_top.cfg_begin_q[2] ),
    .B(_09779_),
    .Y(_09821_));
 sky130_fd_sc_hd__o22a_1 _17487_ (.A1(_09814_),
    .A2(_09792_),
    .B1(_09798_),
    .B2(_09815_),
    .X(_09822_));
 sky130_fd_sc_hd__o221a_1 _17488_ (.A1(_09811_),
    .A2(_09777_),
    .B1(_09795_),
    .B2(\wfg_drive_pat_top.cfg_begin_q[4] ),
    .C1(_09822_),
    .X(_09823_));
 sky130_fd_sc_hd__and4_1 _17489_ (.A(_09819_),
    .B(_09820_),
    .C(_09821_),
    .D(_09823_),
    .X(_09824_));
 sky130_fd_sc_hd__a21oi_4 _17490_ (.A1(_09818_),
    .A2(_09824_),
    .B1(_09803_),
    .Y(_09825_));
 sky130_fd_sc_hd__clkbuf_4 _17491_ (.A(_09825_),
    .X(_09826_));
 sky130_fd_sc_hd__and3b_1 _17492_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[9] ),
    .B(_09804_),
    .C(\wfg_drive_pat_top.patsel1_high_q[9] ),
    .X(_09827_));
 sky130_fd_sc_hd__o21a_1 _17493_ (.A1(_09826_),
    .A2(_09827_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[9].drv.ctrl_en_q_i ),
    .X(_09828_));
 sky130_fd_sc_hd__mux2_1 _17494_ (.A0(_09810_),
    .A1(net176),
    .S(_09828_),
    .X(_09829_));
 sky130_fd_sc_hd__clkbuf_1 _17495_ (.A(_09829_),
    .X(_00606_));
 sky130_fd_sc_hd__nand2_1 _17496_ (.A(\wfg_drive_pat_top.patsel1_high_q[30] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[30].drv.axis_data_ff ),
    .Y(_09830_));
 sky130_fd_sc_hd__a211o_1 _17497_ (.A1(\wfg_drive_pat_top.patsel0_low_q[30] ),
    .A2(_09830_),
    .B1(_09807_),
    .C1(_09808_),
    .X(_09831_));
 sky130_fd_sc_hd__o211a_1 _17498_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[30].drv.axis_data_ff ),
    .A2(_09805_),
    .B1(_09831_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[30].drv.ctrl_en_q_i ),
    .X(_09832_));
 sky130_fd_sc_hd__and3b_1 _17499_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[30] ),
    .B(_09804_),
    .C(\wfg_drive_pat_top.patsel1_high_q[30] ),
    .X(_09833_));
 sky130_fd_sc_hd__o21a_1 _17500_ (.A1(_09826_),
    .A2(_09833_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[30].drv.ctrl_en_q_i ),
    .X(_09834_));
 sky130_fd_sc_hd__mux2_1 _17501_ (.A0(_09832_),
    .A1(net168),
    .S(_09834_),
    .X(_09835_));
 sky130_fd_sc_hd__clkbuf_1 _17502_ (.A(_09835_),
    .X(_00605_));
 sky130_fd_sc_hd__nand2_1 _17503_ (.A(\wfg_drive_pat_top.patsel1_high_q[2] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[2].drv.axis_data_ff ),
    .Y(_09836_));
 sky130_fd_sc_hd__a211o_1 _17504_ (.A1(\wfg_drive_pat_top.patsel0_low_q[2] ),
    .A2(_09836_),
    .B1(_09807_),
    .C1(_09808_),
    .X(_09837_));
 sky130_fd_sc_hd__o211a_1 _17505_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[2].drv.axis_data_ff ),
    .A2(_09805_),
    .B1(_09837_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[2].drv.ctrl_en_q_i ),
    .X(_09838_));
 sky130_fd_sc_hd__and3b_1 _17506_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[2] ),
    .B(_09804_),
    .C(\wfg_drive_pat_top.patsel1_high_q[2] ),
    .X(_09839_));
 sky130_fd_sc_hd__o21a_1 _17507_ (.A1(_09826_),
    .A2(_09839_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[2].drv.ctrl_en_q_i ),
    .X(_09840_));
 sky130_fd_sc_hd__mux2_1 _17508_ (.A0(_09838_),
    .A1(net167),
    .S(_09840_),
    .X(_09841_));
 sky130_fd_sc_hd__clkbuf_1 _17509_ (.A(_09841_),
    .X(_00604_));
 sky130_fd_sc_hd__nand2_1 _17510_ (.A(\wfg_drive_pat_top.patsel1_high_q[28] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[28].drv.axis_data_ff ),
    .Y(_09842_));
 sky130_fd_sc_hd__a211o_1 _17511_ (.A1(\wfg_drive_pat_top.patsel0_low_q[28] ),
    .A2(_09842_),
    .B1(_09807_),
    .C1(_09808_),
    .X(_09843_));
 sky130_fd_sc_hd__o211a_1 _17512_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[28].drv.axis_data_ff ),
    .A2(_09805_),
    .B1(_09843_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[28].drv.ctrl_en_q_i ),
    .X(_09844_));
 sky130_fd_sc_hd__and3b_1 _17513_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[28] ),
    .B(_09804_),
    .C(\wfg_drive_pat_top.patsel1_high_q[28] ),
    .X(_09845_));
 sky130_fd_sc_hd__o21a_1 _17514_ (.A1(_09826_),
    .A2(_09845_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[28].drv.ctrl_en_q_i ),
    .X(_09846_));
 sky130_fd_sc_hd__mux2_1 _17515_ (.A0(_09844_),
    .A1(net165),
    .S(_09846_),
    .X(_09847_));
 sky130_fd_sc_hd__clkbuf_1 _17516_ (.A(_09847_),
    .X(_00603_));
 sky130_fd_sc_hd__nand2_1 _17517_ (.A(\wfg_drive_pat_top.patsel1_high_q[27] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[27].drv.axis_data_ff ),
    .Y(_09848_));
 sky130_fd_sc_hd__a211o_1 _17518_ (.A1(\wfg_drive_pat_top.patsel0_low_q[27] ),
    .A2(_09848_),
    .B1(_09807_),
    .C1(_09808_),
    .X(_09849_));
 sky130_fd_sc_hd__o211a_1 _17519_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[27].drv.axis_data_ff ),
    .A2(_09805_),
    .B1(_09849_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[27].drv.ctrl_en_q_i ),
    .X(_09850_));
 sky130_fd_sc_hd__and3b_1 _17520_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[27] ),
    .B(_09804_),
    .C(\wfg_drive_pat_top.patsel1_high_q[27] ),
    .X(_09851_));
 sky130_fd_sc_hd__o21a_1 _17521_ (.A1(_09826_),
    .A2(_09851_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[27].drv.ctrl_en_q_i ),
    .X(_09852_));
 sky130_fd_sc_hd__mux2_1 _17522_ (.A0(_09850_),
    .A1(net164),
    .S(_09852_),
    .X(_09853_));
 sky130_fd_sc_hd__clkbuf_1 _17523_ (.A(_09853_),
    .X(_00602_));
 sky130_fd_sc_hd__nand2_1 _17524_ (.A(\wfg_drive_pat_top.patsel1_high_q[26] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[26].drv.axis_data_ff ),
    .Y(_09854_));
 sky130_fd_sc_hd__a211o_1 _17525_ (.A1(\wfg_drive_pat_top.patsel0_low_q[26] ),
    .A2(_09854_),
    .B1(_09807_),
    .C1(_09808_),
    .X(_09855_));
 sky130_fd_sc_hd__o211a_1 _17526_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[26].drv.axis_data_ff ),
    .A2(_09805_),
    .B1(_09855_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[26].drv.ctrl_en_q_i ),
    .X(_09856_));
 sky130_fd_sc_hd__clkbuf_4 _17527_ (.A(_09803_),
    .X(_09857_));
 sky130_fd_sc_hd__and3b_1 _17528_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[26] ),
    .B(_09857_),
    .C(\wfg_drive_pat_top.patsel1_high_q[26] ),
    .X(_09858_));
 sky130_fd_sc_hd__o21a_1 _17529_ (.A1(_09826_),
    .A2(_09858_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[26].drv.ctrl_en_q_i ),
    .X(_09859_));
 sky130_fd_sc_hd__mux2_1 _17530_ (.A0(_09856_),
    .A1(net163),
    .S(_09859_),
    .X(_09860_));
 sky130_fd_sc_hd__clkbuf_1 _17531_ (.A(_09860_),
    .X(_00601_));
 sky130_fd_sc_hd__nand2_1 _17532_ (.A(\wfg_drive_pat_top.patsel1_high_q[25] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[25].drv.axis_data_ff ),
    .Y(_09861_));
 sky130_fd_sc_hd__a211o_1 _17533_ (.A1(\wfg_drive_pat_top.patsel0_low_q[25] ),
    .A2(_09861_),
    .B1(_09807_),
    .C1(_09808_),
    .X(_09862_));
 sky130_fd_sc_hd__o211a_1 _17534_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[25].drv.axis_data_ff ),
    .A2(_09805_),
    .B1(_09862_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[25].drv.ctrl_en_q_i ),
    .X(_09863_));
 sky130_fd_sc_hd__and3b_1 _17535_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[25] ),
    .B(_09857_),
    .C(\wfg_drive_pat_top.patsel1_high_q[25] ),
    .X(_09864_));
 sky130_fd_sc_hd__o21a_1 _17536_ (.A1(_09826_),
    .A2(_09864_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[25].drv.ctrl_en_q_i ),
    .X(_09865_));
 sky130_fd_sc_hd__mux2_1 _17537_ (.A0(_09863_),
    .A1(net162),
    .S(_09865_),
    .X(_09866_));
 sky130_fd_sc_hd__clkbuf_1 _17538_ (.A(_09866_),
    .X(_00600_));
 sky130_fd_sc_hd__nand2_1 _17539_ (.A(\wfg_drive_pat_top.patsel1_high_q[24] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[24].drv.axis_data_ff ),
    .Y(_09867_));
 sky130_fd_sc_hd__a211o_1 _17540_ (.A1(\wfg_drive_pat_top.patsel0_low_q[24] ),
    .A2(_09867_),
    .B1(_09807_),
    .C1(_09808_),
    .X(_09868_));
 sky130_fd_sc_hd__o211a_1 _17541_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[24].drv.axis_data_ff ),
    .A2(_09805_),
    .B1(_09868_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[24].drv.ctrl_en_q_i ),
    .X(_09869_));
 sky130_fd_sc_hd__and3b_1 _17542_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[24] ),
    .B(_09857_),
    .C(\wfg_drive_pat_top.patsel1_high_q[24] ),
    .X(_09870_));
 sky130_fd_sc_hd__o21a_1 _17543_ (.A1(_09826_),
    .A2(_09870_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[24].drv.ctrl_en_q_i ),
    .X(_09871_));
 sky130_fd_sc_hd__mux2_1 _17544_ (.A0(_09869_),
    .A1(net161),
    .S(_09871_),
    .X(_09872_));
 sky130_fd_sc_hd__clkbuf_1 _17545_ (.A(_09872_),
    .X(_00599_));
 sky130_fd_sc_hd__nand2_1 _17546_ (.A(\wfg_drive_pat_top.patsel1_high_q[23] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[23].drv.axis_data_ff ),
    .Y(_09873_));
 sky130_fd_sc_hd__a211o_1 _17547_ (.A1(\wfg_drive_pat_top.patsel0_low_q[23] ),
    .A2(_09873_),
    .B1(_09807_),
    .C1(_09808_),
    .X(_09874_));
 sky130_fd_sc_hd__o211a_1 _17548_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[23].drv.axis_data_ff ),
    .A2(_09805_),
    .B1(_09874_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[23].drv.ctrl_en_q_i ),
    .X(_09875_));
 sky130_fd_sc_hd__and3b_1 _17549_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[23] ),
    .B(_09857_),
    .C(\wfg_drive_pat_top.patsel1_high_q[23] ),
    .X(_09876_));
 sky130_fd_sc_hd__o21a_1 _17550_ (.A1(_09826_),
    .A2(_09876_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[23].drv.ctrl_en_q_i ),
    .X(_09877_));
 sky130_fd_sc_hd__mux2_1 _17551_ (.A0(_09875_),
    .A1(net160),
    .S(_09877_),
    .X(_09878_));
 sky130_fd_sc_hd__clkbuf_1 _17552_ (.A(_09878_),
    .X(_00598_));
 sky130_fd_sc_hd__nand2_1 _17553_ (.A(\wfg_drive_pat_top.patsel1_high_q[22] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[22].drv.axis_data_ff ),
    .Y(_09879_));
 sky130_fd_sc_hd__a211o_1 _17554_ (.A1(\wfg_drive_pat_top.patsel0_low_q[22] ),
    .A2(_09879_),
    .B1(_09807_),
    .C1(_09808_),
    .X(_09880_));
 sky130_fd_sc_hd__o211a_1 _17555_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[22].drv.axis_data_ff ),
    .A2(_09805_),
    .B1(_09880_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[22].drv.ctrl_en_q_i ),
    .X(_09881_));
 sky130_fd_sc_hd__and3b_1 _17556_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[22] ),
    .B(_09857_),
    .C(\wfg_drive_pat_top.patsel1_high_q[22] ),
    .X(_09882_));
 sky130_fd_sc_hd__o21a_1 _17557_ (.A1(_09826_),
    .A2(_09882_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[22].drv.ctrl_en_q_i ),
    .X(_09883_));
 sky130_fd_sc_hd__mux2_1 _17558_ (.A0(_09881_),
    .A1(net159),
    .S(_09883_),
    .X(_09884_));
 sky130_fd_sc_hd__clkbuf_1 _17559_ (.A(_09884_),
    .X(_00597_));
 sky130_fd_sc_hd__clkbuf_4 _17560_ (.A(_09804_),
    .X(_09885_));
 sky130_fd_sc_hd__nand2_1 _17561_ (.A(\wfg_drive_pat_top.patsel1_high_q[21] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[21].drv.axis_data_ff ),
    .Y(_09886_));
 sky130_fd_sc_hd__clkbuf_4 _17562_ (.A(_09801_),
    .X(_09887_));
 sky130_fd_sc_hd__clkbuf_4 _17563_ (.A(_09791_),
    .X(_09888_));
 sky130_fd_sc_hd__a211o_1 _17564_ (.A1(\wfg_drive_pat_top.patsel0_low_q[21] ),
    .A2(_09886_),
    .B1(_09887_),
    .C1(_09888_),
    .X(_09889_));
 sky130_fd_sc_hd__o211a_1 _17565_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[21].drv.axis_data_ff ),
    .A2(_09885_),
    .B1(_09889_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[21].drv.ctrl_en_q_i ),
    .X(_09890_));
 sky130_fd_sc_hd__clkbuf_4 _17566_ (.A(_09825_),
    .X(_09891_));
 sky130_fd_sc_hd__and3b_1 _17567_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[21] ),
    .B(_09857_),
    .C(\wfg_drive_pat_top.patsel1_high_q[21] ),
    .X(_09892_));
 sky130_fd_sc_hd__o21a_1 _17568_ (.A1(_09891_),
    .A2(_09892_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[21].drv.ctrl_en_q_i ),
    .X(_09893_));
 sky130_fd_sc_hd__mux2_1 _17569_ (.A0(_09890_),
    .A1(net158),
    .S(_09893_),
    .X(_09894_));
 sky130_fd_sc_hd__clkbuf_1 _17570_ (.A(_09894_),
    .X(_00596_));
 sky130_fd_sc_hd__nand2_1 _17571_ (.A(\wfg_drive_pat_top.patsel1_high_q[20] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[20].drv.axis_data_ff ),
    .Y(_09895_));
 sky130_fd_sc_hd__a211o_1 _17572_ (.A1(\wfg_drive_pat_top.patsel0_low_q[20] ),
    .A2(_09895_),
    .B1(_09887_),
    .C1(_09888_),
    .X(_09896_));
 sky130_fd_sc_hd__o211a_1 _17573_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[20].drv.axis_data_ff ),
    .A2(_09885_),
    .B1(_09896_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[20].drv.ctrl_en_q_i ),
    .X(_09897_));
 sky130_fd_sc_hd__and3b_1 _17574_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[20] ),
    .B(_09857_),
    .C(\wfg_drive_pat_top.patsel1_high_q[20] ),
    .X(_09898_));
 sky130_fd_sc_hd__o21a_1 _17575_ (.A1(_09891_),
    .A2(_09898_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[20].drv.ctrl_en_q_i ),
    .X(_09899_));
 sky130_fd_sc_hd__mux2_1 _17576_ (.A0(_09897_),
    .A1(net157),
    .S(_09899_),
    .X(_09900_));
 sky130_fd_sc_hd__clkbuf_1 _17577_ (.A(_09900_),
    .X(_00595_));
 sky130_fd_sc_hd__nand2_1 _17578_ (.A(\wfg_drive_pat_top.patsel1_high_q[1] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[1].drv.axis_data_ff ),
    .Y(_09901_));
 sky130_fd_sc_hd__a211o_1 _17579_ (.A1(\wfg_drive_pat_top.patsel0_low_q[1] ),
    .A2(_09901_),
    .B1(_09887_),
    .C1(_09888_),
    .X(_09902_));
 sky130_fd_sc_hd__o211a_1 _17580_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[1].drv.axis_data_ff ),
    .A2(_09885_),
    .B1(_09902_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[1].drv.ctrl_en_q_i ),
    .X(_09903_));
 sky130_fd_sc_hd__and3b_1 _17581_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[1] ),
    .B(_09857_),
    .C(\wfg_drive_pat_top.patsel1_high_q[1] ),
    .X(_09904_));
 sky130_fd_sc_hd__o21a_1 _17582_ (.A1(_09891_),
    .A2(_09904_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[1].drv.ctrl_en_q_i ),
    .X(_09905_));
 sky130_fd_sc_hd__mux2_1 _17583_ (.A0(_09903_),
    .A1(net156),
    .S(_09905_),
    .X(_09906_));
 sky130_fd_sc_hd__clkbuf_1 _17584_ (.A(_09906_),
    .X(_00594_));
 sky130_fd_sc_hd__nand2_1 _17585_ (.A(\wfg_drive_pat_top.patsel1_high_q[18] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[18].drv.axis_data_ff ),
    .Y(_09907_));
 sky130_fd_sc_hd__a211o_1 _17586_ (.A1(\wfg_drive_pat_top.patsel0_low_q[18] ),
    .A2(_09907_),
    .B1(_09887_),
    .C1(_09888_),
    .X(_09908_));
 sky130_fd_sc_hd__o211a_1 _17587_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[18].drv.axis_data_ff ),
    .A2(_09885_),
    .B1(_09908_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[18].drv.ctrl_en_q_i ),
    .X(_09909_));
 sky130_fd_sc_hd__and3b_1 _17588_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[18] ),
    .B(_09857_),
    .C(\wfg_drive_pat_top.patsel1_high_q[18] ),
    .X(_09910_));
 sky130_fd_sc_hd__o21a_1 _17589_ (.A1(_09891_),
    .A2(_09910_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[18].drv.ctrl_en_q_i ),
    .X(_09911_));
 sky130_fd_sc_hd__mux2_1 _17590_ (.A0(_09909_),
    .A1(net154),
    .S(_09911_),
    .X(_09912_));
 sky130_fd_sc_hd__clkbuf_1 _17591_ (.A(_09912_),
    .X(_00593_));
 sky130_fd_sc_hd__nand2_1 _17592_ (.A(\wfg_drive_pat_top.patsel1_high_q[17] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[17].drv.axis_data_ff ),
    .Y(_09913_));
 sky130_fd_sc_hd__a211o_1 _17593_ (.A1(\wfg_drive_pat_top.patsel0_low_q[17] ),
    .A2(_09913_),
    .B1(_09887_),
    .C1(_09888_),
    .X(_09914_));
 sky130_fd_sc_hd__o211a_1 _17594_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[17].drv.axis_data_ff ),
    .A2(_09885_),
    .B1(_09914_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[17].drv.ctrl_en_q_i ),
    .X(_09915_));
 sky130_fd_sc_hd__and3b_1 _17595_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[17] ),
    .B(_09857_),
    .C(\wfg_drive_pat_top.patsel1_high_q[17] ),
    .X(_09916_));
 sky130_fd_sc_hd__o21a_1 _17596_ (.A1(_09891_),
    .A2(_09916_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[17].drv.ctrl_en_q_i ),
    .X(_09917_));
 sky130_fd_sc_hd__mux2_1 _17597_ (.A0(_09915_),
    .A1(net153),
    .S(_09917_),
    .X(_09918_));
 sky130_fd_sc_hd__clkbuf_1 _17598_ (.A(_09918_),
    .X(_00592_));
 sky130_fd_sc_hd__nand2_1 _17599_ (.A(\wfg_drive_pat_top.patsel1_high_q[16] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[16].drv.axis_data_ff ),
    .Y(_09919_));
 sky130_fd_sc_hd__a211o_1 _17600_ (.A1(\wfg_drive_pat_top.patsel0_low_q[16] ),
    .A2(_09919_),
    .B1(_09887_),
    .C1(_09888_),
    .X(_09920_));
 sky130_fd_sc_hd__o211a_1 _17601_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[16].drv.axis_data_ff ),
    .A2(_09885_),
    .B1(_09920_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[16].drv.ctrl_en_q_i ),
    .X(_09921_));
 sky130_fd_sc_hd__buf_2 _17602_ (.A(_09802_),
    .X(_09922_));
 sky130_fd_sc_hd__and3b_1 _17603_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[16] ),
    .B(_09922_),
    .C(\wfg_drive_pat_top.patsel1_high_q[16] ),
    .X(_09923_));
 sky130_fd_sc_hd__o21a_1 _17604_ (.A1(_09891_),
    .A2(_09923_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[16].drv.ctrl_en_q_i ),
    .X(_09924_));
 sky130_fd_sc_hd__mux2_1 _17605_ (.A0(_09921_),
    .A1(net152),
    .S(_09924_),
    .X(_09925_));
 sky130_fd_sc_hd__clkbuf_1 _17606_ (.A(_09925_),
    .X(_00591_));
 sky130_fd_sc_hd__nand2_1 _17607_ (.A(\wfg_drive_pat_top.patsel1_high_q[15] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[15].drv.axis_data_ff ),
    .Y(_09926_));
 sky130_fd_sc_hd__a211o_1 _17608_ (.A1(\wfg_drive_pat_top.patsel0_low_q[15] ),
    .A2(_09926_),
    .B1(_09887_),
    .C1(_09888_),
    .X(_09927_));
 sky130_fd_sc_hd__o211a_1 _17609_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[15].drv.axis_data_ff ),
    .A2(_09885_),
    .B1(_09927_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[15].drv.ctrl_en_q_i ),
    .X(_09928_));
 sky130_fd_sc_hd__and3b_1 _17610_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[15] ),
    .B(_09922_),
    .C(\wfg_drive_pat_top.patsel1_high_q[15] ),
    .X(_09929_));
 sky130_fd_sc_hd__o21a_1 _17611_ (.A1(_09891_),
    .A2(_09929_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[15].drv.ctrl_en_q_i ),
    .X(_09930_));
 sky130_fd_sc_hd__mux2_1 _17612_ (.A0(_09928_),
    .A1(net151),
    .S(_09930_),
    .X(_09931_));
 sky130_fd_sc_hd__clkbuf_1 _17613_ (.A(_09931_),
    .X(_00590_));
 sky130_fd_sc_hd__nand2_1 _17614_ (.A(\wfg_drive_pat_top.patsel1_high_q[14] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[14].drv.axis_data_ff ),
    .Y(_09932_));
 sky130_fd_sc_hd__a211o_1 _17615_ (.A1(\wfg_drive_pat_top.patsel0_low_q[14] ),
    .A2(_09932_),
    .B1(_09887_),
    .C1(_09888_),
    .X(_09933_));
 sky130_fd_sc_hd__o211a_1 _17616_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[14].drv.axis_data_ff ),
    .A2(_09885_),
    .B1(_09933_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[14].drv.ctrl_en_q_i ),
    .X(_09934_));
 sky130_fd_sc_hd__and3b_1 _17617_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[14] ),
    .B(_09922_),
    .C(\wfg_drive_pat_top.patsel1_high_q[14] ),
    .X(_09935_));
 sky130_fd_sc_hd__o21a_1 _17618_ (.A1(_09891_),
    .A2(_09935_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[14].drv.ctrl_en_q_i ),
    .X(_09936_));
 sky130_fd_sc_hd__mux2_1 _17619_ (.A0(_09934_),
    .A1(net150),
    .S(_09936_),
    .X(_09937_));
 sky130_fd_sc_hd__clkbuf_1 _17620_ (.A(_09937_),
    .X(_00589_));
 sky130_fd_sc_hd__nand2_1 _17621_ (.A(\wfg_drive_pat_top.patsel1_high_q[13] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[13].drv.axis_data_ff ),
    .Y(_09938_));
 sky130_fd_sc_hd__a211o_1 _17622_ (.A1(\wfg_drive_pat_top.patsel0_low_q[13] ),
    .A2(_09938_),
    .B1(_09887_),
    .C1(_09888_),
    .X(_09939_));
 sky130_fd_sc_hd__o211a_1 _17623_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[13].drv.axis_data_ff ),
    .A2(_09885_),
    .B1(_09939_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[13].drv.ctrl_en_q_i ),
    .X(_09940_));
 sky130_fd_sc_hd__and3b_1 _17624_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[13] ),
    .B(_09922_),
    .C(\wfg_drive_pat_top.patsel1_high_q[13] ),
    .X(_09941_));
 sky130_fd_sc_hd__o21a_1 _17625_ (.A1(_09891_),
    .A2(_09941_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[13].drv.ctrl_en_q_i ),
    .X(_09942_));
 sky130_fd_sc_hd__mux2_1 _17626_ (.A0(_09940_),
    .A1(net149),
    .S(_09942_),
    .X(_09943_));
 sky130_fd_sc_hd__clkbuf_1 _17627_ (.A(_09943_),
    .X(_00564_));
 sky130_fd_sc_hd__nand2_1 _17628_ (.A(\wfg_drive_pat_top.patsel1_high_q[12] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[12].drv.axis_data_ff ),
    .Y(_09944_));
 sky130_fd_sc_hd__a211o_1 _17629_ (.A1(\wfg_drive_pat_top.patsel0_low_q[12] ),
    .A2(_09944_),
    .B1(_09887_),
    .C1(_09888_),
    .X(_09945_));
 sky130_fd_sc_hd__o211a_1 _17630_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[12].drv.axis_data_ff ),
    .A2(_09885_),
    .B1(_09945_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[12].drv.ctrl_en_q_i ),
    .X(_09946_));
 sky130_fd_sc_hd__and3b_1 _17631_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[12] ),
    .B(_09922_),
    .C(\wfg_drive_pat_top.patsel1_high_q[12] ),
    .X(_09947_));
 sky130_fd_sc_hd__o21a_1 _17632_ (.A1(_09891_),
    .A2(_09947_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[12].drv.ctrl_en_q_i ),
    .X(_09948_));
 sky130_fd_sc_hd__mux2_1 _17633_ (.A0(_09946_),
    .A1(net148),
    .S(_09948_),
    .X(_09949_));
 sky130_fd_sc_hd__clkbuf_1 _17634_ (.A(_09949_),
    .X(_00563_));
 sky130_fd_sc_hd__buf_4 _17635_ (.A(_09804_),
    .X(_09950_));
 sky130_fd_sc_hd__nand2_1 _17636_ (.A(\wfg_drive_pat_top.patsel1_high_q[11] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[11].drv.axis_data_ff ),
    .Y(_09951_));
 sky130_fd_sc_hd__buf_4 _17637_ (.A(_09801_),
    .X(_09952_));
 sky130_fd_sc_hd__buf_4 _17638_ (.A(_09791_),
    .X(_09953_));
 sky130_fd_sc_hd__a211o_1 _17639_ (.A1(\wfg_drive_pat_top.patsel0_low_q[11] ),
    .A2(_09951_),
    .B1(_09952_),
    .C1(_09953_),
    .X(_09954_));
 sky130_fd_sc_hd__o211a_1 _17640_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[11].drv.axis_data_ff ),
    .A2(_09950_),
    .B1(_09954_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[11].drv.ctrl_en_q_i ),
    .X(_09955_));
 sky130_fd_sc_hd__buf_4 _17641_ (.A(_09825_),
    .X(_09956_));
 sky130_fd_sc_hd__and3b_1 _17642_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[11] ),
    .B(_09922_),
    .C(\wfg_drive_pat_top.patsel1_high_q[11] ),
    .X(_09957_));
 sky130_fd_sc_hd__o21a_1 _17643_ (.A1(_09956_),
    .A2(_09957_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[11].drv.ctrl_en_q_i ),
    .X(_09958_));
 sky130_fd_sc_hd__mux2_1 _17644_ (.A0(_09955_),
    .A1(net147),
    .S(_09958_),
    .X(_09959_));
 sky130_fd_sc_hd__clkbuf_1 _17645_ (.A(_09959_),
    .X(_00562_));
 sky130_fd_sc_hd__nand2_1 _17646_ (.A(\wfg_drive_pat_top.patsel1_high_q[10] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[10].drv.axis_data_ff ),
    .Y(_09960_));
 sky130_fd_sc_hd__a211o_1 _17647_ (.A1(\wfg_drive_pat_top.patsel0_low_q[10] ),
    .A2(_09960_),
    .B1(_09952_),
    .C1(_09953_),
    .X(_09961_));
 sky130_fd_sc_hd__o211a_1 _17648_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[10].drv.axis_data_ff ),
    .A2(_09950_),
    .B1(_09961_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[10].drv.ctrl_en_q_i ),
    .X(_09962_));
 sky130_fd_sc_hd__and3b_1 _17649_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[10] ),
    .B(_09922_),
    .C(\wfg_drive_pat_top.patsel1_high_q[10] ),
    .X(_09963_));
 sky130_fd_sc_hd__o21a_1 _17650_ (.A1(_09956_),
    .A2(_09963_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[10].drv.ctrl_en_q_i ),
    .X(_09964_));
 sky130_fd_sc_hd__mux2_1 _17651_ (.A0(_09962_),
    .A1(net146),
    .S(_09964_),
    .X(_09965_));
 sky130_fd_sc_hd__clkbuf_1 _17652_ (.A(_09965_),
    .X(_00561_));
 sky130_fd_sc_hd__nand2_1 _17653_ (.A(\wfg_drive_pat_top.patsel1_high_q[0] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[0].drv.axis_data_ff ),
    .Y(_09966_));
 sky130_fd_sc_hd__a211o_1 _17654_ (.A1(\wfg_drive_pat_top.patsel0_low_q[0] ),
    .A2(_09966_),
    .B1(_09952_),
    .C1(_09953_),
    .X(_09967_));
 sky130_fd_sc_hd__o211a_1 _17655_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[0].drv.axis_data_ff ),
    .A2(_09950_),
    .B1(_09967_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[0].drv.ctrl_en_q_i ),
    .X(_09968_));
 sky130_fd_sc_hd__and3b_1 _17656_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[0] ),
    .B(_09922_),
    .C(\wfg_drive_pat_top.patsel1_high_q[0] ),
    .X(_09969_));
 sky130_fd_sc_hd__o21a_1 _17657_ (.A1(_09956_),
    .A2(_09969_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[0].drv.ctrl_en_q_i ),
    .X(_09970_));
 sky130_fd_sc_hd__mux2_1 _17658_ (.A0(_09968_),
    .A1(net145),
    .S(_09970_),
    .X(_09971_));
 sky130_fd_sc_hd__clkbuf_1 _17659_ (.A(_09971_),
    .X(_00560_));
 sky130_fd_sc_hd__nand2_1 _17660_ (.A(\wfg_drive_pat_top.patsel1_high_q[8] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[8].drv.axis_data_ff ),
    .Y(_09972_));
 sky130_fd_sc_hd__a211o_1 _17661_ (.A1(\wfg_drive_pat_top.patsel0_low_q[8] ),
    .A2(_09972_),
    .B1(_09952_),
    .C1(_09953_),
    .X(_09973_));
 sky130_fd_sc_hd__o211a_1 _17662_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[8].drv.axis_data_ff ),
    .A2(_09950_),
    .B1(_09973_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[8].drv.ctrl_en_q_i ),
    .X(_09974_));
 sky130_fd_sc_hd__and3b_1 _17663_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[8] ),
    .B(_09922_),
    .C(\wfg_drive_pat_top.patsel1_high_q[8] ),
    .X(_09975_));
 sky130_fd_sc_hd__o21a_1 _17664_ (.A1(_09956_),
    .A2(_09975_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[8].drv.ctrl_en_q_i ),
    .X(_09976_));
 sky130_fd_sc_hd__mux2_1 _17665_ (.A0(_09974_),
    .A1(net175),
    .S(_09976_),
    .X(_09977_));
 sky130_fd_sc_hd__clkbuf_1 _17666_ (.A(_09977_),
    .X(_00559_));
 sky130_fd_sc_hd__nand2_1 _17667_ (.A(\wfg_drive_pat_top.patsel1_high_q[7] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[7].drv.axis_data_ff ),
    .Y(_09978_));
 sky130_fd_sc_hd__a211o_1 _17668_ (.A1(\wfg_drive_pat_top.patsel0_low_q[7] ),
    .A2(_09978_),
    .B1(_09952_),
    .C1(_09953_),
    .X(_09979_));
 sky130_fd_sc_hd__o211a_1 _17669_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[7].drv.axis_data_ff ),
    .A2(_09950_),
    .B1(_09979_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[7].drv.ctrl_en_q_i ),
    .X(_09980_));
 sky130_fd_sc_hd__and3b_1 _17670_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[7] ),
    .B(_09922_),
    .C(\wfg_drive_pat_top.patsel1_high_q[7] ),
    .X(_09981_));
 sky130_fd_sc_hd__o21a_1 _17671_ (.A1(_09956_),
    .A2(_09981_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[7].drv.ctrl_en_q_i ),
    .X(_09982_));
 sky130_fd_sc_hd__mux2_1 _17672_ (.A0(_09980_),
    .A1(net174),
    .S(_09982_),
    .X(_09983_));
 sky130_fd_sc_hd__clkbuf_1 _17673_ (.A(_09983_),
    .X(_00558_));
 sky130_fd_sc_hd__nand2_1 _17674_ (.A(\wfg_drive_pat_top.patsel1_high_q[6] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[6].drv.axis_data_ff ),
    .Y(_09984_));
 sky130_fd_sc_hd__a211o_1 _17675_ (.A1(\wfg_drive_pat_top.patsel0_low_q[6] ),
    .A2(_09984_),
    .B1(_09952_),
    .C1(_09953_),
    .X(_09985_));
 sky130_fd_sc_hd__o211a_1 _17676_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[6].drv.axis_data_ff ),
    .A2(_09950_),
    .B1(_09985_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[6].drv.ctrl_en_q_i ),
    .X(_09986_));
 sky130_fd_sc_hd__and3b_1 _17677_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[6] ),
    .B(_09803_),
    .C(\wfg_drive_pat_top.patsel1_high_q[6] ),
    .X(_09987_));
 sky130_fd_sc_hd__o21a_1 _17678_ (.A1(_09956_),
    .A2(_09987_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[6].drv.ctrl_en_q_i ),
    .X(_09988_));
 sky130_fd_sc_hd__mux2_1 _17679_ (.A0(_09986_),
    .A1(net173),
    .S(_09988_),
    .X(_09989_));
 sky130_fd_sc_hd__clkbuf_1 _17680_ (.A(_09989_),
    .X(_00557_));
 sky130_fd_sc_hd__nand2_1 _17681_ (.A(\wfg_drive_pat_top.patsel1_high_q[5] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[5].drv.axis_data_ff ),
    .Y(_09990_));
 sky130_fd_sc_hd__a211o_1 _17682_ (.A1(\wfg_drive_pat_top.patsel0_low_q[5] ),
    .A2(_09990_),
    .B1(_09952_),
    .C1(_09953_),
    .X(_09991_));
 sky130_fd_sc_hd__o211a_1 _17683_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[5].drv.axis_data_ff ),
    .A2(_09950_),
    .B1(_09991_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[5].drv.ctrl_en_q_i ),
    .X(_09992_));
 sky130_fd_sc_hd__and3b_1 _17684_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[5] ),
    .B(_09803_),
    .C(\wfg_drive_pat_top.patsel1_high_q[5] ),
    .X(_09993_));
 sky130_fd_sc_hd__o21a_1 _17685_ (.A1(_09956_),
    .A2(_09993_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[5].drv.ctrl_en_q_i ),
    .X(_09994_));
 sky130_fd_sc_hd__mux2_1 _17686_ (.A0(_09992_),
    .A1(net172),
    .S(_09994_),
    .X(_09995_));
 sky130_fd_sc_hd__clkbuf_1 _17687_ (.A(_09995_),
    .X(_00556_));
 sky130_fd_sc_hd__nand2_1 _17688_ (.A(\wfg_drive_pat_top.patsel1_high_q[4] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[4].drv.axis_data_ff ),
    .Y(_09996_));
 sky130_fd_sc_hd__a211o_1 _17689_ (.A1(\wfg_drive_pat_top.patsel0_low_q[4] ),
    .A2(_09996_),
    .B1(_09952_),
    .C1(_09953_),
    .X(_09997_));
 sky130_fd_sc_hd__o211a_1 _17690_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[4].drv.axis_data_ff ),
    .A2(_09950_),
    .B1(_09997_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[4].drv.ctrl_en_q_i ),
    .X(_09998_));
 sky130_fd_sc_hd__and3b_1 _17691_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[4] ),
    .B(_09803_),
    .C(\wfg_drive_pat_top.patsel1_high_q[4] ),
    .X(_09999_));
 sky130_fd_sc_hd__o21a_1 _17692_ (.A1(_09956_),
    .A2(_09999_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[4].drv.ctrl_en_q_i ),
    .X(_10000_));
 sky130_fd_sc_hd__mux2_1 _17693_ (.A0(_09998_),
    .A1(net171),
    .S(_10000_),
    .X(_10001_));
 sky130_fd_sc_hd__clkbuf_1 _17694_ (.A(_10001_),
    .X(_00555_));
 sky130_fd_sc_hd__nand2_1 _17695_ (.A(\wfg_drive_pat_top.patsel1_high_q[3] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[3].drv.axis_data_ff ),
    .Y(_10002_));
 sky130_fd_sc_hd__a211o_1 _17696_ (.A1(\wfg_drive_pat_top.patsel0_low_q[3] ),
    .A2(_10002_),
    .B1(_09952_),
    .C1(_09953_),
    .X(_10003_));
 sky130_fd_sc_hd__o211a_1 _17697_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[3].drv.axis_data_ff ),
    .A2(_09950_),
    .B1(_10003_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[3].drv.ctrl_en_q_i ),
    .X(_10004_));
 sky130_fd_sc_hd__and3b_1 _17698_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[3] ),
    .B(_09803_),
    .C(\wfg_drive_pat_top.patsel1_high_q[3] ),
    .X(_10005_));
 sky130_fd_sc_hd__o21a_1 _17699_ (.A1(_09956_),
    .A2(_10005_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[3].drv.ctrl_en_q_i ),
    .X(_10006_));
 sky130_fd_sc_hd__mux2_1 _17700_ (.A0(_10004_),
    .A1(net170),
    .S(_10006_),
    .X(_10007_));
 sky130_fd_sc_hd__clkbuf_1 _17701_ (.A(_10007_),
    .X(_00554_));
 sky130_fd_sc_hd__nand2_1 _17702_ (.A(\wfg_drive_pat_top.patsel1_high_q[31] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[31].drv.axis_data_ff ),
    .Y(_10008_));
 sky130_fd_sc_hd__a211o_1 _17703_ (.A1(\wfg_drive_pat_top.patsel0_low_q[31] ),
    .A2(_10008_),
    .B1(_09952_),
    .C1(_09953_),
    .X(_10009_));
 sky130_fd_sc_hd__o211a_1 _17704_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[31].drv.axis_data_ff ),
    .A2(_09950_),
    .B1(_10009_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[31].drv.ctrl_en_q_i ),
    .X(_10010_));
 sky130_fd_sc_hd__and3b_1 _17705_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[31] ),
    .B(_09803_),
    .C(\wfg_drive_pat_top.patsel1_high_q[31] ),
    .X(_10011_));
 sky130_fd_sc_hd__o21a_1 _17706_ (.A1(_09956_),
    .A2(_10011_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[31].drv.ctrl_en_q_i ),
    .X(_10012_));
 sky130_fd_sc_hd__mux2_1 _17707_ (.A0(_10010_),
    .A1(net169),
    .S(_10012_),
    .X(_10013_));
 sky130_fd_sc_hd__clkbuf_1 _17708_ (.A(_10013_),
    .X(_00553_));
 sky130_fd_sc_hd__nand2_1 _17709_ (.A(\wfg_drive_pat_top.patsel1_high_q[29] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[29].drv.axis_data_ff ),
    .Y(_10014_));
 sky130_fd_sc_hd__a211o_1 _17710_ (.A1(\wfg_drive_pat_top.patsel0_low_q[29] ),
    .A2(_10014_),
    .B1(_09801_),
    .C1(_09791_),
    .X(_10015_));
 sky130_fd_sc_hd__o211a_1 _17711_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[29].drv.axis_data_ff ),
    .A2(_09804_),
    .B1(_10015_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[29].drv.ctrl_en_q_i ),
    .X(_10016_));
 sky130_fd_sc_hd__and3b_1 _17712_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[29] ),
    .B(_09803_),
    .C(\wfg_drive_pat_top.patsel1_high_q[29] ),
    .X(_10017_));
 sky130_fd_sc_hd__o21a_1 _17713_ (.A1(_09825_),
    .A2(_10017_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[29].drv.ctrl_en_q_i ),
    .X(_10018_));
 sky130_fd_sc_hd__mux2_1 _17714_ (.A0(_10016_),
    .A1(net166),
    .S(_10018_),
    .X(_10019_));
 sky130_fd_sc_hd__clkbuf_1 _17715_ (.A(_10019_),
    .X(_00552_));
 sky130_fd_sc_hd__nand2_1 _17716_ (.A(\wfg_drive_pat_top.patsel1_high_q[19] ),
    .B(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[19].drv.axis_data_ff ),
    .Y(_10020_));
 sky130_fd_sc_hd__a211o_1 _17717_ (.A1(\wfg_drive_pat_top.patsel0_low_q[19] ),
    .A2(_10020_),
    .B1(_09801_),
    .C1(_09791_),
    .X(_10021_));
 sky130_fd_sc_hd__o211a_1 _17718_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[19].drv.axis_data_ff ),
    .A2(_09804_),
    .B1(_10021_),
    .C1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[19].drv.ctrl_en_q_i ),
    .X(_10022_));
 sky130_fd_sc_hd__and3b_1 _17719_ (.A_N(\wfg_drive_pat_top.patsel0_low_q[19] ),
    .B(_09803_),
    .C(\wfg_drive_pat_top.patsel1_high_q[19] ),
    .X(_10023_));
 sky130_fd_sc_hd__o21a_1 _17720_ (.A1(_09825_),
    .A2(_10023_),
    .B1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[19].drv.ctrl_en_q_i ),
    .X(_10024_));
 sky130_fd_sc_hd__mux2_1 _17721_ (.A0(_10022_),
    .A1(net155),
    .S(_10024_),
    .X(_10025_));
 sky130_fd_sc_hd__clkbuf_1 _17722_ (.A(_10025_),
    .X(_00551_));
 sky130_fd_sc_hd__buf_2 _17723_ (.A(_06357_),
    .X(_10026_));
 sky130_fd_sc_hd__buf_4 _17724_ (.A(_06358_),
    .X(_10027_));
 sky130_fd_sc_hd__and2_2 _17725_ (.A(\wfg_interconnect_top.stimulus_0[17] ),
    .B(_10027_),
    .X(_10028_));
 sky130_fd_sc_hd__buf_2 _17726_ (.A(_10028_),
    .X(_10029_));
 sky130_fd_sc_hd__a21o_1 _17727_ (.A1(\wfg_interconnect_top.stimulus_1[31] ),
    .A2(_10026_),
    .B1(_10029_),
    .X(_10030_));
 sky130_fd_sc_hd__a22o_1 _17728_ (.A1(\wfg_interconnect_top.stimulus_1[32] ),
    .A2(_05977_),
    .B1(_10027_),
    .B2(\wfg_interconnect_top.stimulus_0[32] ),
    .X(_10031_));
 sky130_fd_sc_hd__mux2_1 _17729_ (.A0(_02708_),
    .A1(_02709_),
    .S(_09782_),
    .X(_10032_));
 sky130_fd_sc_hd__clkbuf_1 _17730_ (.A(_10032_),
    .X(\wfg_drive_pat_top.wfg_drive_pat.wfg_sync_i ));
 sky130_fd_sc_hd__and2_4 _17731_ (.A(_10031_),
    .B(\wfg_drive_pat_top.wfg_drive_pat.wfg_sync_i ),
    .X(_10033_));
 sky130_fd_sc_hd__clkbuf_4 _17732_ (.A(_10033_),
    .X(_10034_));
 sky130_fd_sc_hd__mux2_1 _17733_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[31].drv.axis_data_ff ),
    .A1(_10030_),
    .S(_10034_),
    .X(_10035_));
 sky130_fd_sc_hd__clkbuf_1 _17734_ (.A(_10035_),
    .X(_00550_));
 sky130_fd_sc_hd__a21o_1 _17735_ (.A1(\wfg_interconnect_top.stimulus_1[30] ),
    .A2(_10026_),
    .B1(_10029_),
    .X(_10036_));
 sky130_fd_sc_hd__mux2_1 _17736_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[30].drv.axis_data_ff ),
    .A1(_10036_),
    .S(_10034_),
    .X(_10037_));
 sky130_fd_sc_hd__clkbuf_1 _17737_ (.A(_10037_),
    .X(_00549_));
 sky130_fd_sc_hd__a21o_1 _17738_ (.A1(\wfg_interconnect_top.stimulus_1[29] ),
    .A2(_10026_),
    .B1(_10029_),
    .X(_10038_));
 sky130_fd_sc_hd__mux2_1 _17739_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[29].drv.axis_data_ff ),
    .A1(_10038_),
    .S(_10034_),
    .X(_10039_));
 sky130_fd_sc_hd__clkbuf_1 _17740_ (.A(_10039_),
    .X(_00548_));
 sky130_fd_sc_hd__a21o_1 _17741_ (.A1(\wfg_interconnect_top.stimulus_1[28] ),
    .A2(_10026_),
    .B1(_10029_),
    .X(_10040_));
 sky130_fd_sc_hd__mux2_1 _17742_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[28].drv.axis_data_ff ),
    .A1(_10040_),
    .S(_10034_),
    .X(_10041_));
 sky130_fd_sc_hd__clkbuf_1 _17743_ (.A(_10041_),
    .X(_00547_));
 sky130_fd_sc_hd__a21o_1 _17744_ (.A1(\wfg_interconnect_top.stimulus_1[27] ),
    .A2(_10026_),
    .B1(_10029_),
    .X(_10042_));
 sky130_fd_sc_hd__mux2_1 _17745_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[27].drv.axis_data_ff ),
    .A1(_10042_),
    .S(_10034_),
    .X(_10043_));
 sky130_fd_sc_hd__clkbuf_1 _17746_ (.A(_10043_),
    .X(_00546_));
 sky130_fd_sc_hd__a21o_1 _17747_ (.A1(\wfg_interconnect_top.stimulus_1[26] ),
    .A2(_10026_),
    .B1(_10029_),
    .X(_10044_));
 sky130_fd_sc_hd__mux2_1 _17748_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[26].drv.axis_data_ff ),
    .A1(_10044_),
    .S(_10034_),
    .X(_10045_));
 sky130_fd_sc_hd__clkbuf_1 _17749_ (.A(_10045_),
    .X(_00545_));
 sky130_fd_sc_hd__a21o_1 _17750_ (.A1(\wfg_interconnect_top.stimulus_1[25] ),
    .A2(_10026_),
    .B1(_10029_),
    .X(_10046_));
 sky130_fd_sc_hd__mux2_1 _17751_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[25].drv.axis_data_ff ),
    .A1(_10046_),
    .S(_10034_),
    .X(_10047_));
 sky130_fd_sc_hd__clkbuf_1 _17752_ (.A(_10047_),
    .X(_00544_));
 sky130_fd_sc_hd__a21o_1 _17753_ (.A1(\wfg_interconnect_top.stimulus_1[24] ),
    .A2(_10026_),
    .B1(_10029_),
    .X(_10048_));
 sky130_fd_sc_hd__mux2_1 _17754_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[24].drv.axis_data_ff ),
    .A1(_10048_),
    .S(_10034_),
    .X(_10049_));
 sky130_fd_sc_hd__clkbuf_1 _17755_ (.A(_10049_),
    .X(_00543_));
 sky130_fd_sc_hd__a21o_1 _17756_ (.A1(\wfg_interconnect_top.stimulus_1[23] ),
    .A2(_10026_),
    .B1(_10029_),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _17757_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[23].drv.axis_data_ff ),
    .A1(_01293_),
    .S(_10034_),
    .X(_01294_));
 sky130_fd_sc_hd__clkbuf_1 _17758_ (.A(_01294_),
    .X(_00542_));
 sky130_fd_sc_hd__a21o_1 _17759_ (.A1(\wfg_interconnect_top.stimulus_1[22] ),
    .A2(_10026_),
    .B1(_10029_),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _17760_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[22].drv.axis_data_ff ),
    .A1(_01295_),
    .S(_10034_),
    .X(_01296_));
 sky130_fd_sc_hd__clkbuf_1 _17761_ (.A(_01296_),
    .X(_00541_));
 sky130_fd_sc_hd__a21o_1 _17762_ (.A1(\wfg_interconnect_top.stimulus_1[21] ),
    .A2(_06357_),
    .B1(_10028_),
    .X(_01297_));
 sky130_fd_sc_hd__clkbuf_4 _17763_ (.A(_10033_),
    .X(_01298_));
 sky130_fd_sc_hd__mux2_1 _17764_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[21].drv.axis_data_ff ),
    .A1(_01297_),
    .S(_01298_),
    .X(_01299_));
 sky130_fd_sc_hd__clkbuf_1 _17765_ (.A(_01299_),
    .X(_00540_));
 sky130_fd_sc_hd__a21o_1 _17766_ (.A1(\wfg_interconnect_top.stimulus_1[20] ),
    .A2(_06357_),
    .B1(_10028_),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_1 _17767_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[20].drv.axis_data_ff ),
    .A1(_01300_),
    .S(_01298_),
    .X(_01301_));
 sky130_fd_sc_hd__clkbuf_1 _17768_ (.A(_01301_),
    .X(_00539_));
 sky130_fd_sc_hd__a21o_1 _17769_ (.A1(\wfg_interconnect_top.stimulus_1[19] ),
    .A2(_06357_),
    .B1(_10028_),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _17770_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[19].drv.axis_data_ff ),
    .A1(_01302_),
    .S(_01298_),
    .X(_01303_));
 sky130_fd_sc_hd__clkbuf_1 _17771_ (.A(_01303_),
    .X(_00538_));
 sky130_fd_sc_hd__a21o_1 _17772_ (.A1(\wfg_interconnect_top.stimulus_1[18] ),
    .A2(_06357_),
    .B1(_10028_),
    .X(_01304_));
 sky130_fd_sc_hd__mux2_1 _17773_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[18].drv.axis_data_ff ),
    .A1(_01304_),
    .S(_01298_),
    .X(_01305_));
 sky130_fd_sc_hd__clkbuf_1 _17774_ (.A(_01305_),
    .X(_00537_));
 sky130_fd_sc_hd__a21o_1 _17775_ (.A1(\wfg_interconnect_top.stimulus_1[17] ),
    .A2(_06357_),
    .B1(_10028_),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _17776_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[17].drv.axis_data_ff ),
    .A1(_01306_),
    .S(_01298_),
    .X(_01307_));
 sky130_fd_sc_hd__clkbuf_1 _17777_ (.A(_01307_),
    .X(_00536_));
 sky130_fd_sc_hd__clkbuf_4 _17778_ (.A(_10027_),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _17779_ (.A0(\wfg_interconnect_top.stimulus_1[16] ),
    .A1(\wfg_interconnect_top.stimulus_0[16] ),
    .S(_01308_),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _17780_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[16].drv.axis_data_ff ),
    .A1(_01309_),
    .S(_01298_),
    .X(_01310_));
 sky130_fd_sc_hd__clkbuf_1 _17781_ (.A(_01310_),
    .X(_00535_));
 sky130_fd_sc_hd__mux2_1 _17782_ (.A0(\wfg_interconnect_top.stimulus_1[15] ),
    .A1(\wfg_interconnect_top.stimulus_0[15] ),
    .S(_01308_),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _17783_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[15].drv.axis_data_ff ),
    .A1(_01311_),
    .S(_01298_),
    .X(_01312_));
 sky130_fd_sc_hd__clkbuf_1 _17784_ (.A(_01312_),
    .X(_00534_));
 sky130_fd_sc_hd__mux2_1 _17785_ (.A0(\wfg_interconnect_top.stimulus_1[14] ),
    .A1(\wfg_interconnect_top.stimulus_0[14] ),
    .S(_01308_),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _17786_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[14].drv.axis_data_ff ),
    .A1(_01313_),
    .S(_01298_),
    .X(_01314_));
 sky130_fd_sc_hd__clkbuf_1 _17787_ (.A(_01314_),
    .X(_00533_));
 sky130_fd_sc_hd__mux2_1 _17788_ (.A0(\wfg_interconnect_top.stimulus_1[13] ),
    .A1(\wfg_interconnect_top.stimulus_0[13] ),
    .S(_01308_),
    .X(_01315_));
 sky130_fd_sc_hd__mux2_1 _17789_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[13].drv.axis_data_ff ),
    .A1(_01315_),
    .S(_01298_),
    .X(_01316_));
 sky130_fd_sc_hd__clkbuf_1 _17790_ (.A(_01316_),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_1 _17791_ (.A0(\wfg_interconnect_top.stimulus_1[12] ),
    .A1(\wfg_interconnect_top.stimulus_0[12] ),
    .S(_01308_),
    .X(_01317_));
 sky130_fd_sc_hd__mux2_1 _17792_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[12].drv.axis_data_ff ),
    .A1(_01317_),
    .S(_01298_),
    .X(_01318_));
 sky130_fd_sc_hd__clkbuf_1 _17793_ (.A(_01318_),
    .X(_00531_));
 sky130_fd_sc_hd__mux2_1 _17794_ (.A0(\wfg_interconnect_top.stimulus_1[11] ),
    .A1(\wfg_interconnect_top.stimulus_0[11] ),
    .S(_01308_),
    .X(_01319_));
 sky130_fd_sc_hd__clkbuf_4 _17795_ (.A(_10033_),
    .X(_01320_));
 sky130_fd_sc_hd__mux2_1 _17796_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[11].drv.axis_data_ff ),
    .A1(_01319_),
    .S(_01320_),
    .X(_01321_));
 sky130_fd_sc_hd__clkbuf_1 _17797_ (.A(_01321_),
    .X(_00530_));
 sky130_fd_sc_hd__mux2_1 _17798_ (.A0(\wfg_interconnect_top.stimulus_1[10] ),
    .A1(\wfg_interconnect_top.stimulus_0[10] ),
    .S(_01308_),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_1 _17799_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[10].drv.axis_data_ff ),
    .A1(_01322_),
    .S(_01320_),
    .X(_01323_));
 sky130_fd_sc_hd__clkbuf_1 _17800_ (.A(_01323_),
    .X(_00529_));
 sky130_fd_sc_hd__mux2_1 _17801_ (.A0(\wfg_interconnect_top.stimulus_1[9] ),
    .A1(\wfg_interconnect_top.stimulus_0[9] ),
    .S(_01308_),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_1 _17802_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[9].drv.axis_data_ff ),
    .A1(_01324_),
    .S(_01320_),
    .X(_01325_));
 sky130_fd_sc_hd__clkbuf_1 _17803_ (.A(_01325_),
    .X(_00528_));
 sky130_fd_sc_hd__mux2_1 _17804_ (.A0(\wfg_interconnect_top.stimulus_1[8] ),
    .A1(\wfg_interconnect_top.stimulus_0[8] ),
    .S(_01308_),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_1 _17805_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[8].drv.axis_data_ff ),
    .A1(_01326_),
    .S(_01320_),
    .X(_01327_));
 sky130_fd_sc_hd__clkbuf_1 _17806_ (.A(_01327_),
    .X(_00527_));
 sky130_fd_sc_hd__mux2_1 _17807_ (.A0(\wfg_interconnect_top.stimulus_1[7] ),
    .A1(\wfg_interconnect_top.stimulus_0[7] ),
    .S(_01308_),
    .X(_01328_));
 sky130_fd_sc_hd__mux2_1 _17808_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[7].drv.axis_data_ff ),
    .A1(_01328_),
    .S(_01320_),
    .X(_01329_));
 sky130_fd_sc_hd__clkbuf_1 _17809_ (.A(_01329_),
    .X(_00526_));
 sky130_fd_sc_hd__mux2_1 _17810_ (.A0(\wfg_interconnect_top.stimulus_1[6] ),
    .A1(\wfg_interconnect_top.stimulus_0[6] ),
    .S(_10027_),
    .X(_01330_));
 sky130_fd_sc_hd__mux2_1 _17811_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[6].drv.axis_data_ff ),
    .A1(_01330_),
    .S(_01320_),
    .X(_01331_));
 sky130_fd_sc_hd__clkbuf_1 _17812_ (.A(_01331_),
    .X(_00525_));
 sky130_fd_sc_hd__mux2_1 _17813_ (.A0(\wfg_interconnect_top.stimulus_1[5] ),
    .A1(\wfg_interconnect_top.stimulus_0[5] ),
    .S(_10027_),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_1 _17814_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[5].drv.axis_data_ff ),
    .A1(_01332_),
    .S(_01320_),
    .X(_01333_));
 sky130_fd_sc_hd__clkbuf_1 _17815_ (.A(_01333_),
    .X(_00524_));
 sky130_fd_sc_hd__mux2_1 _17816_ (.A0(\wfg_interconnect_top.stimulus_1[4] ),
    .A1(\wfg_interconnect_top.stimulus_0[4] ),
    .S(_10027_),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _17817_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[4].drv.axis_data_ff ),
    .A1(_01334_),
    .S(_01320_),
    .X(_01335_));
 sky130_fd_sc_hd__clkbuf_1 _17818_ (.A(_01335_),
    .X(_00523_));
 sky130_fd_sc_hd__mux2_1 _17819_ (.A0(\wfg_interconnect_top.stimulus_1[3] ),
    .A1(\wfg_interconnect_top.stimulus_0[3] ),
    .S(_10027_),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _17820_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[3].drv.axis_data_ff ),
    .A1(_01336_),
    .S(_01320_),
    .X(_01337_));
 sky130_fd_sc_hd__clkbuf_1 _17821_ (.A(_01337_),
    .X(_00522_));
 sky130_fd_sc_hd__mux2_1 _17822_ (.A0(\wfg_interconnect_top.stimulus_1[2] ),
    .A1(\wfg_interconnect_top.stimulus_0[2] ),
    .S(_10027_),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _17823_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[2].drv.axis_data_ff ),
    .A1(_01338_),
    .S(_01320_),
    .X(_01339_));
 sky130_fd_sc_hd__clkbuf_1 _17824_ (.A(_01339_),
    .X(_00521_));
 sky130_fd_sc_hd__mux2_1 _17825_ (.A0(\wfg_interconnect_top.stimulus_1[1] ),
    .A1(\wfg_interconnect_top.stimulus_0[1] ),
    .S(_10027_),
    .X(_01340_));
 sky130_fd_sc_hd__mux2_1 _17826_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[1].drv.axis_data_ff ),
    .A1(_01340_),
    .S(_10033_),
    .X(_01341_));
 sky130_fd_sc_hd__clkbuf_1 _17827_ (.A(_01341_),
    .X(_00520_));
 sky130_fd_sc_hd__mux2_1 _17828_ (.A0(\wfg_interconnect_top.stimulus_1[0] ),
    .A1(\wfg_interconnect_top.stimulus_0[0] ),
    .S(_10027_),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _17829_ (.A0(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[0].drv.axis_data_ff ),
    .A1(_01342_),
    .S(_10033_),
    .X(_01343_));
 sky130_fd_sc_hd__clkbuf_1 _17830_ (.A(_01343_),
    .X(_00519_));
 sky130_fd_sc_hd__and3_1 _17831_ (.A(\wfg_core_top.wfg_core.subcycle_pls_cnt[2] ),
    .B(\wfg_core_top.wfg_core.subcycle_pls_cnt[1] ),
    .C(\wfg_core_top.wfg_core.subcycle_pls_cnt[0] ),
    .X(_01344_));
 sky130_fd_sc_hd__and3_1 _17832_ (.A(\wfg_core_top.wfg_core.subcycle_pls_cnt[4] ),
    .B(\wfg_core_top.wfg_core.subcycle_pls_cnt[3] ),
    .C(_01344_),
    .X(_01345_));
 sky130_fd_sc_hd__and2_1 _17833_ (.A(\wfg_core_top.wfg_core.subcycle_pls_cnt[5] ),
    .B(_01345_),
    .X(_01346_));
 sky130_fd_sc_hd__and2b_1 _17834_ (.A_N(\wfg_core_top.wfg_core.subcycle_dly ),
    .B(\wfg_core_top.wfg_core.temp_subcycle ),
    .X(_01347_));
 sky130_fd_sc_hd__clkbuf_2 _17835_ (.A(_01347_),
    .X(_01348_));
 sky130_fd_sc_hd__and3b_1 _17836_ (.A_N(_02708_),
    .B(_01348_),
    .C(\wfg_core_top.active_o ),
    .X(_01349_));
 sky130_fd_sc_hd__and3_1 _17837_ (.A(\wfg_core_top.wfg_core.subcycle_pls_cnt[6] ),
    .B(_01346_),
    .C(_01349_),
    .X(_01350_));
 sky130_fd_sc_hd__inv_4 _17838_ (.A(\wfg_core_top.active_o ),
    .Y(_01351_));
 sky130_fd_sc_hd__or2_1 _17839_ (.A(_01351_),
    .B(_02708_),
    .X(_01352_));
 sky130_fd_sc_hd__a31oi_1 _17840_ (.A1(\wfg_core_top.wfg_core.subcycle_pls_cnt[6] ),
    .A2(_01346_),
    .A3(_01348_),
    .B1(_01352_),
    .Y(_01353_));
 sky130_fd_sc_hd__mux2_1 _17841_ (.A0(_01350_),
    .A1(_01353_),
    .S(\wfg_core_top.wfg_core.subcycle_pls_cnt[7] ),
    .X(_01354_));
 sky130_fd_sc_hd__clkbuf_1 _17842_ (.A(_01354_),
    .X(_00491_));
 sky130_fd_sc_hd__a31o_1 _17843_ (.A1(\wfg_core_top.wfg_core.subcycle_pls_cnt[5] ),
    .A2(_01345_),
    .A3(_01349_),
    .B1(\wfg_core_top.wfg_core.subcycle_pls_cnt[6] ),
    .X(_01355_));
 sky130_fd_sc_hd__and2_1 _17844_ (.A(_01353_),
    .B(_01355_),
    .X(_01356_));
 sky130_fd_sc_hd__clkbuf_1 _17845_ (.A(_01356_),
    .X(_00490_));
 sky130_fd_sc_hd__o21ai_1 _17846_ (.A1(\wfg_core_top.wfg_core.subcycle_pls_cnt[5] ),
    .A2(_01345_),
    .B1(_01349_),
    .Y(_01357_));
 sky130_fd_sc_hd__nor2_1 _17847_ (.A(_01348_),
    .B(_01352_),
    .Y(_01358_));
 sky130_fd_sc_hd__a2bb2o_1 _17848_ (.A1_N(_01346_),
    .A2_N(_01357_),
    .B1(_01358_),
    .B2(\wfg_core_top.wfg_core.subcycle_pls_cnt[5] ),
    .X(_00489_));
 sky130_fd_sc_hd__inv_2 _17849_ (.A(_01345_),
    .Y(_01359_));
 sky130_fd_sc_hd__a21o_1 _17850_ (.A1(\wfg_core_top.wfg_core.subcycle_pls_cnt[3] ),
    .A2(_01344_),
    .B1(\wfg_core_top.wfg_core.subcycle_pls_cnt[4] ),
    .X(_01360_));
 sky130_fd_sc_hd__a32o_1 _17851_ (.A1(_01359_),
    .A2(_01349_),
    .A3(_01360_),
    .B1(_01358_),
    .B2(\wfg_core_top.wfg_core.subcycle_pls_cnt[4] ),
    .X(_00488_));
 sky130_fd_sc_hd__a21oi_1 _17852_ (.A1(_01344_),
    .A2(_01348_),
    .B1(\wfg_core_top.wfg_core.subcycle_pls_cnt[3] ),
    .Y(_01361_));
 sky130_fd_sc_hd__a311oi_1 _17853_ (.A1(\wfg_core_top.wfg_core.subcycle_pls_cnt[3] ),
    .A2(_01344_),
    .A3(_01348_),
    .B1(_01352_),
    .C1(_01361_),
    .Y(_00487_));
 sky130_fd_sc_hd__inv_2 _17854_ (.A(_01344_),
    .Y(_01362_));
 sky130_fd_sc_hd__a21o_1 _17855_ (.A1(\wfg_core_top.wfg_core.subcycle_pls_cnt[1] ),
    .A2(\wfg_core_top.wfg_core.subcycle_pls_cnt[0] ),
    .B1(\wfg_core_top.wfg_core.subcycle_pls_cnt[2] ),
    .X(_01363_));
 sky130_fd_sc_hd__a32o_1 _17856_ (.A1(_01362_),
    .A2(_01349_),
    .A3(_01363_),
    .B1(_01358_),
    .B2(\wfg_core_top.wfg_core.subcycle_pls_cnt[2] ),
    .X(_00486_));
 sky130_fd_sc_hd__a21oi_1 _17857_ (.A1(\wfg_core_top.wfg_core.subcycle_pls_cnt[0] ),
    .A2(_01348_),
    .B1(\wfg_core_top.wfg_core.subcycle_pls_cnt[1] ),
    .Y(_01364_));
 sky130_fd_sc_hd__a31o_1 _17858_ (.A1(\wfg_core_top.wfg_core.subcycle_pls_cnt[1] ),
    .A2(\wfg_core_top.wfg_core.subcycle_pls_cnt[0] ),
    .A3(_01348_),
    .B1(_01352_),
    .X(_01365_));
 sky130_fd_sc_hd__nor2_1 _17859_ (.A(_01364_),
    .B(_01365_),
    .Y(_00485_));
 sky130_fd_sc_hd__mux2_1 _17860_ (.A0(_01349_),
    .A1(_01358_),
    .S(\wfg_core_top.wfg_core.subcycle_pls_cnt[0] ),
    .X(_01366_));
 sky130_fd_sc_hd__clkbuf_1 _17861_ (.A(_01366_),
    .X(_00484_));
 sky130_fd_sc_hd__or3_1 _17862_ (.A(\wfg_core_top.wfg_core.sync_count[2] ),
    .B(\wfg_core_top.wfg_core.sync_count[1] ),
    .C(\wfg_core_top.wfg_core.sync_count[0] ),
    .X(_01367_));
 sky130_fd_sc_hd__or2_1 _17863_ (.A(\wfg_core_top.wfg_core.sync_count[3] ),
    .B(_01367_),
    .X(_01368_));
 sky130_fd_sc_hd__or3_1 _17864_ (.A(\wfg_core_top.wfg_core.sync_count[5] ),
    .B(\wfg_core_top.wfg_core.sync_count[4] ),
    .C(_01368_),
    .X(_01369_));
 sky130_fd_sc_hd__or2_1 _17865_ (.A(\wfg_core_top.wfg_core.sync_count[6] ),
    .B(_01369_),
    .X(_01370_));
 sky130_fd_sc_hd__or2_1 _17866_ (.A(\wfg_core_top.wfg_core.sync_count[7] ),
    .B(_01370_),
    .X(_01371_));
 sky130_fd_sc_hd__buf_2 _17867_ (.A(_01371_),
    .X(_01372_));
 sky130_fd_sc_hd__or3_1 _17868_ (.A(\wfg_core_top.wfg_core.subcycle_count[2] ),
    .B(\wfg_core_top.wfg_core.subcycle_count[1] ),
    .C(\wfg_core_top.wfg_core.subcycle_count[0] ),
    .X(_01373_));
 sky130_fd_sc_hd__or2_1 _17869_ (.A(\wfg_core_top.wfg_core.subcycle_count[3] ),
    .B(_01373_),
    .X(_01374_));
 sky130_fd_sc_hd__or3_1 _17870_ (.A(\wfg_core_top.wfg_core.subcycle_count[5] ),
    .B(\wfg_core_top.wfg_core.subcycle_count[4] ),
    .C(_01374_),
    .X(_01375_));
 sky130_fd_sc_hd__or2_1 _17871_ (.A(\wfg_core_top.wfg_core.subcycle_count[6] ),
    .B(_01375_),
    .X(_01376_));
 sky130_fd_sc_hd__or3_1 _17872_ (.A(\wfg_core_top.wfg_core.subcycle_count[8] ),
    .B(\wfg_core_top.wfg_core.subcycle_count[7] ),
    .C(_01376_),
    .X(_01377_));
 sky130_fd_sc_hd__or2_2 _17873_ (.A(\wfg_core_top.wfg_core.subcycle_count[9] ),
    .B(_01377_),
    .X(_01378_));
 sky130_fd_sc_hd__or3_1 _17874_ (.A(\wfg_core_top.wfg_core.subcycle_count[11] ),
    .B(\wfg_core_top.wfg_core.subcycle_count[10] ),
    .C(_01378_),
    .X(_01379_));
 sky130_fd_sc_hd__or2_1 _17875_ (.A(\wfg_core_top.wfg_core.subcycle_count[12] ),
    .B(_01379_),
    .X(_01380_));
 sky130_fd_sc_hd__or2_1 _17876_ (.A(\wfg_core_top.wfg_core.subcycle_count[13] ),
    .B(_01380_),
    .X(_01381_));
 sky130_fd_sc_hd__or2_1 _17877_ (.A(\wfg_core_top.wfg_core.subcycle_count[14] ),
    .B(_01381_),
    .X(_01382_));
 sky130_fd_sc_hd__or2_1 _17878_ (.A(\wfg_core_top.wfg_core.subcycle_count[15] ),
    .B(_01382_),
    .X(_01383_));
 sky130_fd_sc_hd__clkbuf_4 _17879_ (.A(_01383_),
    .X(_01384_));
 sky130_fd_sc_hd__nor2_1 _17880_ (.A(_01372_),
    .B(_01384_),
    .Y(_01385_));
 sky130_fd_sc_hd__o21ai_1 _17881_ (.A1(\wfg_core_top.wfg_core.temp_sync ),
    .A2(_01385_),
    .B1(\wfg_core_top.active_o ),
    .Y(_01386_));
 sky130_fd_sc_hd__a21oi_1 _17882_ (.A1(\wfg_core_top.wfg_core.temp_sync ),
    .A2(_01385_),
    .B1(_01386_),
    .Y(_00481_));
 sky130_fd_sc_hd__nor2_4 _17883_ (.A(_01351_),
    .B(_01384_),
    .Y(_01387_));
 sky130_fd_sc_hd__and2_1 _17884_ (.A(\wfg_core_top.active_o ),
    .B(_01384_),
    .X(_01388_));
 sky130_fd_sc_hd__buf_2 _17885_ (.A(_01388_),
    .X(_01389_));
 sky130_fd_sc_hd__mux2_1 _17886_ (.A0(_01387_),
    .A1(_01389_),
    .S(\wfg_core_top.wfg_core.temp_subcycle ),
    .X(_01390_));
 sky130_fd_sc_hd__clkbuf_1 _17887_ (.A(_01390_),
    .X(_00480_));
 sky130_fd_sc_hd__inv_2 _17888_ (.A(\wfg_core_top.cfg_sync_q[7] ),
    .Y(_01391_));
 sky130_fd_sc_hd__nand2_1 _17889_ (.A(\wfg_core_top.wfg_core.sync_count[7] ),
    .B(_01370_),
    .Y(_01392_));
 sky130_fd_sc_hd__o21ai_1 _17890_ (.A1(_01391_),
    .A2(_01372_),
    .B1(_01392_),
    .Y(_01393_));
 sky130_fd_sc_hd__a22o_1 _17891_ (.A1(\wfg_core_top.wfg_core.sync_count[7] ),
    .A2(_01389_),
    .B1(_01387_),
    .B2(_01393_),
    .X(_00479_));
 sky130_fd_sc_hd__clkbuf_4 _17892_ (.A(_01384_),
    .X(_01394_));
 sky130_fd_sc_hd__and2_1 _17893_ (.A(\wfg_core_top.wfg_core.sync_count[6] ),
    .B(_01369_),
    .X(_01395_));
 sky130_fd_sc_hd__inv_2 _17894_ (.A(_01370_),
    .Y(_01396_));
 sky130_fd_sc_hd__o221a_1 _17895_ (.A1(\wfg_core_top.cfg_sync_q[6] ),
    .A2(_01372_),
    .B1(_01395_),
    .B2(_01396_),
    .C1(_01387_),
    .X(_01397_));
 sky130_fd_sc_hd__a31o_1 _17896_ (.A1(\wfg_core_top.active_o ),
    .A2(\wfg_core_top.wfg_core.sync_count[6] ),
    .A3(_01394_),
    .B1(_01397_),
    .X(_00478_));
 sky130_fd_sc_hd__o21ai_1 _17897_ (.A1(\wfg_core_top.wfg_core.sync_count[4] ),
    .A2(_01368_),
    .B1(\wfg_core_top.wfg_core.sync_count[5] ),
    .Y(_01398_));
 sky130_fd_sc_hd__o2bb2a_1 _17898_ (.A1_N(_01369_),
    .A2_N(_01398_),
    .B1(_01372_),
    .B2(\wfg_core_top.cfg_sync_q[5] ),
    .X(_01399_));
 sky130_fd_sc_hd__a22o_1 _17899_ (.A1(\wfg_core_top.wfg_core.sync_count[5] ),
    .A2(_01389_),
    .B1(_01387_),
    .B2(_01399_),
    .X(_00477_));
 sky130_fd_sc_hd__or2_1 _17900_ (.A(\wfg_core_top.cfg_sync_q[4] ),
    .B(_01372_),
    .X(_01400_));
 sky130_fd_sc_hd__xnor2_1 _17901_ (.A(\wfg_core_top.wfg_core.sync_count[4] ),
    .B(_01368_),
    .Y(_01401_));
 sky130_fd_sc_hd__a32o_1 _17902_ (.A1(_01387_),
    .A2(_01400_),
    .A3(_01401_),
    .B1(_01389_),
    .B2(\wfg_core_top.wfg_core.sync_count[4] ),
    .X(_00476_));
 sky130_fd_sc_hd__nand2_1 _17903_ (.A(\wfg_core_top.wfg_core.sync_count[3] ),
    .B(_01367_),
    .Y(_01402_));
 sky130_fd_sc_hd__o2bb2a_1 _17904_ (.A1_N(_01368_),
    .A2_N(_01402_),
    .B1(_01372_),
    .B2(\wfg_core_top.cfg_sync_q[3] ),
    .X(_01403_));
 sky130_fd_sc_hd__a22o_1 _17905_ (.A1(\wfg_core_top.wfg_core.sync_count[3] ),
    .A2(_01389_),
    .B1(_01387_),
    .B2(_01403_),
    .X(_00475_));
 sky130_fd_sc_hd__o21ai_1 _17906_ (.A1(\wfg_core_top.wfg_core.sync_count[1] ),
    .A2(\wfg_core_top.wfg_core.sync_count[0] ),
    .B1(\wfg_core_top.wfg_core.sync_count[2] ),
    .Y(_01404_));
 sky130_fd_sc_hd__o2bb2a_1 _17907_ (.A1_N(_01367_),
    .A2_N(_01404_),
    .B1(_01372_),
    .B2(\wfg_core_top.cfg_sync_q[2] ),
    .X(_01405_));
 sky130_fd_sc_hd__a22o_1 _17908_ (.A1(\wfg_core_top.wfg_core.sync_count[2] ),
    .A2(_01389_),
    .B1(_01387_),
    .B2(_01405_),
    .X(_00474_));
 sky130_fd_sc_hd__and2_1 _17909_ (.A(\wfg_core_top.wfg_core.sync_count[1] ),
    .B(\wfg_core_top.wfg_core.sync_count[0] ),
    .X(_01406_));
 sky130_fd_sc_hd__nor2_1 _17910_ (.A(\wfg_core_top.wfg_core.sync_count[1] ),
    .B(\wfg_core_top.wfg_core.sync_count[0] ),
    .Y(_01407_));
 sky130_fd_sc_hd__o22a_1 _17911_ (.A1(\wfg_core_top.cfg_sync_q[1] ),
    .A2(_01372_),
    .B1(_01406_),
    .B2(_01407_),
    .X(_01408_));
 sky130_fd_sc_hd__a22o_1 _17912_ (.A1(\wfg_core_top.wfg_core.sync_count[1] ),
    .A2(_01389_),
    .B1(_01387_),
    .B2(_01408_),
    .X(_00473_));
 sky130_fd_sc_hd__o21ba_1 _17913_ (.A1(\wfg_core_top.cfg_sync_q[0] ),
    .A2(_01372_),
    .B1_N(\wfg_core_top.wfg_core.sync_count[0] ),
    .X(_01409_));
 sky130_fd_sc_hd__a22o_1 _17914_ (.A1(\wfg_core_top.wfg_core.sync_count[0] ),
    .A2(_01389_),
    .B1(_01387_),
    .B2(_01409_),
    .X(_00472_));
 sky130_fd_sc_hd__inv_2 _17915_ (.A(\wfg_stim_mem_top.ctrl_en_q ),
    .Y(net111));
 sky130_fd_sc_hd__a32o_1 _17916_ (.A1(\wfg_stim_mem_top.wfg_stim_mem.cur_state[3] ),
    .A2(_05976_),
    .A3(_05978_),
    .B1(\wfg_stim_mem_top.wfg_stim_mem.cur_state[0] ),
    .B2(net111),
    .X(_00001_));
 sky130_fd_sc_hd__or4_1 _17917_ (.A(\wfg_subcore_top.wbs_ack_o ),
    .B(\wfg_core_top.wbs_ack_o ),
    .C(\wfg_interconnect_top.wbs_ack_o ),
    .D(\wfg_stim_sine_top.wbs_ack_o ),
    .X(_01410_));
 sky130_fd_sc_hd__or4_4 _17918_ (.A(\wfg_stim_mem_top.wbs_ack_o ),
    .B(\wfg_drive_spi_top.wbs_ack_o ),
    .C(\wfg_drive_pat_top.wbs_ack_o ),
    .D(_01410_),
    .X(_01411_));
 sky130_fd_sc_hd__clkbuf_1 _17919_ (.A(_01411_),
    .X(net112));
 sky130_fd_sc_hd__inv_2 _17920_ (.A(net59),
    .Y(_01412_));
 sky130_fd_sc_hd__or4_4 _17921_ (.A(net62),
    .B(net64),
    .C(net63),
    .D(net46),
    .X(_01413_));
 sky130_fd_sc_hd__or4_4 _17922_ (.A(net48),
    .B(net47),
    .C(net52),
    .D(_01413_),
    .X(_01414_));
 sky130_fd_sc_hd__or4_4 _17923_ (.A(net45),
    .B(net50),
    .C(net49),
    .D(net51),
    .X(_01415_));
 sky130_fd_sc_hd__or4_2 _17924_ (.A(net35),
    .B(net34),
    .C(_01414_),
    .D(_01415_),
    .X(_01416_));
 sky130_fd_sc_hd__inv_2 _17925_ (.A(net61),
    .Y(_01417_));
 sky130_fd_sc_hd__or4_1 _17926_ (.A(net41),
    .B(net40),
    .C(net43),
    .D(net42),
    .X(_01418_));
 sky130_fd_sc_hd__or4_1 _17927_ (.A(net37),
    .B(net36),
    .C(net39),
    .D(net38),
    .X(_01419_));
 sky130_fd_sc_hd__or2_2 _17928_ (.A(_01418_),
    .B(_01419_),
    .X(_01420_));
 sky130_fd_sc_hd__inv_2 _17929_ (.A(_01420_),
    .Y(_01421_));
 sky130_fd_sc_hd__and2_1 _17930_ (.A(net60),
    .B(_01421_),
    .X(_01422_));
 sky130_fd_sc_hd__and4bb_1 _17931_ (.A_N(_01412_),
    .B_N(_01416_),
    .C(_01417_),
    .D(_01422_),
    .X(_01423_));
 sky130_fd_sc_hd__or2_2 _17932_ (.A(net60),
    .B(_01420_),
    .X(_01424_));
 sky130_fd_sc_hd__or3_2 _17933_ (.A(net59),
    .B(_01417_),
    .C(_01416_),
    .X(_01425_));
 sky130_fd_sc_hd__nor2_1 _17934_ (.A(_01424_),
    .B(_01425_),
    .Y(_01426_));
 sky130_fd_sc_hd__clkbuf_4 _17935_ (.A(_01426_),
    .X(_01427_));
 sky130_fd_sc_hd__or3_4 _17936_ (.A(_01412_),
    .B(_01417_),
    .C(_01416_),
    .X(_01428_));
 sky130_fd_sc_hd__nor2_4 _17937_ (.A(_01424_),
    .B(_01428_),
    .Y(_01429_));
 sky130_fd_sc_hd__clkbuf_4 _17938_ (.A(_01429_),
    .X(_01430_));
 sky130_fd_sc_hd__nand2_4 _17939_ (.A(net60),
    .B(_01421_),
    .Y(_01431_));
 sky130_fd_sc_hd__nor2_4 _17940_ (.A(_01431_),
    .B(_01425_),
    .Y(_01432_));
 sky130_fd_sc_hd__nor2_4 _17941_ (.A(_01431_),
    .B(_01428_),
    .Y(_01433_));
 sky130_fd_sc_hd__clkbuf_4 _17942_ (.A(_01433_),
    .X(_01434_));
 sky130_fd_sc_hd__a22o_1 _17943_ (.A1(\wfg_drive_spi_top.wbs_dat_o[0] ),
    .A2(_01432_),
    .B1(_01434_),
    .B2(\wfg_drive_pat_top.wbs_dat_o[0] ),
    .X(_01435_));
 sky130_fd_sc_hd__a221o_1 _17944_ (.A1(\wfg_stim_sine_top.wbs_dat_o[0] ),
    .A2(_01427_),
    .B1(_01430_),
    .B2(\wfg_stim_mem_top.wbs_dat_o[0] ),
    .C1(_01435_),
    .X(_01436_));
 sky130_fd_sc_hd__or4_1 _17945_ (.A(net63),
    .B(net35),
    .C(net34),
    .D(net46),
    .X(_01437_));
 sky130_fd_sc_hd__or4_1 _17946_ (.A(net45),
    .B(net48),
    .C(net47),
    .D(net50),
    .X(_01438_));
 sky130_fd_sc_hd__or4_4 _17947_ (.A(net49),
    .B(net52),
    .C(net51),
    .D(_01438_),
    .X(_01439_));
 sky130_fd_sc_hd__or4_1 _17948_ (.A(net62),
    .B(net64),
    .C(_01437_),
    .D(_01439_),
    .X(_01440_));
 sky130_fd_sc_hd__or2_1 _17949_ (.A(_01417_),
    .B(_01440_),
    .X(_01441_));
 sky130_fd_sc_hd__nor2_1 _17950_ (.A(net61),
    .B(_01440_),
    .Y(_01442_));
 sky130_fd_sc_hd__nand2_1 _17951_ (.A(_01422_),
    .B(_01442_),
    .Y(_01443_));
 sky130_fd_sc_hd__o21a_2 _17952_ (.A1(_01420_),
    .A2(_01441_),
    .B1(_01443_),
    .X(_01444_));
 sky130_fd_sc_hd__clkbuf_4 _17953_ (.A(_01444_),
    .X(_01445_));
 sky130_fd_sc_hd__and4b_2 _17954_ (.A_N(_01416_),
    .B(_01417_),
    .C(_01412_),
    .D(_01422_),
    .X(_01446_));
 sky130_fd_sc_hd__clkbuf_4 _17955_ (.A(_01446_),
    .X(_01447_));
 sky130_fd_sc_hd__a22o_1 _17956_ (.A1(\wfg_core_top.wbs_dat_o[0] ),
    .A2(_01445_),
    .B1(_01447_),
    .B2(\wfg_subcore_top.wbs_dat_o[0] ),
    .X(_01448_));
 sky130_fd_sc_hd__a211o_2 _17957_ (.A1(\wfg_interconnect_top.wbs_dat_o[0] ),
    .A2(_01423_),
    .B1(_01436_),
    .C1(_01448_),
    .X(net113));
 sky130_fd_sc_hd__a22o_1 _17958_ (.A1(\wfg_core_top.wbs_dat_o[1] ),
    .A2(_01445_),
    .B1(_01447_),
    .B2(\wfg_subcore_top.wbs_dat_o[1] ),
    .X(_01449_));
 sky130_fd_sc_hd__a22o_1 _17959_ (.A1(\wfg_drive_spi_top.wbs_dat_o[1] ),
    .A2(_01432_),
    .B1(_01434_),
    .B2(\wfg_drive_pat_top.wbs_dat_o[1] ),
    .X(_01450_));
 sky130_fd_sc_hd__a221o_1 _17960_ (.A1(\wfg_stim_sine_top.wbs_dat_o[1] ),
    .A2(_01427_),
    .B1(_01430_),
    .B2(\wfg_stim_mem_top.wbs_dat_o[1] ),
    .C1(_01450_),
    .X(_01451_));
 sky130_fd_sc_hd__a211o_2 _17961_ (.A1(\wfg_interconnect_top.wbs_dat_o[1] ),
    .A2(_01423_),
    .B1(_01449_),
    .C1(_01451_),
    .X(net124));
 sky130_fd_sc_hd__a22o_1 _17962_ (.A1(\wfg_core_top.wbs_dat_o[2] ),
    .A2(_01445_),
    .B1(_01447_),
    .B2(\wfg_subcore_top.wbs_dat_o[2] ),
    .X(_01452_));
 sky130_fd_sc_hd__clkbuf_4 _17963_ (.A(_01433_),
    .X(_01453_));
 sky130_fd_sc_hd__a22o_1 _17964_ (.A1(\wfg_drive_pat_top.wbs_dat_o[2] ),
    .A2(_01453_),
    .B1(_01430_),
    .B2(\wfg_stim_mem_top.wbs_dat_o[2] ),
    .X(_01454_));
 sky130_fd_sc_hd__a21o_1 _17965_ (.A1(\wfg_stim_sine_top.wbs_dat_o[2] ),
    .A2(_01427_),
    .B1(_01454_),
    .X(_01455_));
 sky130_fd_sc_hd__a211o_2 _17966_ (.A1(\wfg_drive_spi_top.wbs_dat_o[2] ),
    .A2(_01432_),
    .B1(_01452_),
    .C1(_01455_),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_4 _17967_ (.A(_01427_),
    .X(_01456_));
 sky130_fd_sc_hd__a22o_1 _17968_ (.A1(\wfg_drive_pat_top.wbs_dat_o[3] ),
    .A2(_01434_),
    .B1(_01429_),
    .B2(\wfg_stim_mem_top.wbs_dat_o[3] ),
    .X(_01457_));
 sky130_fd_sc_hd__a21o_1 _17969_ (.A1(\wfg_drive_spi_top.wbs_dat_o[3] ),
    .A2(_01432_),
    .B1(_01457_),
    .X(_01458_));
 sky130_fd_sc_hd__a22o_1 _17970_ (.A1(\wfg_core_top.wbs_dat_o[3] ),
    .A2(_01445_),
    .B1(_01447_),
    .B2(\wfg_subcore_top.wbs_dat_o[3] ),
    .X(_01459_));
 sky130_fd_sc_hd__a211o_1 _17971_ (.A1(\wfg_stim_sine_top.wbs_dat_o[3] ),
    .A2(_01456_),
    .B1(_01458_),
    .C1(_01459_),
    .X(net138));
 sky130_fd_sc_hd__a22o_1 _17972_ (.A1(\wfg_core_top.wbs_dat_o[4] ),
    .A2(_01445_),
    .B1(_01447_),
    .B2(\wfg_subcore_top.wbs_dat_o[4] ),
    .X(_01460_));
 sky130_fd_sc_hd__a22o_1 _17973_ (.A1(\wfg_drive_pat_top.wbs_dat_o[4] ),
    .A2(_01453_),
    .B1(_01429_),
    .B2(\wfg_stim_mem_top.wbs_dat_o[4] ),
    .X(_01461_));
 sky130_fd_sc_hd__a21o_1 _17974_ (.A1(\wfg_stim_sine_top.wbs_dat_o[4] ),
    .A2(_01427_),
    .B1(_01461_),
    .X(_01462_));
 sky130_fd_sc_hd__a211o_1 _17975_ (.A1(\wfg_drive_spi_top.wbs_dat_o[4] ),
    .A2(_01432_),
    .B1(_01460_),
    .C1(_01462_),
    .X(net139));
 sky130_fd_sc_hd__a22o_1 _17976_ (.A1(\wfg_drive_pat_top.wbs_dat_o[5] ),
    .A2(_01434_),
    .B1(_01429_),
    .B2(\wfg_stim_mem_top.wbs_dat_o[5] ),
    .X(_01463_));
 sky130_fd_sc_hd__a21o_1 _17977_ (.A1(\wfg_drive_spi_top.wbs_dat_o[5] ),
    .A2(_01432_),
    .B1(_01463_),
    .X(_01464_));
 sky130_fd_sc_hd__a22o_1 _17978_ (.A1(\wfg_core_top.wbs_dat_o[5] ),
    .A2(_01445_),
    .B1(_01447_),
    .B2(\wfg_subcore_top.wbs_dat_o[5] ),
    .X(_01465_));
 sky130_fd_sc_hd__a211o_1 _17979_ (.A1(\wfg_stim_sine_top.wbs_dat_o[5] ),
    .A2(_01456_),
    .B1(_01464_),
    .C1(_01465_),
    .X(net140));
 sky130_fd_sc_hd__a22o_1 _17980_ (.A1(\wfg_core_top.wbs_dat_o[6] ),
    .A2(_01445_),
    .B1(_01447_),
    .B2(\wfg_subcore_top.wbs_dat_o[6] ),
    .X(_01466_));
 sky130_fd_sc_hd__a22o_1 _17981_ (.A1(\wfg_drive_pat_top.wbs_dat_o[6] ),
    .A2(_01453_),
    .B1(_01429_),
    .B2(\wfg_stim_mem_top.wbs_dat_o[6] ),
    .X(_01467_));
 sky130_fd_sc_hd__a21o_1 _17982_ (.A1(\wfg_stim_sine_top.wbs_dat_o[6] ),
    .A2(_01427_),
    .B1(_01467_),
    .X(_01468_));
 sky130_fd_sc_hd__a211o_1 _17983_ (.A1(\wfg_drive_spi_top.wbs_dat_o[6] ),
    .A2(_01432_),
    .B1(_01466_),
    .C1(_01468_),
    .X(net141));
 sky130_fd_sc_hd__a22o_1 _17984_ (.A1(\wfg_drive_pat_top.wbs_dat_o[7] ),
    .A2(_01434_),
    .B1(_01429_),
    .B2(\wfg_stim_mem_top.wbs_dat_o[7] ),
    .X(_01469_));
 sky130_fd_sc_hd__a21o_1 _17985_ (.A1(\wfg_drive_spi_top.wbs_dat_o[7] ),
    .A2(_01432_),
    .B1(_01469_),
    .X(_01470_));
 sky130_fd_sc_hd__a22o_1 _17986_ (.A1(\wfg_core_top.wbs_dat_o[7] ),
    .A2(_01445_),
    .B1(_01447_),
    .B2(\wfg_subcore_top.wbs_dat_o[7] ),
    .X(_01471_));
 sky130_fd_sc_hd__a211o_1 _17987_ (.A1(\wfg_stim_sine_top.wbs_dat_o[7] ),
    .A2(_01456_),
    .B1(_01470_),
    .C1(_01471_),
    .X(net142));
 sky130_fd_sc_hd__buf_2 _17988_ (.A(_01430_),
    .X(_01472_));
 sky130_fd_sc_hd__and2_1 _17989_ (.A(\wfg_drive_pat_top.wbs_dat_o[8] ),
    .B(_01434_),
    .X(_01473_));
 sky130_fd_sc_hd__a221o_1 _17990_ (.A1(\wfg_core_top.wbs_dat_o[8] ),
    .A2(_01445_),
    .B1(_01447_),
    .B2(\wfg_subcore_top.wbs_dat_o[8] ),
    .C1(_01473_),
    .X(_01474_));
 sky130_fd_sc_hd__a221o_1 _17991_ (.A1(\wfg_stim_sine_top.wbs_dat_o[8] ),
    .A2(_01456_),
    .B1(_01472_),
    .B2(\wfg_stim_mem_top.wbs_dat_o[8] ),
    .C1(_01474_),
    .X(net143));
 sky130_fd_sc_hd__and2_1 _17992_ (.A(\wfg_drive_pat_top.wbs_dat_o[9] ),
    .B(_01434_),
    .X(_01475_));
 sky130_fd_sc_hd__a221o_1 _17993_ (.A1(\wfg_core_top.wbs_dat_o[9] ),
    .A2(_01445_),
    .B1(_01447_),
    .B2(\wfg_subcore_top.wbs_dat_o[9] ),
    .C1(_01475_),
    .X(_01476_));
 sky130_fd_sc_hd__a221o_1 _17994_ (.A1(\wfg_stim_sine_top.wbs_dat_o[9] ),
    .A2(_01456_),
    .B1(_01472_),
    .B2(\wfg_stim_mem_top.wbs_dat_o[9] ),
    .C1(_01476_),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_4 _17995_ (.A(_01444_),
    .X(_01477_));
 sky130_fd_sc_hd__buf_2 _17996_ (.A(_01446_),
    .X(_01478_));
 sky130_fd_sc_hd__and2_1 _17997_ (.A(\wfg_drive_pat_top.wbs_dat_o[10] ),
    .B(_01434_),
    .X(_01479_));
 sky130_fd_sc_hd__a221o_1 _17998_ (.A1(\wfg_core_top.wbs_dat_o[10] ),
    .A2(_01477_),
    .B1(_01478_),
    .B2(\wfg_subcore_top.wbs_dat_o[10] ),
    .C1(_01479_),
    .X(_01480_));
 sky130_fd_sc_hd__a221o_1 _17999_ (.A1(\wfg_stim_sine_top.wbs_dat_o[10] ),
    .A2(_01456_),
    .B1(_01472_),
    .B2(\wfg_stim_mem_top.wbs_dat_o[10] ),
    .C1(_01480_),
    .X(net114));
 sky130_fd_sc_hd__and2_1 _18000_ (.A(\wfg_drive_pat_top.wbs_dat_o[11] ),
    .B(_01434_),
    .X(_01481_));
 sky130_fd_sc_hd__a221o_1 _18001_ (.A1(\wfg_core_top.wbs_dat_o[11] ),
    .A2(_01477_),
    .B1(_01478_),
    .B2(\wfg_subcore_top.wbs_dat_o[11] ),
    .C1(_01481_),
    .X(_01482_));
 sky130_fd_sc_hd__a221o_1 _18002_ (.A1(\wfg_stim_sine_top.wbs_dat_o[11] ),
    .A2(_01456_),
    .B1(_01472_),
    .B2(\wfg_stim_mem_top.wbs_dat_o[11] ),
    .C1(_01482_),
    .X(net115));
 sky130_fd_sc_hd__and2_1 _18003_ (.A(\wfg_drive_pat_top.wbs_dat_o[12] ),
    .B(_01434_),
    .X(_01483_));
 sky130_fd_sc_hd__a221o_1 _18004_ (.A1(\wfg_core_top.wbs_dat_o[12] ),
    .A2(_01477_),
    .B1(_01478_),
    .B2(\wfg_subcore_top.wbs_dat_o[12] ),
    .C1(_01483_),
    .X(_01484_));
 sky130_fd_sc_hd__a221o_1 _18005_ (.A1(\wfg_stim_sine_top.wbs_dat_o[12] ),
    .A2(_01456_),
    .B1(_01472_),
    .B2(\wfg_stim_mem_top.wbs_dat_o[12] ),
    .C1(_01484_),
    .X(net116));
 sky130_fd_sc_hd__and2_1 _18006_ (.A(\wfg_drive_pat_top.wbs_dat_o[13] ),
    .B(_01433_),
    .X(_01485_));
 sky130_fd_sc_hd__a221o_1 _18007_ (.A1(\wfg_core_top.wbs_dat_o[13] ),
    .A2(_01477_),
    .B1(_01478_),
    .B2(\wfg_subcore_top.wbs_dat_o[13] ),
    .C1(_01485_),
    .X(_01486_));
 sky130_fd_sc_hd__a221o_1 _18008_ (.A1(\wfg_stim_sine_top.wbs_dat_o[13] ),
    .A2(_01456_),
    .B1(_01472_),
    .B2(\wfg_stim_mem_top.wbs_dat_o[13] ),
    .C1(_01486_),
    .X(net117));
 sky130_fd_sc_hd__and2_1 _18009_ (.A(\wfg_drive_pat_top.wbs_dat_o[14] ),
    .B(_01433_),
    .X(_01487_));
 sky130_fd_sc_hd__a221o_1 _18010_ (.A1(\wfg_core_top.wbs_dat_o[14] ),
    .A2(_01477_),
    .B1(_01478_),
    .B2(\wfg_subcore_top.wbs_dat_o[14] ),
    .C1(_01487_),
    .X(_01488_));
 sky130_fd_sc_hd__a221o_1 _18011_ (.A1(\wfg_stim_sine_top.wbs_dat_o[14] ),
    .A2(_01456_),
    .B1(_01472_),
    .B2(\wfg_stim_mem_top.wbs_dat_o[14] ),
    .C1(_01488_),
    .X(net118));
 sky130_fd_sc_hd__and2_1 _18012_ (.A(\wfg_drive_pat_top.wbs_dat_o[15] ),
    .B(_01433_),
    .X(_01489_));
 sky130_fd_sc_hd__a221o_1 _18013_ (.A1(\wfg_core_top.wbs_dat_o[15] ),
    .A2(_01477_),
    .B1(_01478_),
    .B2(\wfg_subcore_top.wbs_dat_o[15] ),
    .C1(_01489_),
    .X(_01490_));
 sky130_fd_sc_hd__a221o_1 _18014_ (.A1(\wfg_stim_sine_top.wbs_dat_o[15] ),
    .A2(_01427_),
    .B1(_01472_),
    .B2(\wfg_stim_mem_top.wbs_dat_o[15] ),
    .C1(_01490_),
    .X(net119));
 sky130_fd_sc_hd__and2_1 _18015_ (.A(\wfg_drive_pat_top.wbs_dat_o[16] ),
    .B(_01433_),
    .X(_01491_));
 sky130_fd_sc_hd__a221o_1 _18016_ (.A1(\wfg_core_top.wbs_dat_o[16] ),
    .A2(_01477_),
    .B1(_01478_),
    .B2(\wfg_subcore_top.wbs_dat_o[16] ),
    .C1(_01491_),
    .X(_01492_));
 sky130_fd_sc_hd__a221o_2 _18017_ (.A1(\wfg_stim_sine_top.wbs_dat_o[16] ),
    .A2(_01427_),
    .B1(_01472_),
    .B2(\wfg_stim_mem_top.wbs_dat_o[16] ),
    .C1(_01492_),
    .X(net120));
 sky130_fd_sc_hd__and2_1 _18018_ (.A(\wfg_drive_pat_top.wbs_dat_o[17] ),
    .B(_01433_),
    .X(_01493_));
 sky130_fd_sc_hd__a221o_1 _18019_ (.A1(\wfg_core_top.wbs_dat_o[17] ),
    .A2(_01477_),
    .B1(_01478_),
    .B2(\wfg_subcore_top.wbs_dat_o[17] ),
    .C1(_01493_),
    .X(_01494_));
 sky130_fd_sc_hd__a221o_2 _18020_ (.A1(\wfg_stim_sine_top.wbs_dat_o[17] ),
    .A2(_01427_),
    .B1(_01472_),
    .B2(\wfg_stim_mem_top.wbs_dat_o[17] ),
    .C1(_01494_),
    .X(net121));
 sky130_fd_sc_hd__a22o_1 _18021_ (.A1(\wfg_subcore_top.wbs_dat_o[18] ),
    .A2(_01478_),
    .B1(_01453_),
    .B2(\wfg_drive_pat_top.wbs_dat_o[18] ),
    .X(_01495_));
 sky130_fd_sc_hd__a22o_1 _18022_ (.A1(\wfg_core_top.wbs_dat_o[18] ),
    .A2(_01477_),
    .B1(_01430_),
    .B2(\wfg_stim_mem_top.wbs_dat_o[18] ),
    .X(_01496_));
 sky130_fd_sc_hd__or2_1 _18023_ (.A(_01495_),
    .B(_01496_),
    .X(_01497_));
 sky130_fd_sc_hd__clkbuf_1 _18024_ (.A(_01497_),
    .X(net122));
 sky130_fd_sc_hd__a22o_1 _18025_ (.A1(\wfg_subcore_top.wbs_dat_o[19] ),
    .A2(_01478_),
    .B1(_01453_),
    .B2(\wfg_drive_pat_top.wbs_dat_o[19] ),
    .X(_01498_));
 sky130_fd_sc_hd__a22o_1 _18026_ (.A1(\wfg_core_top.wbs_dat_o[19] ),
    .A2(_01477_),
    .B1(_01430_),
    .B2(\wfg_stim_mem_top.wbs_dat_o[19] ),
    .X(_01499_));
 sky130_fd_sc_hd__or2_1 _18027_ (.A(_01498_),
    .B(_01499_),
    .X(_01500_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18028_ (.A(_01500_),
    .X(net123));
 sky130_fd_sc_hd__a22o_1 _18029_ (.A1(\wfg_subcore_top.wbs_dat_o[20] ),
    .A2(_01446_),
    .B1(_01453_),
    .B2(\wfg_drive_pat_top.wbs_dat_o[20] ),
    .X(_01501_));
 sky130_fd_sc_hd__a22o_1 _18030_ (.A1(\wfg_core_top.wbs_dat_o[20] ),
    .A2(_01444_),
    .B1(_01430_),
    .B2(\wfg_stim_mem_top.wbs_dat_o[20] ),
    .X(_01502_));
 sky130_fd_sc_hd__or2_1 _18031_ (.A(_01501_),
    .B(_01502_),
    .X(_01503_));
 sky130_fd_sc_hd__clkbuf_1 _18032_ (.A(_01503_),
    .X(net125));
 sky130_fd_sc_hd__a22o_1 _18033_ (.A1(\wfg_subcore_top.wbs_dat_o[21] ),
    .A2(_01446_),
    .B1(_01453_),
    .B2(\wfg_drive_pat_top.wbs_dat_o[21] ),
    .X(_01504_));
 sky130_fd_sc_hd__a22o_1 _18034_ (.A1(\wfg_core_top.wbs_dat_o[21] ),
    .A2(_01444_),
    .B1(_01430_),
    .B2(\wfg_stim_mem_top.wbs_dat_o[21] ),
    .X(_01505_));
 sky130_fd_sc_hd__or2_1 _18035_ (.A(_01504_),
    .B(_01505_),
    .X(_01506_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18036_ (.A(_01506_),
    .X(net126));
 sky130_fd_sc_hd__a22o_1 _18037_ (.A1(\wfg_subcore_top.wbs_dat_o[22] ),
    .A2(_01446_),
    .B1(_01453_),
    .B2(\wfg_drive_pat_top.wbs_dat_o[22] ),
    .X(_01507_));
 sky130_fd_sc_hd__a22o_1 _18038_ (.A1(\wfg_core_top.wbs_dat_o[22] ),
    .A2(_01444_),
    .B1(_01430_),
    .B2(\wfg_stim_mem_top.wbs_dat_o[22] ),
    .X(_01508_));
 sky130_fd_sc_hd__or2_1 _18039_ (.A(_01507_),
    .B(_01508_),
    .X(_01509_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18040_ (.A(_01509_),
    .X(net127));
 sky130_fd_sc_hd__a22o_1 _18041_ (.A1(\wfg_subcore_top.wbs_dat_o[23] ),
    .A2(_01446_),
    .B1(_01453_),
    .B2(\wfg_drive_pat_top.wbs_dat_o[23] ),
    .X(_01510_));
 sky130_fd_sc_hd__a22o_1 _18042_ (.A1(\wfg_core_top.wbs_dat_o[23] ),
    .A2(_01444_),
    .B1(_01430_),
    .B2(\wfg_stim_mem_top.wbs_dat_o[23] ),
    .X(_01511_));
 sky130_fd_sc_hd__or2_1 _18043_ (.A(_01510_),
    .B(_01511_),
    .X(_01512_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18044_ (.A(_01512_),
    .X(net128));
 sky130_fd_sc_hd__inv_2 _18045_ (.A(_01441_),
    .Y(_01513_));
 sky130_fd_sc_hd__and3_4 _18046_ (.A(net59),
    .B(_01422_),
    .C(_01513_),
    .X(_01514_));
 sky130_fd_sc_hd__and2_1 _18047_ (.A(\wfg_drive_pat_top.wbs_dat_o[24] ),
    .B(_01514_),
    .X(_01515_));
 sky130_fd_sc_hd__clkbuf_1 _18048_ (.A(_01515_),
    .X(net129));
 sky130_fd_sc_hd__and2_1 _18049_ (.A(\wfg_drive_pat_top.wbs_dat_o[25] ),
    .B(_01514_),
    .X(_01516_));
 sky130_fd_sc_hd__clkbuf_1 _18050_ (.A(_01516_),
    .X(net130));
 sky130_fd_sc_hd__and2_1 _18051_ (.A(\wfg_drive_pat_top.wbs_dat_o[26] ),
    .B(_01514_),
    .X(_01517_));
 sky130_fd_sc_hd__clkbuf_1 _18052_ (.A(_01517_),
    .X(net131));
 sky130_fd_sc_hd__and2_1 _18053_ (.A(\wfg_drive_pat_top.wbs_dat_o[27] ),
    .B(_01514_),
    .X(_01518_));
 sky130_fd_sc_hd__clkbuf_1 _18054_ (.A(_01518_),
    .X(net132));
 sky130_fd_sc_hd__and2_1 _18055_ (.A(\wfg_drive_pat_top.wbs_dat_o[28] ),
    .B(_01514_),
    .X(_01519_));
 sky130_fd_sc_hd__clkbuf_1 _18056_ (.A(_01519_),
    .X(net133));
 sky130_fd_sc_hd__and2_1 _18057_ (.A(\wfg_drive_pat_top.wbs_dat_o[29] ),
    .B(_01514_),
    .X(_01520_));
 sky130_fd_sc_hd__clkbuf_1 _18058_ (.A(_01520_),
    .X(net134));
 sky130_fd_sc_hd__and2_1 _18059_ (.A(\wfg_drive_pat_top.wbs_dat_o[30] ),
    .B(_01514_),
    .X(_01521_));
 sky130_fd_sc_hd__clkbuf_1 _18060_ (.A(_01521_),
    .X(net136));
 sky130_fd_sc_hd__and2_1 _18061_ (.A(\wfg_drive_pat_top.wbs_dat_o[31] ),
    .B(_01514_),
    .X(_01522_));
 sky130_fd_sc_hd__clkbuf_1 _18062_ (.A(_01522_),
    .X(net137));
 sky130_fd_sc_hd__inv_2 _18063_ (.A(\wfg_core_top.wfg_core.subcycle_count[0] ),
    .Y(_01523_));
 sky130_fd_sc_hd__buf_2 _18064_ (.A(\wfg_core_top.active_o ),
    .X(_01524_));
 sky130_fd_sc_hd__o211a_1 _18065_ (.A1(\wfg_core_top.cfg_subcycle_q[8] ),
    .A2(_01394_),
    .B1(_01523_),
    .C1(_01524_),
    .X(_00004_));
 sky130_fd_sc_hd__and2_1 _18066_ (.A(\wfg_core_top.wfg_core.subcycle_count[1] ),
    .B(\wfg_core_top.wfg_core.subcycle_count[0] ),
    .X(_01525_));
 sky130_fd_sc_hd__nor2_1 _18067_ (.A(\wfg_core_top.wfg_core.subcycle_count[1] ),
    .B(\wfg_core_top.wfg_core.subcycle_count[0] ),
    .Y(_01526_));
 sky130_fd_sc_hd__o221a_1 _18068_ (.A1(\wfg_core_top.cfg_subcycle_q[9] ),
    .A2(_01394_),
    .B1(_01525_),
    .B2(_01526_),
    .C1(_01524_),
    .X(_00011_));
 sky130_fd_sc_hd__o21a_1 _18069_ (.A1(\wfg_core_top.wfg_core.subcycle_count[1] ),
    .A2(\wfg_core_top.wfg_core.subcycle_count[0] ),
    .B1(\wfg_core_top.wfg_core.subcycle_count[2] ),
    .X(_01527_));
 sky130_fd_sc_hd__inv_2 _18070_ (.A(_01373_),
    .Y(_01528_));
 sky130_fd_sc_hd__o221a_1 _18071_ (.A1(\wfg_core_top.cfg_subcycle_q[10] ),
    .A2(_01394_),
    .B1(_01527_),
    .B2(_01528_),
    .C1(_01524_),
    .X(_00012_));
 sky130_fd_sc_hd__and2_1 _18072_ (.A(\wfg_core_top.wfg_core.subcycle_count[3] ),
    .B(_01373_),
    .X(_01529_));
 sky130_fd_sc_hd__inv_2 _18073_ (.A(_01374_),
    .Y(_01530_));
 sky130_fd_sc_hd__o221a_1 _18074_ (.A1(\wfg_core_top.cfg_subcycle_q[11] ),
    .A2(_01394_),
    .B1(_01529_),
    .B2(_01530_),
    .C1(_01524_),
    .X(_00013_));
 sky130_fd_sc_hd__and2_1 _18075_ (.A(\wfg_core_top.wfg_core.subcycle_count[4] ),
    .B(_01374_),
    .X(_01531_));
 sky130_fd_sc_hd__nor2_1 _18076_ (.A(\wfg_core_top.wfg_core.subcycle_count[4] ),
    .B(_01374_),
    .Y(_01532_));
 sky130_fd_sc_hd__o221a_1 _18077_ (.A1(\wfg_core_top.cfg_subcycle_q[12] ),
    .A2(_01394_),
    .B1(_01531_),
    .B2(_01532_),
    .C1(_01524_),
    .X(_00014_));
 sky130_fd_sc_hd__o21a_1 _18078_ (.A1(\wfg_core_top.wfg_core.subcycle_count[4] ),
    .A2(_01374_),
    .B1(\wfg_core_top.wfg_core.subcycle_count[5] ),
    .X(_01533_));
 sky130_fd_sc_hd__inv_2 _18079_ (.A(_01375_),
    .Y(_01534_));
 sky130_fd_sc_hd__o221a_1 _18080_ (.A1(\wfg_core_top.cfg_subcycle_q[13] ),
    .A2(_01394_),
    .B1(_01533_),
    .B2(_01534_),
    .C1(_01524_),
    .X(_00015_));
 sky130_fd_sc_hd__nand2_1 _18081_ (.A(\wfg_core_top.wfg_core.subcycle_count[6] ),
    .B(_01375_),
    .Y(_01535_));
 sky130_fd_sc_hd__nand2_1 _18082_ (.A(_01376_),
    .B(_01535_),
    .Y(_01536_));
 sky130_fd_sc_hd__o211a_1 _18083_ (.A1(\wfg_core_top.cfg_subcycle_q[14] ),
    .A2(_01394_),
    .B1(_01536_),
    .C1(_01524_),
    .X(_00016_));
 sky130_fd_sc_hd__and2_1 _18084_ (.A(\wfg_core_top.wfg_core.subcycle_count[7] ),
    .B(_01376_),
    .X(_01537_));
 sky130_fd_sc_hd__nor2_1 _18085_ (.A(\wfg_core_top.wfg_core.subcycle_count[7] ),
    .B(_01376_),
    .Y(_01538_));
 sky130_fd_sc_hd__o221a_1 _18086_ (.A1(\wfg_core_top.cfg_subcycle_q[15] ),
    .A2(_01394_),
    .B1(_01537_),
    .B2(_01538_),
    .C1(_01524_),
    .X(_00017_));
 sky130_fd_sc_hd__o21a_1 _18087_ (.A1(\wfg_core_top.wfg_core.subcycle_count[7] ),
    .A2(_01376_),
    .B1(\wfg_core_top.wfg_core.subcycle_count[8] ),
    .X(_01539_));
 sky130_fd_sc_hd__inv_2 _18088_ (.A(_01377_),
    .Y(_01540_));
 sky130_fd_sc_hd__o221a_1 _18089_ (.A1(\wfg_core_top.cfg_subcycle_q[16] ),
    .A2(_01384_),
    .B1(_01539_),
    .B2(_01540_),
    .C1(_01524_),
    .X(_00018_));
 sky130_fd_sc_hd__nand2_1 _18090_ (.A(\wfg_core_top.wfg_core.subcycle_count[9] ),
    .B(_01377_),
    .Y(_01541_));
 sky130_fd_sc_hd__nand2_1 _18091_ (.A(_01378_),
    .B(_01541_),
    .Y(_01542_));
 sky130_fd_sc_hd__o211a_1 _18092_ (.A1(\wfg_core_top.cfg_subcycle_q[17] ),
    .A2(_01394_),
    .B1(_01542_),
    .C1(_01524_),
    .X(_00019_));
 sky130_fd_sc_hd__and2_1 _18093_ (.A(\wfg_core_top.wfg_core.subcycle_count[10] ),
    .B(_01378_),
    .X(_01543_));
 sky130_fd_sc_hd__nor2_1 _18094_ (.A(\wfg_core_top.wfg_core.subcycle_count[10] ),
    .B(_01378_),
    .Y(_01544_));
 sky130_fd_sc_hd__o221a_1 _18095_ (.A1(\wfg_core_top.cfg_subcycle_q[18] ),
    .A2(_01384_),
    .B1(_01543_),
    .B2(_01544_),
    .C1(\wfg_core_top.active_o ),
    .X(_00005_));
 sky130_fd_sc_hd__o21a_1 _18096_ (.A1(\wfg_core_top.wfg_core.subcycle_count[10] ),
    .A2(_01378_),
    .B1(\wfg_core_top.wfg_core.subcycle_count[11] ),
    .X(_01545_));
 sky130_fd_sc_hd__inv_2 _18097_ (.A(_01379_),
    .Y(_01546_));
 sky130_fd_sc_hd__o221a_1 _18098_ (.A1(\wfg_core_top.cfg_subcycle_q[19] ),
    .A2(_01384_),
    .B1(_01545_),
    .B2(_01546_),
    .C1(\wfg_core_top.active_o ),
    .X(_00006_));
 sky130_fd_sc_hd__nand2_1 _18099_ (.A(\wfg_core_top.wfg_core.subcycle_count[12] ),
    .B(_01379_),
    .Y(_01547_));
 sky130_fd_sc_hd__a2bb2o_1 _18100_ (.A1_N(\wfg_core_top.cfg_subcycle_q[20] ),
    .A2_N(_01384_),
    .B1(_01547_),
    .B2(_01380_),
    .X(_01548_));
 sky130_fd_sc_hd__nor2_1 _18101_ (.A(_01351_),
    .B(_01548_),
    .Y(_00007_));
 sky130_fd_sc_hd__nand2_1 _18102_ (.A(\wfg_core_top.wfg_core.subcycle_count[13] ),
    .B(_01380_),
    .Y(_01549_));
 sky130_fd_sc_hd__a2bb2o_1 _18103_ (.A1_N(\wfg_core_top.cfg_subcycle_q[21] ),
    .A2_N(_01384_),
    .B1(_01549_),
    .B2(_01381_),
    .X(_01550_));
 sky130_fd_sc_hd__nor2_1 _18104_ (.A(_01351_),
    .B(_01550_),
    .Y(_00008_));
 sky130_fd_sc_hd__o21ba_1 _18105_ (.A1(\wfg_core_top.cfg_subcycle_q[22] ),
    .A2(\wfg_core_top.wfg_core.subcycle_count[15] ),
    .B1_N(_01382_),
    .X(_01551_));
 sky130_fd_sc_hd__a21oi_1 _18106_ (.A1(\wfg_core_top.wfg_core.subcycle_count[14] ),
    .A2(_01381_),
    .B1(_01551_),
    .Y(_01552_));
 sky130_fd_sc_hd__nor2_1 _18107_ (.A(_01351_),
    .B(_01552_),
    .Y(_00009_));
 sky130_fd_sc_hd__and3_1 _18108_ (.A(\wfg_core_top.active_o ),
    .B(\wfg_core_top.wfg_core.subcycle_count[15] ),
    .C(_01382_),
    .X(_01553_));
 sky130_fd_sc_hd__a21o_1 _18109_ (.A1(\wfg_core_top.cfg_subcycle_q[23] ),
    .A2(_01387_),
    .B1(_01553_),
    .X(_00010_));
 sky130_fd_sc_hd__clkbuf_4 _18110_ (.A(_09751_),
    .X(_01554_));
 sky130_fd_sc_hd__inv_2 _18111_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_count[0] ),
    .Y(_01555_));
 sky130_fd_sc_hd__clkbuf_4 _18112_ (.A(\wfg_subcore_top.active_o ),
    .X(_01556_));
 sky130_fd_sc_hd__o211a_1 _18113_ (.A1(\wfg_subcore_top.cfg_subcycle_q[8] ),
    .A2(_01554_),
    .B1(_01555_),
    .C1(_01556_),
    .X(_00024_));
 sky130_fd_sc_hd__and2_1 _18114_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_count[1] ),
    .B(\wfg_subcore_top.wfg_subcore.subcycle_count[0] ),
    .X(_01557_));
 sky130_fd_sc_hd__nor2_1 _18115_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_count[1] ),
    .B(\wfg_subcore_top.wfg_subcore.subcycle_count[0] ),
    .Y(_01558_));
 sky130_fd_sc_hd__o221a_1 _18116_ (.A1(\wfg_subcore_top.cfg_subcycle_q[9] ),
    .A2(_01554_),
    .B1(_01557_),
    .B2(_01558_),
    .C1(_01556_),
    .X(_00031_));
 sky130_fd_sc_hd__o21a_1 _18117_ (.A1(\wfg_subcore_top.wfg_subcore.subcycle_count[1] ),
    .A2(\wfg_subcore_top.wfg_subcore.subcycle_count[0] ),
    .B1(\wfg_subcore_top.wfg_subcore.subcycle_count[2] ),
    .X(_01559_));
 sky130_fd_sc_hd__inv_2 _18118_ (.A(_09740_),
    .Y(_01560_));
 sky130_fd_sc_hd__o221a_1 _18119_ (.A1(\wfg_subcore_top.cfg_subcycle_q[10] ),
    .A2(_01554_),
    .B1(_01559_),
    .B2(_01560_),
    .C1(_01556_),
    .X(_00032_));
 sky130_fd_sc_hd__and2_1 _18120_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_count[3] ),
    .B(_09740_),
    .X(_01561_));
 sky130_fd_sc_hd__inv_2 _18121_ (.A(_09741_),
    .Y(_01562_));
 sky130_fd_sc_hd__o221a_1 _18122_ (.A1(\wfg_subcore_top.cfg_subcycle_q[11] ),
    .A2(_01554_),
    .B1(_01561_),
    .B2(_01562_),
    .C1(_01556_),
    .X(_00033_));
 sky130_fd_sc_hd__and2_1 _18123_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_count[4] ),
    .B(_09741_),
    .X(_01563_));
 sky130_fd_sc_hd__nor2_1 _18124_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_count[4] ),
    .B(_09741_),
    .Y(_01564_));
 sky130_fd_sc_hd__o221a_1 _18125_ (.A1(\wfg_subcore_top.cfg_subcycle_q[12] ),
    .A2(_01554_),
    .B1(_01563_),
    .B2(_01564_),
    .C1(_01556_),
    .X(_00034_));
 sky130_fd_sc_hd__o21a_1 _18126_ (.A1(\wfg_subcore_top.wfg_subcore.subcycle_count[4] ),
    .A2(_09741_),
    .B1(\wfg_subcore_top.wfg_subcore.subcycle_count[5] ),
    .X(_01565_));
 sky130_fd_sc_hd__inv_2 _18127_ (.A(_09742_),
    .Y(_01566_));
 sky130_fd_sc_hd__o221a_1 _18128_ (.A1(\wfg_subcore_top.cfg_subcycle_q[13] ),
    .A2(_01554_),
    .B1(_01565_),
    .B2(_01566_),
    .C1(_01556_),
    .X(_00035_));
 sky130_fd_sc_hd__nand2_1 _18129_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_count[6] ),
    .B(_09742_),
    .Y(_01567_));
 sky130_fd_sc_hd__nand2_1 _18130_ (.A(_09743_),
    .B(_01567_),
    .Y(_01568_));
 sky130_fd_sc_hd__o211a_1 _18131_ (.A1(\wfg_subcore_top.cfg_subcycle_q[14] ),
    .A2(_01554_),
    .B1(_01568_),
    .C1(_01556_),
    .X(_00036_));
 sky130_fd_sc_hd__and2_1 _18132_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_count[7] ),
    .B(_09743_),
    .X(_01569_));
 sky130_fd_sc_hd__nor2_1 _18133_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_count[7] ),
    .B(_09743_),
    .Y(_01570_));
 sky130_fd_sc_hd__o221a_1 _18134_ (.A1(\wfg_subcore_top.cfg_subcycle_q[15] ),
    .A2(_01554_),
    .B1(_01569_),
    .B2(_01570_),
    .C1(_01556_),
    .X(_00037_));
 sky130_fd_sc_hd__o21a_1 _18135_ (.A1(\wfg_subcore_top.wfg_subcore.subcycle_count[7] ),
    .A2(_09743_),
    .B1(\wfg_subcore_top.wfg_subcore.subcycle_count[8] ),
    .X(_01571_));
 sky130_fd_sc_hd__inv_2 _18136_ (.A(_09744_),
    .Y(_01572_));
 sky130_fd_sc_hd__o221a_1 _18137_ (.A1(\wfg_subcore_top.cfg_subcycle_q[16] ),
    .A2(_01554_),
    .B1(_01571_),
    .B2(_01572_),
    .C1(_01556_),
    .X(_00038_));
 sky130_fd_sc_hd__nand2_1 _18138_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_count[9] ),
    .B(_09744_),
    .Y(_01573_));
 sky130_fd_sc_hd__nand2_1 _18139_ (.A(_09745_),
    .B(_01573_),
    .Y(_01574_));
 sky130_fd_sc_hd__o211a_1 _18140_ (.A1(\wfg_subcore_top.cfg_subcycle_q[17] ),
    .A2(_01554_),
    .B1(_01574_),
    .C1(_01556_),
    .X(_00039_));
 sky130_fd_sc_hd__and2_1 _18141_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_count[10] ),
    .B(_09745_),
    .X(_01575_));
 sky130_fd_sc_hd__nor2_1 _18142_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_count[10] ),
    .B(_09745_),
    .Y(_01576_));
 sky130_fd_sc_hd__o221a_1 _18143_ (.A1(\wfg_subcore_top.cfg_subcycle_q[18] ),
    .A2(_09751_),
    .B1(_01575_),
    .B2(_01576_),
    .C1(\wfg_subcore_top.active_o ),
    .X(_00025_));
 sky130_fd_sc_hd__o21a_1 _18144_ (.A1(\wfg_subcore_top.wfg_subcore.subcycle_count[10] ),
    .A2(_09745_),
    .B1(\wfg_subcore_top.wfg_subcore.subcycle_count[11] ),
    .X(_01577_));
 sky130_fd_sc_hd__inv_2 _18145_ (.A(_09746_),
    .Y(_01578_));
 sky130_fd_sc_hd__o221a_1 _18146_ (.A1(\wfg_subcore_top.cfg_subcycle_q[19] ),
    .A2(_09751_),
    .B1(_01577_),
    .B2(_01578_),
    .C1(\wfg_subcore_top.active_o ),
    .X(_00026_));
 sky130_fd_sc_hd__nand2_1 _18147_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_count[12] ),
    .B(_09746_),
    .Y(_01579_));
 sky130_fd_sc_hd__a2bb2o_1 _18148_ (.A1_N(\wfg_subcore_top.cfg_subcycle_q[20] ),
    .A2_N(_09751_),
    .B1(_01579_),
    .B2(_09747_),
    .X(_01580_));
 sky130_fd_sc_hd__nor2_1 _18149_ (.A(_09712_),
    .B(_01580_),
    .Y(_00027_));
 sky130_fd_sc_hd__nand2_1 _18150_ (.A(\wfg_subcore_top.wfg_subcore.subcycle_count[13] ),
    .B(_09747_),
    .Y(_01581_));
 sky130_fd_sc_hd__a2bb2o_1 _18151_ (.A1_N(\wfg_subcore_top.cfg_subcycle_q[21] ),
    .A2_N(_09751_),
    .B1(_01581_),
    .B2(_09748_),
    .X(_01582_));
 sky130_fd_sc_hd__nor2_1 _18152_ (.A(_09712_),
    .B(_01582_),
    .Y(_00028_));
 sky130_fd_sc_hd__o21ba_1 _18153_ (.A1(\wfg_subcore_top.cfg_subcycle_q[22] ),
    .A2(\wfg_subcore_top.wfg_subcore.subcycle_count[15] ),
    .B1_N(_09749_),
    .X(_01583_));
 sky130_fd_sc_hd__a21oi_1 _18154_ (.A1(\wfg_subcore_top.wfg_subcore.subcycle_count[14] ),
    .A2(_09748_),
    .B1(_01583_),
    .Y(_01584_));
 sky130_fd_sc_hd__nor2_1 _18155_ (.A(_09712_),
    .B(_01584_),
    .Y(_00029_));
 sky130_fd_sc_hd__and3_1 _18156_ (.A(\wfg_subcore_top.active_o ),
    .B(\wfg_subcore_top.wfg_subcore.subcycle_count[15] ),
    .C(_09749_),
    .X(_01585_));
 sky130_fd_sc_hd__a21o_1 _18157_ (.A1(\wfg_subcore_top.cfg_subcycle_q[23] ),
    .A2(_09754_),
    .B1(_01585_),
    .X(_00030_));
 sky130_fd_sc_hd__xor2_1 _18158_ (.A(\wfg_drive_spi_top.wfg_drive_spi.cpol ),
    .B(\wfg_drive_spi_top.wfg_drive_spi.spi_clk ),
    .X(_00021_));
 sky130_fd_sc_hd__xnor2_1 _18159_ (.A(\wfg_drive_spi_top.wfg_drive_spi.cspol ),
    .B(\wfg_drive_spi_top.wfg_drive_spi.spi_cs ),
    .Y(_00020_));
 sky130_fd_sc_hd__mux4_1 _18160_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[7] ),
    .A1(\wfg_drive_spi_top.wfg_drive_spi.spi_data[15] ),
    .A2(\wfg_drive_spi_top.wfg_drive_spi.spi_data[23] ),
    .A3(\wfg_drive_spi_top.wfg_drive_spi.spi_data[31] ),
    .S0(\wfg_drive_spi_top.wfg_drive_spi.byte_cnt[0] ),
    .S1(\wfg_drive_spi_top.wfg_drive_spi.byte_cnt[1] ),
    .X(_01586_));
 sky130_fd_sc_hd__mux2_1 _18161_ (.A0(\wfg_drive_spi_top.wfg_drive_spi.spi_data[0] ),
    .A1(_01586_),
    .S(_02739_),
    .X(_01587_));
 sky130_fd_sc_hd__clkbuf_1 _18162_ (.A(_01587_),
    .X(_00022_));
 sky130_fd_sc_hd__clkinv_4 _18163_ (.A(net98),
    .Y(_01588_));
 sky130_fd_sc_hd__buf_4 _18164_ (.A(_01588_),
    .X(_01589_));
 sky130_fd_sc_hd__clkbuf_4 _18165_ (.A(_01589_),
    .X(_00040_));
 sky130_fd_sc_hd__buf_6 _18166_ (.A(net98),
    .X(_01590_));
 sky130_fd_sc_hd__buf_6 _18167_ (.A(_01590_),
    .X(_01591_));
 sky130_fd_sc_hd__buf_4 _18168_ (.A(_01591_),
    .X(_01592_));
 sky130_fd_sc_hd__inv_2 _18169_ (.A(_01592_),
    .Y(_00041_));
 sky130_fd_sc_hd__inv_2 _18170_ (.A(_01592_),
    .Y(_00042_));
 sky130_fd_sc_hd__inv_2 _18171_ (.A(_01592_),
    .Y(_00043_));
 sky130_fd_sc_hd__inv_2 _18172_ (.A(_01592_),
    .Y(_00044_));
 sky130_fd_sc_hd__inv_2 _18173_ (.A(_01592_),
    .Y(_00045_));
 sky130_fd_sc_hd__inv_2 _18174_ (.A(_01592_),
    .Y(_00046_));
 sky130_fd_sc_hd__inv_2 _18175_ (.A(_01592_),
    .Y(_00047_));
 sky130_fd_sc_hd__inv_2 _18176_ (.A(_01592_),
    .Y(_00048_));
 sky130_fd_sc_hd__inv_2 _18177_ (.A(_01592_),
    .Y(_00049_));
 sky130_fd_sc_hd__inv_2 _18178_ (.A(_01592_),
    .Y(_00050_));
 sky130_fd_sc_hd__buf_4 _18179_ (.A(_01591_),
    .X(_01593_));
 sky130_fd_sc_hd__inv_2 _18180_ (.A(_01593_),
    .Y(_00051_));
 sky130_fd_sc_hd__inv_2 _18181_ (.A(_01593_),
    .Y(_00052_));
 sky130_fd_sc_hd__inv_2 _18182_ (.A(_01593_),
    .Y(_00053_));
 sky130_fd_sc_hd__inv_2 _18183_ (.A(_01593_),
    .Y(_00054_));
 sky130_fd_sc_hd__inv_2 _18184_ (.A(_01593_),
    .Y(_00055_));
 sky130_fd_sc_hd__inv_2 _18185_ (.A(_01593_),
    .Y(_00056_));
 sky130_fd_sc_hd__inv_2 _18186_ (.A(_01593_),
    .Y(_00057_));
 sky130_fd_sc_hd__inv_2 _18187_ (.A(_01593_),
    .Y(_00058_));
 sky130_fd_sc_hd__inv_2 _18188_ (.A(_01593_),
    .Y(_00059_));
 sky130_fd_sc_hd__inv_2 _18189_ (.A(_01593_),
    .Y(_00060_));
 sky130_fd_sc_hd__buf_6 _18190_ (.A(_01591_),
    .X(_01594_));
 sky130_fd_sc_hd__inv_2 _18191_ (.A(_01594_),
    .Y(_00061_));
 sky130_fd_sc_hd__inv_2 _18192_ (.A(_01594_),
    .Y(_00062_));
 sky130_fd_sc_hd__inv_2 _18193_ (.A(_01594_),
    .Y(_00063_));
 sky130_fd_sc_hd__inv_2 _18194_ (.A(_01594_),
    .Y(_00064_));
 sky130_fd_sc_hd__inv_2 _18195_ (.A(_01594_),
    .Y(_00065_));
 sky130_fd_sc_hd__mux2_1 _18196_ (.A0(\wfg_core_top.wfg_core.temp_subcycle ),
    .A1(\wfg_core_top.wfg_core.subcycle_dly ),
    .S(_01590_),
    .X(_01595_));
 sky130_fd_sc_hd__clkbuf_1 _18197_ (.A(_01595_),
    .X(_00482_));
 sky130_fd_sc_hd__mux2_1 _18198_ (.A0(\wfg_core_top.wfg_core.temp_sync ),
    .A1(\wfg_core_top.wfg_core.sync_dly ),
    .S(_01590_),
    .X(_01596_));
 sky130_fd_sc_hd__clkbuf_1 _18199_ (.A(_01596_),
    .X(_00483_));
 sky130_fd_sc_hd__inv_2 _18200_ (.A(_01594_),
    .Y(_00066_));
 sky130_fd_sc_hd__inv_2 _18201_ (.A(_01594_),
    .Y(_00067_));
 sky130_fd_sc_hd__inv_2 _18202_ (.A(_01594_),
    .Y(_00068_));
 sky130_fd_sc_hd__inv_2 _18203_ (.A(_01594_),
    .Y(_00069_));
 sky130_fd_sc_hd__inv_2 _18204_ (.A(_01594_),
    .Y(_00070_));
 sky130_fd_sc_hd__buf_6 _18205_ (.A(_01590_),
    .X(_01597_));
 sky130_fd_sc_hd__buf_6 _18206_ (.A(_01597_),
    .X(_01598_));
 sky130_fd_sc_hd__inv_2 _18207_ (.A(_01598_),
    .Y(_00071_));
 sky130_fd_sc_hd__inv_2 _18208_ (.A(_01598_),
    .Y(_00072_));
 sky130_fd_sc_hd__inv_2 _18209_ (.A(_01598_),
    .Y(_00073_));
 sky130_fd_sc_hd__buf_6 _18210_ (.A(_01588_),
    .X(_01599_));
 sky130_fd_sc_hd__buf_4 _18211_ (.A(_01599_),
    .X(_01600_));
 sky130_fd_sc_hd__buf_8 _18212_ (.A(net96),
    .X(_01601_));
 sky130_fd_sc_hd__or2_2 _18213_ (.A(net33),
    .B(net44),
    .X(_01602_));
 sky130_fd_sc_hd__or2b_1 _18214_ (.A(net58),
    .B_N(net55),
    .X(_01603_));
 sky130_fd_sc_hd__or2_4 _18215_ (.A(_01602_),
    .B(_01603_),
    .X(_01604_));
 sky130_fd_sc_hd__nand2_2 _18216_ (.A(net100),
    .B(net65),
    .Y(_01605_));
 sky130_fd_sc_hd__nand2_1 _18217_ (.A(net99),
    .B(net53),
    .Y(_01606_));
 sky130_fd_sc_hd__or4b_4 _18218_ (.A(net57),
    .B(net56),
    .C(_01606_),
    .D_N(net54),
    .X(_01607_));
 sky130_fd_sc_hd__nor2_2 _18219_ (.A(_01412_),
    .B(_01424_),
    .Y(_01608_));
 sky130_fd_sc_hd__or3_1 _18220_ (.A(net63),
    .B(net35),
    .C(net34),
    .X(_01609_));
 sky130_fd_sc_hd__nor3_1 _18221_ (.A(net62),
    .B(net64),
    .C(_01609_),
    .Y(_01610_));
 sky130_fd_sc_hd__or4_1 _18222_ (.A(net50),
    .B(net49),
    .C(net52),
    .D(net51),
    .X(_01611_));
 sky130_fd_sc_hd__or4_1 _18223_ (.A(net46),
    .B(net45),
    .C(net48),
    .D(net47),
    .X(_01612_));
 sky130_fd_sc_hd__nor2_4 _18224_ (.A(_01611_),
    .B(_01612_),
    .Y(_01613_));
 sky130_fd_sc_hd__and4_1 _18225_ (.A(_01417_),
    .B(_01608_),
    .C(_01610_),
    .D(_01613_),
    .X(_01614_));
 sky130_fd_sc_hd__or4b_1 _18226_ (.A(_01604_),
    .B(_01605_),
    .C(_01607_),
    .D_N(_01614_),
    .X(_01615_));
 sky130_fd_sc_hd__buf_2 _18227_ (.A(_01615_),
    .X(_01616_));
 sky130_fd_sc_hd__clkbuf_4 _18228_ (.A(_01616_),
    .X(_01617_));
 sky130_fd_sc_hd__mux2_1 _18229_ (.A0(_01601_),
    .A1(\wfg_core_top.cfg_subcycle_q[8] ),
    .S(_01617_),
    .X(_01618_));
 sky130_fd_sc_hd__and2_1 _18230_ (.A(_01600_),
    .B(_01618_),
    .X(_01619_));
 sky130_fd_sc_hd__clkbuf_1 _18231_ (.A(_01619_),
    .X(_00492_));
 sky130_fd_sc_hd__buf_6 _18232_ (.A(net97),
    .X(_01620_));
 sky130_fd_sc_hd__mux2_1 _18233_ (.A0(_01620_),
    .A1(\wfg_core_top.cfg_subcycle_q[9] ),
    .S(_01617_),
    .X(_01621_));
 sky130_fd_sc_hd__and2_1 _18234_ (.A(_01600_),
    .B(_01621_),
    .X(_01622_));
 sky130_fd_sc_hd__clkbuf_1 _18235_ (.A(_01622_),
    .X(_00493_));
 sky130_fd_sc_hd__buf_2 _18236_ (.A(_01599_),
    .X(_01623_));
 sky130_fd_sc_hd__buf_6 _18237_ (.A(net67),
    .X(_01624_));
 sky130_fd_sc_hd__mux2_1 _18238_ (.A0(_01624_),
    .A1(\wfg_core_top.cfg_subcycle_q[10] ),
    .S(_01617_),
    .X(_01625_));
 sky130_fd_sc_hd__and2_1 _18239_ (.A(_01623_),
    .B(_01625_),
    .X(_01626_));
 sky130_fd_sc_hd__clkbuf_1 _18240_ (.A(_01626_),
    .X(_00494_));
 sky130_fd_sc_hd__buf_6 _18241_ (.A(net68),
    .X(_01627_));
 sky130_fd_sc_hd__mux2_1 _18242_ (.A0(_01627_),
    .A1(\wfg_core_top.cfg_subcycle_q[11] ),
    .S(_01617_),
    .X(_01628_));
 sky130_fd_sc_hd__and2_1 _18243_ (.A(_01623_),
    .B(_01628_),
    .X(_01629_));
 sky130_fd_sc_hd__clkbuf_1 _18244_ (.A(_01629_),
    .X(_00495_));
 sky130_fd_sc_hd__buf_8 _18245_ (.A(net69),
    .X(_01630_));
 sky130_fd_sc_hd__mux2_1 _18246_ (.A0(_01630_),
    .A1(\wfg_core_top.cfg_subcycle_q[12] ),
    .S(_01617_),
    .X(_01631_));
 sky130_fd_sc_hd__and2_1 _18247_ (.A(_01623_),
    .B(_01631_),
    .X(_01632_));
 sky130_fd_sc_hd__clkbuf_1 _18248_ (.A(_01632_),
    .X(_00496_));
 sky130_fd_sc_hd__buf_8 _18249_ (.A(net70),
    .X(_01633_));
 sky130_fd_sc_hd__mux2_1 _18250_ (.A0(_01633_),
    .A1(\wfg_core_top.cfg_subcycle_q[13] ),
    .S(_01617_),
    .X(_01634_));
 sky130_fd_sc_hd__and2_1 _18251_ (.A(_01623_),
    .B(_01634_),
    .X(_01635_));
 sky130_fd_sc_hd__clkbuf_1 _18252_ (.A(_01635_),
    .X(_00497_));
 sky130_fd_sc_hd__buf_8 _18253_ (.A(net71),
    .X(_01636_));
 sky130_fd_sc_hd__mux2_1 _18254_ (.A0(_01636_),
    .A1(\wfg_core_top.cfg_subcycle_q[14] ),
    .S(_01617_),
    .X(_01637_));
 sky130_fd_sc_hd__and2_1 _18255_ (.A(_01623_),
    .B(_01637_),
    .X(_01638_));
 sky130_fd_sc_hd__clkbuf_1 _18256_ (.A(_01638_),
    .X(_00498_));
 sky130_fd_sc_hd__buf_8 _18257_ (.A(net72),
    .X(_01639_));
 sky130_fd_sc_hd__mux2_1 _18258_ (.A0(_01639_),
    .A1(\wfg_core_top.cfg_subcycle_q[15] ),
    .S(_01617_),
    .X(_01640_));
 sky130_fd_sc_hd__and2_1 _18259_ (.A(_01623_),
    .B(_01640_),
    .X(_01641_));
 sky130_fd_sc_hd__clkbuf_1 _18260_ (.A(_01641_),
    .X(_00499_));
 sky130_fd_sc_hd__mux2_1 _18261_ (.A0(net73),
    .A1(\wfg_core_top.cfg_subcycle_q[16] ),
    .S(_01617_),
    .X(_01642_));
 sky130_fd_sc_hd__and2_1 _18262_ (.A(_01623_),
    .B(_01642_),
    .X(_01643_));
 sky130_fd_sc_hd__clkbuf_1 _18263_ (.A(_01643_),
    .X(_00500_));
 sky130_fd_sc_hd__mux2_1 _18264_ (.A0(net74),
    .A1(\wfg_core_top.cfg_subcycle_q[17] ),
    .S(_01617_),
    .X(_01644_));
 sky130_fd_sc_hd__and2_1 _18265_ (.A(_01623_),
    .B(_01644_),
    .X(_01645_));
 sky130_fd_sc_hd__clkbuf_1 _18266_ (.A(_01645_),
    .X(_00501_));
 sky130_fd_sc_hd__clkbuf_4 _18267_ (.A(_01616_),
    .X(_01646_));
 sky130_fd_sc_hd__mux2_1 _18268_ (.A0(net75),
    .A1(\wfg_core_top.cfg_subcycle_q[18] ),
    .S(_01646_),
    .X(_01647_));
 sky130_fd_sc_hd__and2_1 _18269_ (.A(_01623_),
    .B(_01647_),
    .X(_01648_));
 sky130_fd_sc_hd__clkbuf_1 _18270_ (.A(_01648_),
    .X(_00502_));
 sky130_fd_sc_hd__mux2_1 _18271_ (.A0(net76),
    .A1(\wfg_core_top.cfg_subcycle_q[19] ),
    .S(_01646_),
    .X(_01649_));
 sky130_fd_sc_hd__and2_1 _18272_ (.A(_01623_),
    .B(_01649_),
    .X(_01650_));
 sky130_fd_sc_hd__clkbuf_1 _18273_ (.A(_01650_),
    .X(_00503_));
 sky130_fd_sc_hd__clkbuf_2 _18274_ (.A(_01599_),
    .X(_01651_));
 sky130_fd_sc_hd__mux2_1 _18275_ (.A0(net78),
    .A1(\wfg_core_top.cfg_subcycle_q[20] ),
    .S(_01646_),
    .X(_01652_));
 sky130_fd_sc_hd__and2_1 _18276_ (.A(_01651_),
    .B(_01652_),
    .X(_01653_));
 sky130_fd_sc_hd__clkbuf_1 _18277_ (.A(_01653_),
    .X(_00504_));
 sky130_fd_sc_hd__mux2_1 _18278_ (.A0(net79),
    .A1(\wfg_core_top.cfg_subcycle_q[21] ),
    .S(_01646_),
    .X(_01654_));
 sky130_fd_sc_hd__and2_1 _18279_ (.A(_01651_),
    .B(_01654_),
    .X(_01655_));
 sky130_fd_sc_hd__clkbuf_1 _18280_ (.A(_01655_),
    .X(_00505_));
 sky130_fd_sc_hd__mux2_1 _18281_ (.A0(net80),
    .A1(\wfg_core_top.cfg_subcycle_q[22] ),
    .S(_01646_),
    .X(_01656_));
 sky130_fd_sc_hd__and2_1 _18282_ (.A(_01651_),
    .B(_01656_),
    .X(_01657_));
 sky130_fd_sc_hd__clkbuf_1 _18283_ (.A(_01657_),
    .X(_00506_));
 sky130_fd_sc_hd__mux2_1 _18284_ (.A0(net81),
    .A1(\wfg_core_top.cfg_subcycle_q[23] ),
    .S(_01646_),
    .X(_01658_));
 sky130_fd_sc_hd__and2_1 _18285_ (.A(_01651_),
    .B(_01658_),
    .X(_01659_));
 sky130_fd_sc_hd__clkbuf_1 _18286_ (.A(_01659_),
    .X(_00507_));
 sky130_fd_sc_hd__buf_6 _18287_ (.A(net66),
    .X(_01660_));
 sky130_fd_sc_hd__mux2_1 _18288_ (.A0(_01660_),
    .A1(\wfg_core_top.cfg_sync_q[0] ),
    .S(_01646_),
    .X(_01661_));
 sky130_fd_sc_hd__and2_1 _18289_ (.A(_01651_),
    .B(_01661_),
    .X(_01662_));
 sky130_fd_sc_hd__clkbuf_1 _18290_ (.A(_01662_),
    .X(_00508_));
 sky130_fd_sc_hd__buf_8 _18291_ (.A(net77),
    .X(_01663_));
 sky130_fd_sc_hd__mux2_1 _18292_ (.A0(_01663_),
    .A1(\wfg_core_top.cfg_sync_q[1] ),
    .S(_01646_),
    .X(_01664_));
 sky130_fd_sc_hd__and2_1 _18293_ (.A(_01651_),
    .B(_01664_),
    .X(_01665_));
 sky130_fd_sc_hd__clkbuf_1 _18294_ (.A(_01665_),
    .X(_00509_));
 sky130_fd_sc_hd__buf_6 _18295_ (.A(net88),
    .X(_01666_));
 sky130_fd_sc_hd__mux2_1 _18296_ (.A0(_01666_),
    .A1(\wfg_core_top.cfg_sync_q[2] ),
    .S(_01646_),
    .X(_01667_));
 sky130_fd_sc_hd__and2_1 _18297_ (.A(_01651_),
    .B(_01667_),
    .X(_01668_));
 sky130_fd_sc_hd__clkbuf_1 _18298_ (.A(_01668_),
    .X(_00510_));
 sky130_fd_sc_hd__clkbuf_8 _18299_ (.A(net91),
    .X(_01669_));
 sky130_fd_sc_hd__mux2_1 _18300_ (.A0(_01669_),
    .A1(\wfg_core_top.cfg_sync_q[3] ),
    .S(_01646_),
    .X(_01670_));
 sky130_fd_sc_hd__and2_1 _18301_ (.A(_01651_),
    .B(_01670_),
    .X(_01671_));
 sky130_fd_sc_hd__clkbuf_1 _18302_ (.A(_01671_),
    .X(_00511_));
 sky130_fd_sc_hd__buf_6 _18303_ (.A(net92),
    .X(_01672_));
 sky130_fd_sc_hd__mux2_1 _18304_ (.A0(_01672_),
    .A1(\wfg_core_top.cfg_sync_q[4] ),
    .S(_01616_),
    .X(_01673_));
 sky130_fd_sc_hd__and2_1 _18305_ (.A(_01651_),
    .B(_01673_),
    .X(_01674_));
 sky130_fd_sc_hd__clkbuf_1 _18306_ (.A(_01674_),
    .X(_00512_));
 sky130_fd_sc_hd__buf_6 _18307_ (.A(net93),
    .X(_01675_));
 sky130_fd_sc_hd__mux2_1 _18308_ (.A0(_01675_),
    .A1(\wfg_core_top.cfg_sync_q[5] ),
    .S(_01616_),
    .X(_01676_));
 sky130_fd_sc_hd__and2_1 _18309_ (.A(_01651_),
    .B(_01676_),
    .X(_01677_));
 sky130_fd_sc_hd__clkbuf_1 _18310_ (.A(_01677_),
    .X(_00513_));
 sky130_fd_sc_hd__buf_4 _18311_ (.A(_01599_),
    .X(_01678_));
 sky130_fd_sc_hd__buf_6 _18312_ (.A(net94),
    .X(_01679_));
 sky130_fd_sc_hd__mux2_1 _18313_ (.A0(_01679_),
    .A1(\wfg_core_top.cfg_sync_q[6] ),
    .S(_01616_),
    .X(_01680_));
 sky130_fd_sc_hd__and2_1 _18314_ (.A(_01678_),
    .B(_01680_),
    .X(_01681_));
 sky130_fd_sc_hd__clkbuf_1 _18315_ (.A(_01681_),
    .X(_00514_));
 sky130_fd_sc_hd__buf_6 _18316_ (.A(net95),
    .X(_01682_));
 sky130_fd_sc_hd__mux2_1 _18317_ (.A0(_01682_),
    .A1(\wfg_core_top.cfg_sync_q[7] ),
    .S(_01616_),
    .X(_01683_));
 sky130_fd_sc_hd__and2_1 _18318_ (.A(_01678_),
    .B(_01683_),
    .X(_01684_));
 sky130_fd_sc_hd__clkbuf_1 _18319_ (.A(_01684_),
    .X(_00515_));
 sky130_fd_sc_hd__buf_2 _18320_ (.A(_01588_),
    .X(_01685_));
 sky130_fd_sc_hd__clkbuf_4 _18321_ (.A(_01607_),
    .X(_01686_));
 sky130_fd_sc_hd__nand2_1 _18322_ (.A(_01442_),
    .B(_01608_),
    .Y(_01687_));
 sky130_fd_sc_hd__or2_2 _18323_ (.A(_01686_),
    .B(_01687_),
    .X(_01688_));
 sky130_fd_sc_hd__or2_2 _18324_ (.A(net55),
    .B(_01602_),
    .X(_01689_));
 sky130_fd_sc_hd__or2_4 _18325_ (.A(net58),
    .B(_01689_),
    .X(_01690_));
 sky130_fd_sc_hd__buf_4 _18326_ (.A(_01690_),
    .X(_01691_));
 sky130_fd_sc_hd__or4_1 _18327_ (.A(net66),
    .B(_01605_),
    .C(_01688_),
    .D(_01691_),
    .X(_01692_));
 sky130_fd_sc_hd__o31ai_1 _18328_ (.A1(_01605_),
    .A2(_01688_),
    .A3(_01691_),
    .B1(_01351_),
    .Y(_01693_));
 sky130_fd_sc_hd__and3_1 _18329_ (.A(_01685_),
    .B(_01692_),
    .C(_01693_),
    .X(_01694_));
 sky130_fd_sc_hd__clkbuf_1 _18330_ (.A(_01694_),
    .X(_00516_));
 sky130_fd_sc_hd__or2_2 _18331_ (.A(net59),
    .B(_01443_),
    .X(_01695_));
 sky130_fd_sc_hd__nor2_2 _18332_ (.A(_01695_),
    .B(_01686_),
    .Y(_01696_));
 sky130_fd_sc_hd__and2_1 _18333_ (.A(net65),
    .B(_01588_),
    .X(_01697_));
 sky130_fd_sc_hd__and3b_1 _18334_ (.A_N(\wfg_subcore_top.wbs_ack_o ),
    .B(_01696_),
    .C(_01697_),
    .X(_01698_));
 sky130_fd_sc_hd__clkbuf_1 _18335_ (.A(_01698_),
    .X(_00517_));
 sky130_fd_sc_hd__inv_2 _18336_ (.A(_01598_),
    .Y(_00074_));
 sky130_fd_sc_hd__inv_2 _18337_ (.A(_01598_),
    .Y(_00075_));
 sky130_fd_sc_hd__inv_2 _18338_ (.A(_01598_),
    .Y(_00076_));
 sky130_fd_sc_hd__inv_2 _18339_ (.A(_01598_),
    .Y(_00077_));
 sky130_fd_sc_hd__or3b_1 _18340_ (.A(\wfg_core_top.wbs_ack_o ),
    .B(_01688_),
    .C_N(_01697_),
    .X(_01699_));
 sky130_fd_sc_hd__clkinv_2 _18341_ (.A(_01699_),
    .Y(_00518_));
 sky130_fd_sc_hd__inv_2 _18342_ (.A(_01598_),
    .Y(_00078_));
 sky130_fd_sc_hd__inv_2 _18343_ (.A(_01598_),
    .Y(_00079_));
 sky130_fd_sc_hd__inv_2 _18344_ (.A(_01598_),
    .Y(_00080_));
 sky130_fd_sc_hd__buf_4 _18345_ (.A(_01597_),
    .X(_01700_));
 sky130_fd_sc_hd__inv_2 _18346_ (.A(_01700_),
    .Y(_00081_));
 sky130_fd_sc_hd__inv_2 _18347_ (.A(_01700_),
    .Y(_00082_));
 sky130_fd_sc_hd__inv_2 _18348_ (.A(_01700_),
    .Y(_00083_));
 sky130_fd_sc_hd__inv_2 _18349_ (.A(_01700_),
    .Y(_00084_));
 sky130_fd_sc_hd__inv_2 _18350_ (.A(_01700_),
    .Y(_00085_));
 sky130_fd_sc_hd__inv_2 _18351_ (.A(_01700_),
    .Y(_00086_));
 sky130_fd_sc_hd__inv_2 _18352_ (.A(_01700_),
    .Y(_00087_));
 sky130_fd_sc_hd__inv_2 _18353_ (.A(_01700_),
    .Y(_00088_));
 sky130_fd_sc_hd__inv_2 _18354_ (.A(_01700_),
    .Y(_00089_));
 sky130_fd_sc_hd__inv_2 _18355_ (.A(_01700_),
    .Y(_00090_));
 sky130_fd_sc_hd__buf_4 _18356_ (.A(_01597_),
    .X(_01701_));
 sky130_fd_sc_hd__inv_2 _18357_ (.A(_01701_),
    .Y(_00091_));
 sky130_fd_sc_hd__inv_2 _18358_ (.A(_01701_),
    .Y(_00092_));
 sky130_fd_sc_hd__inv_2 _18359_ (.A(_01701_),
    .Y(_00093_));
 sky130_fd_sc_hd__inv_2 _18360_ (.A(_01701_),
    .Y(_00094_));
 sky130_fd_sc_hd__inv_2 _18361_ (.A(_01701_),
    .Y(_00095_));
 sky130_fd_sc_hd__inv_2 _18362_ (.A(_01701_),
    .Y(_00096_));
 sky130_fd_sc_hd__inv_2 _18363_ (.A(_01701_),
    .Y(_00097_));
 sky130_fd_sc_hd__inv_2 _18364_ (.A(_01701_),
    .Y(_00098_));
 sky130_fd_sc_hd__inv_2 _18365_ (.A(_01701_),
    .Y(_00099_));
 sky130_fd_sc_hd__inv_2 _18366_ (.A(_01701_),
    .Y(_00100_));
 sky130_fd_sc_hd__buf_4 _18367_ (.A(_01597_),
    .X(_01702_));
 sky130_fd_sc_hd__inv_2 _18368_ (.A(_01702_),
    .Y(_00101_));
 sky130_fd_sc_hd__inv_2 _18369_ (.A(_01702_),
    .Y(_00102_));
 sky130_fd_sc_hd__inv_2 _18370_ (.A(_01702_),
    .Y(_00103_));
 sky130_fd_sc_hd__inv_2 _18371_ (.A(_01702_),
    .Y(_00104_));
 sky130_fd_sc_hd__inv_2 _18372_ (.A(_01702_),
    .Y(_00105_));
 sky130_fd_sc_hd__inv_2 _18373_ (.A(_01702_),
    .Y(_00106_));
 sky130_fd_sc_hd__inv_2 _18374_ (.A(_01702_),
    .Y(_00107_));
 sky130_fd_sc_hd__inv_2 _18375_ (.A(_01702_),
    .Y(_00108_));
 sky130_fd_sc_hd__inv_2 _18376_ (.A(_01702_),
    .Y(_00109_));
 sky130_fd_sc_hd__inv_2 _18377_ (.A(_01702_),
    .Y(_00110_));
 sky130_fd_sc_hd__buf_6 _18378_ (.A(_01597_),
    .X(_01703_));
 sky130_fd_sc_hd__inv_2 _18379_ (.A(_01703_),
    .Y(_00111_));
 sky130_fd_sc_hd__inv_2 _18380_ (.A(_01703_),
    .Y(_00112_));
 sky130_fd_sc_hd__inv_2 _18381_ (.A(_01703_),
    .Y(_00113_));
 sky130_fd_sc_hd__inv_2 _18382_ (.A(_01703_),
    .Y(_00114_));
 sky130_fd_sc_hd__inv_2 _18383_ (.A(_01703_),
    .Y(_00115_));
 sky130_fd_sc_hd__inv_2 _18384_ (.A(_01703_),
    .Y(_00116_));
 sky130_fd_sc_hd__inv_2 _18385_ (.A(_01703_),
    .Y(_00117_));
 sky130_fd_sc_hd__inv_2 _18386_ (.A(_01703_),
    .Y(_00118_));
 sky130_fd_sc_hd__inv_2 _18387_ (.A(_01703_),
    .Y(_00119_));
 sky130_fd_sc_hd__inv_2 _18388_ (.A(_01703_),
    .Y(_00120_));
 sky130_fd_sc_hd__buf_4 _18389_ (.A(_01597_),
    .X(_01704_));
 sky130_fd_sc_hd__inv_2 _18390_ (.A(_01704_),
    .Y(_00121_));
 sky130_fd_sc_hd__inv_2 _18391_ (.A(_01704_),
    .Y(_00122_));
 sky130_fd_sc_hd__inv_2 _18392_ (.A(_01704_),
    .Y(_00123_));
 sky130_fd_sc_hd__inv_2 _18393_ (.A(_01704_),
    .Y(_00124_));
 sky130_fd_sc_hd__and2b_1 _18394_ (.A_N(net100),
    .B(net65),
    .X(_01705_));
 sky130_fd_sc_hd__buf_4 _18395_ (.A(_01705_),
    .X(_01706_));
 sky130_fd_sc_hd__nand2_2 _18396_ (.A(_01696_),
    .B(_01706_),
    .Y(_01707_));
 sky130_fd_sc_hd__buf_2 _18397_ (.A(_01707_),
    .X(_01708_));
 sky130_fd_sc_hd__nor2_8 _18398_ (.A(net58),
    .B(_01689_),
    .Y(_01709_));
 sky130_fd_sc_hd__nor2_2 _18399_ (.A(_01695_),
    .B(_01709_),
    .Y(_01710_));
 sky130_fd_sc_hd__or3_1 _18400_ (.A(\wfg_subcore_top.cfg_sync_q[0] ),
    .B(_01695_),
    .C(_01709_),
    .X(_01711_));
 sky130_fd_sc_hd__or2_1 _18401_ (.A(_01695_),
    .B(_01686_),
    .X(_01712_));
 sky130_fd_sc_hd__or2b_2 _18402_ (.A(net100),
    .B_N(net65),
    .X(_01713_));
 sky130_fd_sc_hd__nor2_2 _18403_ (.A(_01712_),
    .B(_01713_),
    .Y(_01714_));
 sky130_fd_sc_hd__o211a_1 _18404_ (.A1(\wfg_subcore_top.active_o ),
    .A2(_01710_),
    .B1(_01711_),
    .C1(_01714_),
    .X(_01715_));
 sky130_fd_sc_hd__a21oi_1 _18405_ (.A1(\wfg_subcore_top.wbs_dat_o[0] ),
    .A2(_01708_),
    .B1(_01715_),
    .Y(_01716_));
 sky130_fd_sc_hd__nor2_1 _18406_ (.A(_01591_),
    .B(_01716_),
    .Y(_00565_));
 sky130_fd_sc_hd__buf_2 _18407_ (.A(_01714_),
    .X(_01717_));
 sky130_fd_sc_hd__buf_2 _18408_ (.A(_01710_),
    .X(_01718_));
 sky130_fd_sc_hd__a21o_1 _18409_ (.A1(\wfg_subcore_top.cfg_sync_q[1] ),
    .A2(_01718_),
    .B1(_01708_),
    .X(_01719_));
 sky130_fd_sc_hd__o211a_1 _18410_ (.A1(\wfg_subcore_top.wbs_dat_o[1] ),
    .A2(_01717_),
    .B1(_01719_),
    .C1(_00040_),
    .X(_00566_));
 sky130_fd_sc_hd__a21o_1 _18411_ (.A1(\wfg_subcore_top.cfg_sync_q[2] ),
    .A2(_01718_),
    .B1(_01708_),
    .X(_01720_));
 sky130_fd_sc_hd__o211a_1 _18412_ (.A1(\wfg_subcore_top.wbs_dat_o[2] ),
    .A2(_01717_),
    .B1(_01720_),
    .C1(_00040_),
    .X(_00567_));
 sky130_fd_sc_hd__a21o_1 _18413_ (.A1(\wfg_subcore_top.cfg_sync_q[3] ),
    .A2(_01718_),
    .B1(_01708_),
    .X(_01721_));
 sky130_fd_sc_hd__o211a_1 _18414_ (.A1(\wfg_subcore_top.wbs_dat_o[3] ),
    .A2(_01717_),
    .B1(_01721_),
    .C1(_00040_),
    .X(_00568_));
 sky130_fd_sc_hd__a21o_1 _18415_ (.A1(\wfg_subcore_top.cfg_sync_q[4] ),
    .A2(_01718_),
    .B1(_01708_),
    .X(_01722_));
 sky130_fd_sc_hd__o211a_1 _18416_ (.A1(\wfg_subcore_top.wbs_dat_o[4] ),
    .A2(_01717_),
    .B1(_01722_),
    .C1(_00040_),
    .X(_00569_));
 sky130_fd_sc_hd__a21o_1 _18417_ (.A1(\wfg_subcore_top.cfg_sync_q[5] ),
    .A2(_01718_),
    .B1(_01708_),
    .X(_01723_));
 sky130_fd_sc_hd__o211a_1 _18418_ (.A1(\wfg_subcore_top.wbs_dat_o[5] ),
    .A2(_01717_),
    .B1(_01723_),
    .C1(_00040_),
    .X(_00570_));
 sky130_fd_sc_hd__a21o_1 _18419_ (.A1(\wfg_subcore_top.cfg_sync_q[6] ),
    .A2(_01718_),
    .B1(_01708_),
    .X(_01724_));
 sky130_fd_sc_hd__o211a_1 _18420_ (.A1(\wfg_subcore_top.wbs_dat_o[6] ),
    .A2(_01717_),
    .B1(_01724_),
    .C1(_00040_),
    .X(_00571_));
 sky130_fd_sc_hd__a21o_1 _18421_ (.A1(\wfg_subcore_top.cfg_sync_q[7] ),
    .A2(_01718_),
    .B1(_01708_),
    .X(_01725_));
 sky130_fd_sc_hd__o211a_1 _18422_ (.A1(\wfg_subcore_top.wbs_dat_o[7] ),
    .A2(_01717_),
    .B1(_01725_),
    .C1(_00040_),
    .X(_00572_));
 sky130_fd_sc_hd__a21o_1 _18423_ (.A1(\wfg_subcore_top.cfg_subcycle_q[8] ),
    .A2(_01718_),
    .B1(_01708_),
    .X(_01726_));
 sky130_fd_sc_hd__o211a_1 _18424_ (.A1(\wfg_subcore_top.wbs_dat_o[8] ),
    .A2(_01717_),
    .B1(_01726_),
    .C1(_00040_),
    .X(_00573_));
 sky130_fd_sc_hd__a21o_1 _18425_ (.A1(\wfg_subcore_top.cfg_subcycle_q[9] ),
    .A2(_01718_),
    .B1(_01708_),
    .X(_01727_));
 sky130_fd_sc_hd__o211a_1 _18426_ (.A1(\wfg_subcore_top.wbs_dat_o[9] ),
    .A2(_01717_),
    .B1(_01727_),
    .C1(_00040_),
    .X(_00574_));
 sky130_fd_sc_hd__buf_2 _18427_ (.A(_01707_),
    .X(_01728_));
 sky130_fd_sc_hd__a21o_1 _18428_ (.A1(\wfg_subcore_top.cfg_subcycle_q[10] ),
    .A2(_01718_),
    .B1(_01728_),
    .X(_01729_));
 sky130_fd_sc_hd__buf_6 _18429_ (.A(_01588_),
    .X(_01730_));
 sky130_fd_sc_hd__buf_2 _18430_ (.A(_01730_),
    .X(_01731_));
 sky130_fd_sc_hd__o211a_1 _18431_ (.A1(\wfg_subcore_top.wbs_dat_o[10] ),
    .A2(_01717_),
    .B1(_01729_),
    .C1(_01731_),
    .X(_00575_));
 sky130_fd_sc_hd__buf_2 _18432_ (.A(_01714_),
    .X(_01732_));
 sky130_fd_sc_hd__buf_2 _18433_ (.A(_01710_),
    .X(_01733_));
 sky130_fd_sc_hd__a21o_1 _18434_ (.A1(\wfg_subcore_top.cfg_subcycle_q[11] ),
    .A2(_01733_),
    .B1(_01728_),
    .X(_01734_));
 sky130_fd_sc_hd__o211a_1 _18435_ (.A1(\wfg_subcore_top.wbs_dat_o[11] ),
    .A2(_01732_),
    .B1(_01734_),
    .C1(_01731_),
    .X(_00576_));
 sky130_fd_sc_hd__a21o_1 _18436_ (.A1(\wfg_subcore_top.cfg_subcycle_q[12] ),
    .A2(_01733_),
    .B1(_01728_),
    .X(_01735_));
 sky130_fd_sc_hd__o211a_1 _18437_ (.A1(\wfg_subcore_top.wbs_dat_o[12] ),
    .A2(_01732_),
    .B1(_01735_),
    .C1(_01731_),
    .X(_00577_));
 sky130_fd_sc_hd__a21o_1 _18438_ (.A1(\wfg_subcore_top.cfg_subcycle_q[13] ),
    .A2(_01733_),
    .B1(_01728_),
    .X(_01736_));
 sky130_fd_sc_hd__o211a_1 _18439_ (.A1(\wfg_subcore_top.wbs_dat_o[13] ),
    .A2(_01732_),
    .B1(_01736_),
    .C1(_01731_),
    .X(_00578_));
 sky130_fd_sc_hd__a21o_1 _18440_ (.A1(\wfg_subcore_top.cfg_subcycle_q[14] ),
    .A2(_01733_),
    .B1(_01728_),
    .X(_01737_));
 sky130_fd_sc_hd__o211a_1 _18441_ (.A1(\wfg_subcore_top.wbs_dat_o[14] ),
    .A2(_01732_),
    .B1(_01737_),
    .C1(_01731_),
    .X(_00579_));
 sky130_fd_sc_hd__a21o_1 _18442_ (.A1(\wfg_subcore_top.cfg_subcycle_q[15] ),
    .A2(_01733_),
    .B1(_01728_),
    .X(_01738_));
 sky130_fd_sc_hd__o211a_1 _18443_ (.A1(\wfg_subcore_top.wbs_dat_o[15] ),
    .A2(_01732_),
    .B1(_01738_),
    .C1(_01731_),
    .X(_00580_));
 sky130_fd_sc_hd__a21o_1 _18444_ (.A1(\wfg_subcore_top.cfg_subcycle_q[16] ),
    .A2(_01733_),
    .B1(_01728_),
    .X(_01739_));
 sky130_fd_sc_hd__o211a_1 _18445_ (.A1(\wfg_subcore_top.wbs_dat_o[16] ),
    .A2(_01732_),
    .B1(_01739_),
    .C1(_01731_),
    .X(_00581_));
 sky130_fd_sc_hd__a21o_1 _18446_ (.A1(\wfg_subcore_top.cfg_subcycle_q[17] ),
    .A2(_01733_),
    .B1(_01728_),
    .X(_01740_));
 sky130_fd_sc_hd__o211a_1 _18447_ (.A1(\wfg_subcore_top.wbs_dat_o[17] ),
    .A2(_01732_),
    .B1(_01740_),
    .C1(_01731_),
    .X(_00582_));
 sky130_fd_sc_hd__a21o_1 _18448_ (.A1(\wfg_subcore_top.cfg_subcycle_q[18] ),
    .A2(_01733_),
    .B1(_01728_),
    .X(_01741_));
 sky130_fd_sc_hd__o211a_1 _18449_ (.A1(\wfg_subcore_top.wbs_dat_o[18] ),
    .A2(_01732_),
    .B1(_01741_),
    .C1(_01731_),
    .X(_00583_));
 sky130_fd_sc_hd__a21o_1 _18450_ (.A1(\wfg_subcore_top.cfg_subcycle_q[19] ),
    .A2(_01733_),
    .B1(_01728_),
    .X(_01742_));
 sky130_fd_sc_hd__o211a_1 _18451_ (.A1(\wfg_subcore_top.wbs_dat_o[19] ),
    .A2(_01732_),
    .B1(_01742_),
    .C1(_01731_),
    .X(_00584_));
 sky130_fd_sc_hd__a21o_1 _18452_ (.A1(\wfg_subcore_top.cfg_subcycle_q[20] ),
    .A2(_01733_),
    .B1(_01707_),
    .X(_01743_));
 sky130_fd_sc_hd__clkbuf_4 _18453_ (.A(_01730_),
    .X(_01744_));
 sky130_fd_sc_hd__o211a_1 _18454_ (.A1(\wfg_subcore_top.wbs_dat_o[20] ),
    .A2(_01732_),
    .B1(_01743_),
    .C1(_01744_),
    .X(_00585_));
 sky130_fd_sc_hd__a21o_1 _18455_ (.A1(\wfg_subcore_top.cfg_subcycle_q[21] ),
    .A2(_01710_),
    .B1(_01707_),
    .X(_01745_));
 sky130_fd_sc_hd__o211a_1 _18456_ (.A1(\wfg_subcore_top.wbs_dat_o[21] ),
    .A2(_01714_),
    .B1(_01745_),
    .C1(_01744_),
    .X(_00586_));
 sky130_fd_sc_hd__a21o_1 _18457_ (.A1(\wfg_subcore_top.cfg_subcycle_q[22] ),
    .A2(_01710_),
    .B1(_01707_),
    .X(_01746_));
 sky130_fd_sc_hd__o211a_1 _18458_ (.A1(\wfg_subcore_top.wbs_dat_o[22] ),
    .A2(_01714_),
    .B1(_01746_),
    .C1(_01744_),
    .X(_00587_));
 sky130_fd_sc_hd__a21o_1 _18459_ (.A1(\wfg_subcore_top.cfg_subcycle_q[23] ),
    .A2(_01710_),
    .B1(_01707_),
    .X(_01747_));
 sky130_fd_sc_hd__o211a_1 _18460_ (.A1(\wfg_subcore_top.wbs_dat_o[23] ),
    .A2(_01714_),
    .B1(_01747_),
    .C1(_01744_),
    .X(_00588_));
 sky130_fd_sc_hd__inv_2 _18461_ (.A(_01704_),
    .Y(_00125_));
 sky130_fd_sc_hd__inv_2 _18462_ (.A(_01704_),
    .Y(_00126_));
 sky130_fd_sc_hd__inv_2 _18463_ (.A(_01704_),
    .Y(_00127_));
 sky130_fd_sc_hd__inv_2 _18464_ (.A(_01704_),
    .Y(_00128_));
 sky130_fd_sc_hd__inv_2 _18465_ (.A(_01704_),
    .Y(_00129_));
 sky130_fd_sc_hd__inv_2 _18466_ (.A(_01704_),
    .Y(_00130_));
 sky130_fd_sc_hd__buf_4 _18467_ (.A(_01597_),
    .X(_01748_));
 sky130_fd_sc_hd__inv_2 _18468_ (.A(_01748_),
    .Y(_00131_));
 sky130_fd_sc_hd__inv_2 _18469_ (.A(_01748_),
    .Y(_00132_));
 sky130_fd_sc_hd__inv_2 _18470_ (.A(_01748_),
    .Y(_00133_));
 sky130_fd_sc_hd__inv_2 _18471_ (.A(_01748_),
    .Y(_00134_));
 sky130_fd_sc_hd__inv_2 _18472_ (.A(_01748_),
    .Y(_00135_));
 sky130_fd_sc_hd__inv_2 _18473_ (.A(_01748_),
    .Y(_00136_));
 sky130_fd_sc_hd__inv_2 _18474_ (.A(_01748_),
    .Y(_00137_));
 sky130_fd_sc_hd__inv_2 _18475_ (.A(_01748_),
    .Y(_00138_));
 sky130_fd_sc_hd__inv_2 _18476_ (.A(_01748_),
    .Y(_00139_));
 sky130_fd_sc_hd__inv_2 _18477_ (.A(_01748_),
    .Y(_00140_));
 sky130_fd_sc_hd__buf_8 _18478_ (.A(_01597_),
    .X(_01749_));
 sky130_fd_sc_hd__inv_2 _18479_ (.A(_01749_),
    .Y(_00141_));
 sky130_fd_sc_hd__inv_2 _18480_ (.A(_01749_),
    .Y(_00142_));
 sky130_fd_sc_hd__clkinv_2 _18481_ (.A(_01607_),
    .Y(_01750_));
 sky130_fd_sc_hd__and3_2 _18482_ (.A(_01433_),
    .B(_01750_),
    .C(_01706_),
    .X(_01751_));
 sky130_fd_sc_hd__buf_4 _18483_ (.A(_01751_),
    .X(_01752_));
 sky130_fd_sc_hd__buf_4 _18484_ (.A(_01752_),
    .X(_01753_));
 sky130_fd_sc_hd__or2_4 _18485_ (.A(_01431_),
    .B(_01428_),
    .X(_01754_));
 sky130_fd_sc_hd__nor2_4 _18486_ (.A(net33),
    .B(net44),
    .Y(_01755_));
 sky130_fd_sc_hd__nand3_4 _18487_ (.A(net55),
    .B(net58),
    .C(_01755_),
    .Y(_01756_));
 sky130_fd_sc_hd__nor2_4 _18488_ (.A(_01754_),
    .B(_01756_),
    .Y(_01757_));
 sky130_fd_sc_hd__buf_4 _18489_ (.A(_01757_),
    .X(_01758_));
 sky130_fd_sc_hd__clkbuf_4 _18490_ (.A(_01758_),
    .X(_01759_));
 sky130_fd_sc_hd__a21oi_4 _18491_ (.A1(_01755_),
    .A2(_01603_),
    .B1(_01754_),
    .Y(_01760_));
 sky130_fd_sc_hd__nor2_2 _18492_ (.A(net55),
    .B(_01602_),
    .Y(_01761_));
 sky130_fd_sc_hd__nand2_2 _18493_ (.A(net58),
    .B(_01761_),
    .Y(_01762_));
 sky130_fd_sc_hd__buf_6 _18494_ (.A(_01762_),
    .X(_01763_));
 sky130_fd_sc_hd__nor2_4 _18495_ (.A(_01754_),
    .B(_01763_),
    .Y(_01764_));
 sky130_fd_sc_hd__a22o_1 _18496_ (.A1(\wfg_drive_pat_top.cfg_begin_q[0] ),
    .A2(_01760_),
    .B1(_01764_),
    .B2(\wfg_drive_pat_top.patsel0_low_q[0] ),
    .X(_01765_));
 sky130_fd_sc_hd__nand2_4 _18497_ (.A(_01433_),
    .B(_01690_),
    .Y(_01766_));
 sky130_fd_sc_hd__buf_4 _18498_ (.A(_01766_),
    .X(_01767_));
 sky130_fd_sc_hd__buf_4 _18499_ (.A(_01767_),
    .X(_01768_));
 sky130_fd_sc_hd__or3_4 _18500_ (.A(_01754_),
    .B(_01686_),
    .C(_01713_),
    .X(_01769_));
 sky130_fd_sc_hd__buf_4 _18501_ (.A(_01769_),
    .X(_01770_));
 sky130_fd_sc_hd__a21o_1 _18502_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[0].drv.ctrl_en_q_i ),
    .A2(_01768_),
    .B1(_01770_),
    .X(_01771_));
 sky130_fd_sc_hd__a211o_1 _18503_ (.A1(\wfg_drive_pat_top.patsel1_high_q[0] ),
    .A2(_01759_),
    .B1(_01765_),
    .C1(_01771_),
    .X(_01772_));
 sky130_fd_sc_hd__o211a_1 _18504_ (.A1(\wfg_drive_pat_top.wbs_dat_o[0] ),
    .A2(_01753_),
    .B1(_01772_),
    .C1(_01744_),
    .X(_00607_));
 sky130_fd_sc_hd__buf_2 _18505_ (.A(_01751_),
    .X(_01773_));
 sky130_fd_sc_hd__clkbuf_4 _18506_ (.A(_01766_),
    .X(_01774_));
 sky130_fd_sc_hd__a21o_1 _18507_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[1].drv.ctrl_en_q_i ),
    .A2(_01774_),
    .B1(_01770_),
    .X(_01775_));
 sky130_fd_sc_hd__clkbuf_4 _18508_ (.A(_01760_),
    .X(_01776_));
 sky130_fd_sc_hd__buf_4 _18509_ (.A(_01764_),
    .X(_01777_));
 sky130_fd_sc_hd__a22o_1 _18510_ (.A1(\wfg_drive_pat_top.cfg_begin_q[1] ),
    .A2(_01776_),
    .B1(_01777_),
    .B2(\wfg_drive_pat_top.patsel0_low_q[1] ),
    .X(_01778_));
 sky130_fd_sc_hd__a211o_1 _18511_ (.A1(\wfg_drive_pat_top.patsel1_high_q[1] ),
    .A2(_01759_),
    .B1(_01775_),
    .C1(_01778_),
    .X(_01779_));
 sky130_fd_sc_hd__o211a_1 _18512_ (.A1(\wfg_drive_pat_top.wbs_dat_o[1] ),
    .A2(_01773_),
    .B1(_01779_),
    .C1(_01744_),
    .X(_00608_));
 sky130_fd_sc_hd__or2_1 _18513_ (.A(\wfg_drive_pat_top.wbs_dat_o[2] ),
    .B(_01751_),
    .X(_01780_));
 sky130_fd_sc_hd__clkbuf_4 _18514_ (.A(_01764_),
    .X(_01781_));
 sky130_fd_sc_hd__a221o_1 _18515_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[2].drv.ctrl_en_q_i ),
    .A2(_01766_),
    .B1(_01757_),
    .B2(\wfg_drive_pat_top.patsel1_high_q[2] ),
    .C1(_01769_),
    .X(_01782_));
 sky130_fd_sc_hd__a221o_2 _18516_ (.A1(\wfg_drive_pat_top.cfg_begin_q[2] ),
    .A2(_01760_),
    .B1(_01781_),
    .B2(\wfg_drive_pat_top.patsel0_low_q[2] ),
    .C1(_01782_),
    .X(_01783_));
 sky130_fd_sc_hd__and3_1 _18517_ (.A(_01685_),
    .B(_01780_),
    .C(_01783_),
    .X(_01784_));
 sky130_fd_sc_hd__clkbuf_1 _18518_ (.A(_01784_),
    .X(_00609_));
 sky130_fd_sc_hd__a21o_1 _18519_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[3].drv.ctrl_en_q_i ),
    .A2(_01774_),
    .B1(_01770_),
    .X(_01785_));
 sky130_fd_sc_hd__a22o_1 _18520_ (.A1(\wfg_drive_pat_top.cfg_begin_q[3] ),
    .A2(_01776_),
    .B1(_01777_),
    .B2(\wfg_drive_pat_top.patsel0_low_q[3] ),
    .X(_01786_));
 sky130_fd_sc_hd__a211o_1 _18521_ (.A1(\wfg_drive_pat_top.patsel1_high_q[3] ),
    .A2(_01759_),
    .B1(_01785_),
    .C1(_01786_),
    .X(_01787_));
 sky130_fd_sc_hd__o211a_1 _18522_ (.A1(\wfg_drive_pat_top.wbs_dat_o[3] ),
    .A2(_01773_),
    .B1(_01787_),
    .C1(_01744_),
    .X(_00610_));
 sky130_fd_sc_hd__a21o_1 _18523_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[4].drv.ctrl_en_q_i ),
    .A2(_01774_),
    .B1(_01770_),
    .X(_01788_));
 sky130_fd_sc_hd__a22o_1 _18524_ (.A1(\wfg_drive_pat_top.cfg_begin_q[4] ),
    .A2(_01776_),
    .B1(_01777_),
    .B2(\wfg_drive_pat_top.patsel0_low_q[4] ),
    .X(_01789_));
 sky130_fd_sc_hd__a211o_1 _18525_ (.A1(\wfg_drive_pat_top.patsel1_high_q[4] ),
    .A2(_01759_),
    .B1(_01788_),
    .C1(_01789_),
    .X(_01790_));
 sky130_fd_sc_hd__o211a_1 _18526_ (.A1(\wfg_drive_pat_top.wbs_dat_o[4] ),
    .A2(_01773_),
    .B1(_01790_),
    .C1(_01744_),
    .X(_00611_));
 sky130_fd_sc_hd__or2_1 _18527_ (.A(\wfg_drive_pat_top.wbs_dat_o[5] ),
    .B(_01751_),
    .X(_01791_));
 sky130_fd_sc_hd__a221o_1 _18528_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[5].drv.ctrl_en_q_i ),
    .A2(_01766_),
    .B1(_01757_),
    .B2(\wfg_drive_pat_top.patsel1_high_q[5] ),
    .C1(_01769_),
    .X(_01792_));
 sky130_fd_sc_hd__a221o_1 _18529_ (.A1(\wfg_drive_pat_top.cfg_begin_q[5] ),
    .A2(_01760_),
    .B1(_01781_),
    .B2(\wfg_drive_pat_top.patsel0_low_q[5] ),
    .C1(_01792_),
    .X(_01793_));
 sky130_fd_sc_hd__and3_1 _18530_ (.A(_01685_),
    .B(_01791_),
    .C(_01793_),
    .X(_01794_));
 sky130_fd_sc_hd__clkbuf_1 _18531_ (.A(_01794_),
    .X(_00612_));
 sky130_fd_sc_hd__a21o_1 _18532_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[6].drv.ctrl_en_q_i ),
    .A2(_01774_),
    .B1(_01770_),
    .X(_01795_));
 sky130_fd_sc_hd__a22o_1 _18533_ (.A1(\wfg_drive_pat_top.cfg_begin_q[6] ),
    .A2(_01776_),
    .B1(_01777_),
    .B2(\wfg_drive_pat_top.patsel0_low_q[6] ),
    .X(_01796_));
 sky130_fd_sc_hd__a211o_1 _18534_ (.A1(\wfg_drive_pat_top.patsel1_high_q[6] ),
    .A2(_01759_),
    .B1(_01795_),
    .C1(_01796_),
    .X(_01797_));
 sky130_fd_sc_hd__o211a_1 _18535_ (.A1(\wfg_drive_pat_top.wbs_dat_o[6] ),
    .A2(_01773_),
    .B1(_01797_),
    .C1(_01744_),
    .X(_00613_));
 sky130_fd_sc_hd__clkbuf_4 _18536_ (.A(_01769_),
    .X(_01798_));
 sky130_fd_sc_hd__a21o_1 _18537_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[7].drv.ctrl_en_q_i ),
    .A2(_01774_),
    .B1(_01798_),
    .X(_01799_));
 sky130_fd_sc_hd__a22o_1 _18538_ (.A1(\wfg_drive_pat_top.cfg_begin_q[7] ),
    .A2(_01776_),
    .B1(_01777_),
    .B2(\wfg_drive_pat_top.patsel0_low_q[7] ),
    .X(_01800_));
 sky130_fd_sc_hd__a211o_1 _18539_ (.A1(\wfg_drive_pat_top.patsel1_high_q[7] ),
    .A2(_01759_),
    .B1(_01799_),
    .C1(_01800_),
    .X(_01801_));
 sky130_fd_sc_hd__o211a_1 _18540_ (.A1(\wfg_drive_pat_top.wbs_dat_o[7] ),
    .A2(_01773_),
    .B1(_01801_),
    .C1(_01744_),
    .X(_00614_));
 sky130_fd_sc_hd__a21o_1 _18541_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[8].drv.ctrl_en_q_i ),
    .A2(_01774_),
    .B1(_01798_),
    .X(_01802_));
 sky130_fd_sc_hd__a22o_1 _18542_ (.A1(\wfg_drive_pat_top.cfg_end_q[8] ),
    .A2(_01776_),
    .B1(_01781_),
    .B2(\wfg_drive_pat_top.patsel0_low_q[8] ),
    .X(_01803_));
 sky130_fd_sc_hd__a211o_1 _18543_ (.A1(\wfg_drive_pat_top.patsel1_high_q[8] ),
    .A2(_01759_),
    .B1(_01802_),
    .C1(_01803_),
    .X(_01804_));
 sky130_fd_sc_hd__clkbuf_4 _18544_ (.A(_01730_),
    .X(_01805_));
 sky130_fd_sc_hd__o211a_1 _18545_ (.A1(\wfg_drive_pat_top.wbs_dat_o[8] ),
    .A2(_01773_),
    .B1(_01804_),
    .C1(_01805_),
    .X(_00615_));
 sky130_fd_sc_hd__a21o_1 _18546_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[9].drv.ctrl_en_q_i ),
    .A2(_01774_),
    .B1(_01798_),
    .X(_01806_));
 sky130_fd_sc_hd__a22o_1 _18547_ (.A1(\wfg_drive_pat_top.cfg_end_q[9] ),
    .A2(_01776_),
    .B1(_01781_),
    .B2(\wfg_drive_pat_top.patsel0_low_q[9] ),
    .X(_01807_));
 sky130_fd_sc_hd__a211o_1 _18548_ (.A1(\wfg_drive_pat_top.patsel1_high_q[9] ),
    .A2(_01759_),
    .B1(_01806_),
    .C1(_01807_),
    .X(_01808_));
 sky130_fd_sc_hd__o211a_1 _18549_ (.A1(\wfg_drive_pat_top.wbs_dat_o[9] ),
    .A2(_01773_),
    .B1(_01808_),
    .C1(_01805_),
    .X(_00616_));
 sky130_fd_sc_hd__a21o_1 _18550_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[10].drv.ctrl_en_q_i ),
    .A2(_01774_),
    .B1(_01798_),
    .X(_01809_));
 sky130_fd_sc_hd__a22o_1 _18551_ (.A1(\wfg_drive_pat_top.cfg_end_q[10] ),
    .A2(_01776_),
    .B1(_01781_),
    .B2(\wfg_drive_pat_top.patsel0_low_q[10] ),
    .X(_01810_));
 sky130_fd_sc_hd__a211o_1 _18552_ (.A1(\wfg_drive_pat_top.patsel1_high_q[10] ),
    .A2(_01759_),
    .B1(_01809_),
    .C1(_01810_),
    .X(_01811_));
 sky130_fd_sc_hd__o211a_1 _18553_ (.A1(\wfg_drive_pat_top.wbs_dat_o[10] ),
    .A2(_01773_),
    .B1(_01811_),
    .C1(_01805_),
    .X(_00617_));
 sky130_fd_sc_hd__a21o_1 _18554_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[11].drv.ctrl_en_q_i ),
    .A2(_01774_),
    .B1(_01798_),
    .X(_01812_));
 sky130_fd_sc_hd__a22o_1 _18555_ (.A1(\wfg_drive_pat_top.cfg_end_q[11] ),
    .A2(_01776_),
    .B1(_01781_),
    .B2(\wfg_drive_pat_top.patsel0_low_q[11] ),
    .X(_01813_));
 sky130_fd_sc_hd__a211o_1 _18556_ (.A1(\wfg_drive_pat_top.patsel1_high_q[11] ),
    .A2(_01759_),
    .B1(_01812_),
    .C1(_01813_),
    .X(_01814_));
 sky130_fd_sc_hd__o211a_1 _18557_ (.A1(\wfg_drive_pat_top.wbs_dat_o[11] ),
    .A2(_01773_),
    .B1(_01814_),
    .C1(_01805_),
    .X(_00618_));
 sky130_fd_sc_hd__clkbuf_4 _18558_ (.A(_01757_),
    .X(_01815_));
 sky130_fd_sc_hd__a21o_1 _18559_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[12].drv.ctrl_en_q_i ),
    .A2(_01774_),
    .B1(_01798_),
    .X(_01816_));
 sky130_fd_sc_hd__a22o_1 _18560_ (.A1(\wfg_drive_pat_top.cfg_end_q[12] ),
    .A2(_01776_),
    .B1(_01781_),
    .B2(\wfg_drive_pat_top.patsel0_low_q[12] ),
    .X(_01817_));
 sky130_fd_sc_hd__a211o_1 _18561_ (.A1(\wfg_drive_pat_top.patsel1_high_q[12] ),
    .A2(_01815_),
    .B1(_01816_),
    .C1(_01817_),
    .X(_01818_));
 sky130_fd_sc_hd__o211a_1 _18562_ (.A1(\wfg_drive_pat_top.wbs_dat_o[12] ),
    .A2(_01773_),
    .B1(_01818_),
    .C1(_01805_),
    .X(_00619_));
 sky130_fd_sc_hd__a21o_1 _18563_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[13].drv.ctrl_en_q_i ),
    .A2(_01767_),
    .B1(_01798_),
    .X(_01819_));
 sky130_fd_sc_hd__a22o_1 _18564_ (.A1(\wfg_drive_pat_top.cfg_end_q[13] ),
    .A2(_01760_),
    .B1(_01781_),
    .B2(\wfg_drive_pat_top.patsel0_low_q[13] ),
    .X(_01820_));
 sky130_fd_sc_hd__a211o_1 _18565_ (.A1(\wfg_drive_pat_top.patsel1_high_q[13] ),
    .A2(_01815_),
    .B1(_01819_),
    .C1(_01820_),
    .X(_01821_));
 sky130_fd_sc_hd__o211a_1 _18566_ (.A1(\wfg_drive_pat_top.wbs_dat_o[13] ),
    .A2(_01752_),
    .B1(_01821_),
    .C1(_01805_),
    .X(_00620_));
 sky130_fd_sc_hd__a21o_1 _18567_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[14].drv.ctrl_en_q_i ),
    .A2(_01767_),
    .B1(_01798_),
    .X(_01822_));
 sky130_fd_sc_hd__a22o_1 _18568_ (.A1(\wfg_drive_pat_top.cfg_end_q[14] ),
    .A2(_01760_),
    .B1(_01781_),
    .B2(\wfg_drive_pat_top.patsel0_low_q[14] ),
    .X(_01823_));
 sky130_fd_sc_hd__a211o_1 _18569_ (.A1(\wfg_drive_pat_top.patsel1_high_q[14] ),
    .A2(_01815_),
    .B1(_01822_),
    .C1(_01823_),
    .X(_01824_));
 sky130_fd_sc_hd__o211a_1 _18570_ (.A1(\wfg_drive_pat_top.wbs_dat_o[14] ),
    .A2(_01752_),
    .B1(_01824_),
    .C1(_01805_),
    .X(_00621_));
 sky130_fd_sc_hd__or2_1 _18571_ (.A(\wfg_drive_pat_top.wbs_dat_o[15] ),
    .B(_01751_),
    .X(_01825_));
 sky130_fd_sc_hd__a221o_1 _18572_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[15].drv.ctrl_en_q_i ),
    .A2(_01766_),
    .B1(_01757_),
    .B2(\wfg_drive_pat_top.patsel1_high_q[15] ),
    .C1(_01769_),
    .X(_01826_));
 sky130_fd_sc_hd__a221o_2 _18573_ (.A1(\wfg_drive_pat_top.cfg_end_q[15] ),
    .A2(_01760_),
    .B1(_01764_),
    .B2(\wfg_drive_pat_top.patsel0_low_q[15] ),
    .C1(_01826_),
    .X(_01827_));
 sky130_fd_sc_hd__and3_1 _18574_ (.A(_01685_),
    .B(_01825_),
    .C(_01827_),
    .X(_01828_));
 sky130_fd_sc_hd__clkbuf_1 _18575_ (.A(_01828_),
    .X(_00622_));
 sky130_fd_sc_hd__a21o_1 _18576_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[16].drv.ctrl_en_q_i ),
    .A2(_01767_),
    .B1(_01798_),
    .X(_01829_));
 sky130_fd_sc_hd__a22o_1 _18577_ (.A1(_09782_),
    .A2(_01760_),
    .B1(_01781_),
    .B2(\wfg_drive_pat_top.patsel0_low_q[16] ),
    .X(_01830_));
 sky130_fd_sc_hd__a211o_1 _18578_ (.A1(\wfg_drive_pat_top.patsel1_high_q[16] ),
    .A2(_01815_),
    .B1(_01829_),
    .C1(_01830_),
    .X(_01831_));
 sky130_fd_sc_hd__o211a_1 _18579_ (.A1(\wfg_drive_pat_top.wbs_dat_o[16] ),
    .A2(_01752_),
    .B1(_01831_),
    .C1(_01805_),
    .X(_00623_));
 sky130_fd_sc_hd__nand2_1 _18580_ (.A(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[17].drv.ctrl_en_q_i ),
    .B(_01768_),
    .Y(_01832_));
 sky130_fd_sc_hd__nand2_1 _18581_ (.A(\wfg_drive_pat_top.patsel1_high_q[17] ),
    .B(_01815_),
    .Y(_01833_));
 sky130_fd_sc_hd__clkbuf_4 _18582_ (.A(_01764_),
    .X(_01834_));
 sky130_fd_sc_hd__clkbuf_4 _18583_ (.A(_01798_),
    .X(_01835_));
 sky130_fd_sc_hd__a21oi_1 _18584_ (.A1(\wfg_drive_pat_top.patsel0_low_q[17] ),
    .A2(_01834_),
    .B1(_01835_),
    .Y(_01836_));
 sky130_fd_sc_hd__buf_8 _18585_ (.A(net98),
    .X(_01837_));
 sky130_fd_sc_hd__a31o_1 _18586_ (.A1(_01832_),
    .A2(_01833_),
    .A3(_01836_),
    .B1(_01837_),
    .X(_01838_));
 sky130_fd_sc_hd__o21ba_1 _18587_ (.A1(\wfg_drive_pat_top.wbs_dat_o[17] ),
    .A2(_01753_),
    .B1_N(_01838_),
    .X(_00624_));
 sky130_fd_sc_hd__nand2_1 _18588_ (.A(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[18].drv.ctrl_en_q_i ),
    .B(_01768_),
    .Y(_01839_));
 sky130_fd_sc_hd__nand2_1 _18589_ (.A(\wfg_drive_pat_top.patsel1_high_q[18] ),
    .B(_01815_),
    .Y(_01840_));
 sky130_fd_sc_hd__a21oi_1 _18590_ (.A1(\wfg_drive_pat_top.patsel0_low_q[18] ),
    .A2(_01834_),
    .B1(_01835_),
    .Y(_01841_));
 sky130_fd_sc_hd__a31o_1 _18591_ (.A1(_01839_),
    .A2(_01840_),
    .A3(_01841_),
    .B1(_01837_),
    .X(_01842_));
 sky130_fd_sc_hd__o21ba_1 _18592_ (.A1(\wfg_drive_pat_top.wbs_dat_o[18] ),
    .A2(_01753_),
    .B1_N(_01842_),
    .X(_00625_));
 sky130_fd_sc_hd__nand2_1 _18593_ (.A(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[19].drv.ctrl_en_q_i ),
    .B(_01768_),
    .Y(_01843_));
 sky130_fd_sc_hd__nand2_1 _18594_ (.A(\wfg_drive_pat_top.patsel1_high_q[19] ),
    .B(_01815_),
    .Y(_01844_));
 sky130_fd_sc_hd__a21oi_1 _18595_ (.A1(\wfg_drive_pat_top.patsel0_low_q[19] ),
    .A2(_01834_),
    .B1(_01835_),
    .Y(_01845_));
 sky130_fd_sc_hd__a31o_1 _18596_ (.A1(_01843_),
    .A2(_01844_),
    .A3(_01845_),
    .B1(_01837_),
    .X(_01846_));
 sky130_fd_sc_hd__o21ba_1 _18597_ (.A1(\wfg_drive_pat_top.wbs_dat_o[19] ),
    .A2(_01753_),
    .B1_N(_01846_),
    .X(_00626_));
 sky130_fd_sc_hd__nand2_1 _18598_ (.A(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[20].drv.ctrl_en_q_i ),
    .B(_01768_),
    .Y(_01847_));
 sky130_fd_sc_hd__nand2_1 _18599_ (.A(\wfg_drive_pat_top.patsel1_high_q[20] ),
    .B(_01815_),
    .Y(_01848_));
 sky130_fd_sc_hd__a21oi_1 _18600_ (.A1(\wfg_drive_pat_top.patsel0_low_q[20] ),
    .A2(_01834_),
    .B1(_01835_),
    .Y(_01849_));
 sky130_fd_sc_hd__a31o_1 _18601_ (.A1(_01847_),
    .A2(_01848_),
    .A3(_01849_),
    .B1(_01837_),
    .X(_01850_));
 sky130_fd_sc_hd__o21ba_1 _18602_ (.A1(\wfg_drive_pat_top.wbs_dat_o[20] ),
    .A2(_01753_),
    .B1_N(_01850_),
    .X(_00627_));
 sky130_fd_sc_hd__a22o_1 _18603_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[21].drv.ctrl_en_q_i ),
    .A2(_01767_),
    .B1(_01758_),
    .B2(\wfg_drive_pat_top.patsel1_high_q[21] ),
    .X(_01851_));
 sky130_fd_sc_hd__a211o_1 _18604_ (.A1(\wfg_drive_pat_top.patsel0_low_q[21] ),
    .A2(_01834_),
    .B1(_01851_),
    .C1(_01835_),
    .X(_01852_));
 sky130_fd_sc_hd__o211a_1 _18605_ (.A1(\wfg_drive_pat_top.wbs_dat_o[21] ),
    .A2(_01752_),
    .B1(_01852_),
    .C1(_01805_),
    .X(_00628_));
 sky130_fd_sc_hd__nand2_1 _18606_ (.A(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[22].drv.ctrl_en_q_i ),
    .B(_01768_),
    .Y(_01853_));
 sky130_fd_sc_hd__nand2_1 _18607_ (.A(\wfg_drive_pat_top.patsel1_high_q[22] ),
    .B(_01815_),
    .Y(_01854_));
 sky130_fd_sc_hd__a21oi_1 _18608_ (.A1(\wfg_drive_pat_top.patsel0_low_q[22] ),
    .A2(_01777_),
    .B1(_01770_),
    .Y(_01855_));
 sky130_fd_sc_hd__a31o_1 _18609_ (.A1(_01853_),
    .A2(_01854_),
    .A3(_01855_),
    .B1(_01837_),
    .X(_01856_));
 sky130_fd_sc_hd__o21ba_1 _18610_ (.A1(\wfg_drive_pat_top.wbs_dat_o[22] ),
    .A2(_01753_),
    .B1_N(_01856_),
    .X(_00629_));
 sky130_fd_sc_hd__a22o_1 _18611_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[23].drv.ctrl_en_q_i ),
    .A2(_01767_),
    .B1(_01758_),
    .B2(\wfg_drive_pat_top.patsel1_high_q[23] ),
    .X(_01857_));
 sky130_fd_sc_hd__a211o_2 _18612_ (.A1(\wfg_drive_pat_top.patsel0_low_q[23] ),
    .A2(_01834_),
    .B1(_01857_),
    .C1(_01835_),
    .X(_01858_));
 sky130_fd_sc_hd__o211a_1 _18613_ (.A1(\wfg_drive_pat_top.wbs_dat_o[23] ),
    .A2(_01752_),
    .B1(_01858_),
    .C1(_01805_),
    .X(_00630_));
 sky130_fd_sc_hd__a22o_1 _18614_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[24].drv.ctrl_en_q_i ),
    .A2(_01767_),
    .B1(_01758_),
    .B2(\wfg_drive_pat_top.patsel1_high_q[24] ),
    .X(_01859_));
 sky130_fd_sc_hd__a211o_1 _18615_ (.A1(\wfg_drive_pat_top.patsel0_low_q[24] ),
    .A2(_01834_),
    .B1(_01859_),
    .C1(_01835_),
    .X(_01860_));
 sky130_fd_sc_hd__buf_4 _18616_ (.A(_01730_),
    .X(_01861_));
 sky130_fd_sc_hd__o211a_1 _18617_ (.A1(\wfg_drive_pat_top.wbs_dat_o[24] ),
    .A2(_01752_),
    .B1(_01860_),
    .C1(_01861_),
    .X(_00631_));
 sky130_fd_sc_hd__a22o_1 _18618_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[25].drv.ctrl_en_q_i ),
    .A2(_01767_),
    .B1(_01758_),
    .B2(\wfg_drive_pat_top.patsel1_high_q[25] ),
    .X(_01862_));
 sky130_fd_sc_hd__a211o_1 _18619_ (.A1(\wfg_drive_pat_top.patsel0_low_q[25] ),
    .A2(_01834_),
    .B1(_01862_),
    .C1(_01835_),
    .X(_01863_));
 sky130_fd_sc_hd__o211a_1 _18620_ (.A1(\wfg_drive_pat_top.wbs_dat_o[25] ),
    .A2(_01752_),
    .B1(_01863_),
    .C1(_01861_),
    .X(_00632_));
 sky130_fd_sc_hd__nand2_1 _18621_ (.A(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[26].drv.ctrl_en_q_i ),
    .B(_01768_),
    .Y(_01864_));
 sky130_fd_sc_hd__nand2_1 _18622_ (.A(\wfg_drive_pat_top.patsel1_high_q[26] ),
    .B(_01815_),
    .Y(_01865_));
 sky130_fd_sc_hd__a21oi_1 _18623_ (.A1(\wfg_drive_pat_top.patsel0_low_q[26] ),
    .A2(_01777_),
    .B1(_01770_),
    .Y(_01866_));
 sky130_fd_sc_hd__a31o_1 _18624_ (.A1(_01864_),
    .A2(_01865_),
    .A3(_01866_),
    .B1(_01837_),
    .X(_01867_));
 sky130_fd_sc_hd__o21ba_1 _18625_ (.A1(\wfg_drive_pat_top.wbs_dat_o[26] ),
    .A2(_01753_),
    .B1_N(_01867_),
    .X(_00633_));
 sky130_fd_sc_hd__a22o_1 _18626_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[27].drv.ctrl_en_q_i ),
    .A2(_01767_),
    .B1(_01758_),
    .B2(\wfg_drive_pat_top.patsel1_high_q[27] ),
    .X(_01868_));
 sky130_fd_sc_hd__a211o_1 _18627_ (.A1(\wfg_drive_pat_top.patsel0_low_q[27] ),
    .A2(_01834_),
    .B1(_01868_),
    .C1(_01835_),
    .X(_01869_));
 sky130_fd_sc_hd__o211a_1 _18628_ (.A1(\wfg_drive_pat_top.wbs_dat_o[27] ),
    .A2(_01752_),
    .B1(_01869_),
    .C1(_01861_),
    .X(_00634_));
 sky130_fd_sc_hd__a22o_1 _18629_ (.A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[28].drv.ctrl_en_q_i ),
    .A2(_01767_),
    .B1(_01758_),
    .B2(\wfg_drive_pat_top.patsel1_high_q[28] ),
    .X(_01870_));
 sky130_fd_sc_hd__a211o_1 _18630_ (.A1(\wfg_drive_pat_top.patsel0_low_q[28] ),
    .A2(_01834_),
    .B1(_01870_),
    .C1(_01835_),
    .X(_01871_));
 sky130_fd_sc_hd__o211a_1 _18631_ (.A1(\wfg_drive_pat_top.wbs_dat_o[28] ),
    .A2(_01752_),
    .B1(_01871_),
    .C1(_01861_),
    .X(_00635_));
 sky130_fd_sc_hd__nand2_1 _18632_ (.A(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[29].drv.ctrl_en_q_i ),
    .B(_01768_),
    .Y(_01872_));
 sky130_fd_sc_hd__nand2_1 _18633_ (.A(\wfg_drive_pat_top.patsel1_high_q[29] ),
    .B(_01758_),
    .Y(_01873_));
 sky130_fd_sc_hd__a21oi_1 _18634_ (.A1(\wfg_drive_pat_top.patsel0_low_q[29] ),
    .A2(_01777_),
    .B1(_01770_),
    .Y(_01874_));
 sky130_fd_sc_hd__a31o_1 _18635_ (.A1(_01872_),
    .A2(_01873_),
    .A3(_01874_),
    .B1(_01590_),
    .X(_01875_));
 sky130_fd_sc_hd__o21ba_1 _18636_ (.A1(\wfg_drive_pat_top.wbs_dat_o[29] ),
    .A2(_01753_),
    .B1_N(_01875_),
    .X(_00636_));
 sky130_fd_sc_hd__nand2_1 _18637_ (.A(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[30].drv.ctrl_en_q_i ),
    .B(_01768_),
    .Y(_01876_));
 sky130_fd_sc_hd__nand2_1 _18638_ (.A(\wfg_drive_pat_top.patsel1_high_q[30] ),
    .B(_01758_),
    .Y(_01877_));
 sky130_fd_sc_hd__a21oi_1 _18639_ (.A1(\wfg_drive_pat_top.patsel0_low_q[30] ),
    .A2(_01777_),
    .B1(_01770_),
    .Y(_01878_));
 sky130_fd_sc_hd__a31o_1 _18640_ (.A1(_01876_),
    .A2(_01877_),
    .A3(_01878_),
    .B1(_01590_),
    .X(_01879_));
 sky130_fd_sc_hd__o21ba_1 _18641_ (.A1(\wfg_drive_pat_top.wbs_dat_o[30] ),
    .A2(_01753_),
    .B1_N(_01879_),
    .X(_00637_));
 sky130_fd_sc_hd__nand2_1 _18642_ (.A(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[31].drv.ctrl_en_q_i ),
    .B(_01768_),
    .Y(_01880_));
 sky130_fd_sc_hd__nand2_1 _18643_ (.A(\wfg_drive_pat_top.patsel1_high_q[31] ),
    .B(_01758_),
    .Y(_01881_));
 sky130_fd_sc_hd__a21oi_1 _18644_ (.A1(\wfg_drive_pat_top.patsel0_low_q[31] ),
    .A2(_01777_),
    .B1(_01770_),
    .Y(_01882_));
 sky130_fd_sc_hd__a31o_1 _18645_ (.A1(_01880_),
    .A2(_01881_),
    .A3(_01882_),
    .B1(_01590_),
    .X(_01883_));
 sky130_fd_sc_hd__o21ba_1 _18646_ (.A1(\wfg_drive_pat_top.wbs_dat_o[31] ),
    .A2(_01753_),
    .B1_N(_01883_),
    .X(_00638_));
 sky130_fd_sc_hd__buf_6 _18647_ (.A(net66),
    .X(_01884_));
 sky130_fd_sc_hd__and3_1 _18648_ (.A(net61),
    .B(_01610_),
    .C(_01613_),
    .X(_01885_));
 sky130_fd_sc_hd__or3b_1 _18649_ (.A(_01412_),
    .B(_01431_),
    .C_N(_01885_),
    .X(_01886_));
 sky130_fd_sc_hd__or3_2 _18650_ (.A(_01886_),
    .B(_01605_),
    .C(_01607_),
    .X(_01887_));
 sky130_fd_sc_hd__or2_4 _18651_ (.A(_01690_),
    .B(_01887_),
    .X(_01888_));
 sky130_fd_sc_hd__buf_4 _18652_ (.A(_01888_),
    .X(_01889_));
 sky130_fd_sc_hd__mux2_1 _18653_ (.A0(_01884_),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[0].drv.ctrl_en_q_i ),
    .S(_01889_),
    .X(_01890_));
 sky130_fd_sc_hd__and2_1 _18654_ (.A(_01678_),
    .B(_01890_),
    .X(_01891_));
 sky130_fd_sc_hd__clkbuf_1 _18655_ (.A(_01891_),
    .X(_00639_));
 sky130_fd_sc_hd__mux2_1 _18656_ (.A0(_01663_),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[1].drv.ctrl_en_q_i ),
    .S(_01889_),
    .X(_01892_));
 sky130_fd_sc_hd__and2_1 _18657_ (.A(_01678_),
    .B(_01892_),
    .X(_01893_));
 sky130_fd_sc_hd__clkbuf_1 _18658_ (.A(_01893_),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_1 _18659_ (.A0(_01666_),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[2].drv.ctrl_en_q_i ),
    .S(_01889_),
    .X(_01894_));
 sky130_fd_sc_hd__and2_1 _18660_ (.A(_01678_),
    .B(_01894_),
    .X(_01895_));
 sky130_fd_sc_hd__clkbuf_1 _18661_ (.A(_01895_),
    .X(_00641_));
 sky130_fd_sc_hd__mux2_1 _18662_ (.A0(_01669_),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[3].drv.ctrl_en_q_i ),
    .S(_01889_),
    .X(_01896_));
 sky130_fd_sc_hd__and2_1 _18663_ (.A(_01678_),
    .B(_01896_),
    .X(_01897_));
 sky130_fd_sc_hd__clkbuf_1 _18664_ (.A(_01897_),
    .X(_00642_));
 sky130_fd_sc_hd__mux2_1 _18665_ (.A0(_01672_),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[4].drv.ctrl_en_q_i ),
    .S(_01889_),
    .X(_01898_));
 sky130_fd_sc_hd__and2_1 _18666_ (.A(_01678_),
    .B(_01898_),
    .X(_01899_));
 sky130_fd_sc_hd__clkbuf_1 _18667_ (.A(_01899_),
    .X(_00643_));
 sky130_fd_sc_hd__mux2_1 _18668_ (.A0(_01675_),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[5].drv.ctrl_en_q_i ),
    .S(_01889_),
    .X(_01900_));
 sky130_fd_sc_hd__and2_1 _18669_ (.A(_01678_),
    .B(_01900_),
    .X(_01901_));
 sky130_fd_sc_hd__clkbuf_1 _18670_ (.A(_01901_),
    .X(_00644_));
 sky130_fd_sc_hd__mux2_1 _18671_ (.A0(_01679_),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[6].drv.ctrl_en_q_i ),
    .S(_01889_),
    .X(_01902_));
 sky130_fd_sc_hd__and2_1 _18672_ (.A(_01678_),
    .B(_01902_),
    .X(_01903_));
 sky130_fd_sc_hd__clkbuf_1 _18673_ (.A(_01903_),
    .X(_00645_));
 sky130_fd_sc_hd__mux2_1 _18674_ (.A0(_01682_),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[7].drv.ctrl_en_q_i ),
    .S(_01889_),
    .X(_01904_));
 sky130_fd_sc_hd__and2_1 _18675_ (.A(_01678_),
    .B(_01904_),
    .X(_01905_));
 sky130_fd_sc_hd__clkbuf_1 _18676_ (.A(_01905_),
    .X(_00646_));
 sky130_fd_sc_hd__buf_2 _18677_ (.A(_01599_),
    .X(_01906_));
 sky130_fd_sc_hd__mux2_1 _18678_ (.A0(_01601_),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[8].drv.ctrl_en_q_i ),
    .S(_01889_),
    .X(_01907_));
 sky130_fd_sc_hd__and2_1 _18679_ (.A(_01906_),
    .B(_01907_),
    .X(_01908_));
 sky130_fd_sc_hd__clkbuf_1 _18680_ (.A(_01908_),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_1 _18681_ (.A0(_01620_),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[9].drv.ctrl_en_q_i ),
    .S(_01889_),
    .X(_01909_));
 sky130_fd_sc_hd__and2_1 _18682_ (.A(_01906_),
    .B(_01909_),
    .X(_01910_));
 sky130_fd_sc_hd__clkbuf_1 _18683_ (.A(_01910_),
    .X(_00648_));
 sky130_fd_sc_hd__buf_4 _18684_ (.A(_01888_),
    .X(_01911_));
 sky130_fd_sc_hd__mux2_1 _18685_ (.A0(_01624_),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[10].drv.ctrl_en_q_i ),
    .S(_01911_),
    .X(_01912_));
 sky130_fd_sc_hd__and2_1 _18686_ (.A(_01906_),
    .B(_01912_),
    .X(_01913_));
 sky130_fd_sc_hd__clkbuf_1 _18687_ (.A(_01913_),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_1 _18688_ (.A0(_01627_),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[11].drv.ctrl_en_q_i ),
    .S(_01911_),
    .X(_01914_));
 sky130_fd_sc_hd__and2_1 _18689_ (.A(_01906_),
    .B(_01914_),
    .X(_01915_));
 sky130_fd_sc_hd__clkbuf_1 _18690_ (.A(_01915_),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_1 _18691_ (.A0(_01630_),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[12].drv.ctrl_en_q_i ),
    .S(_01911_),
    .X(_01916_));
 sky130_fd_sc_hd__and2_1 _18692_ (.A(_01906_),
    .B(_01916_),
    .X(_01917_));
 sky130_fd_sc_hd__clkbuf_1 _18693_ (.A(_01917_),
    .X(_00651_));
 sky130_fd_sc_hd__mux2_1 _18694_ (.A0(_01633_),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[13].drv.ctrl_en_q_i ),
    .S(_01911_),
    .X(_01918_));
 sky130_fd_sc_hd__and2_1 _18695_ (.A(_01906_),
    .B(_01918_),
    .X(_01919_));
 sky130_fd_sc_hd__clkbuf_1 _18696_ (.A(_01919_),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_1 _18697_ (.A0(_01636_),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[14].drv.ctrl_en_q_i ),
    .S(_01911_),
    .X(_01920_));
 sky130_fd_sc_hd__and2_1 _18698_ (.A(_01906_),
    .B(_01920_),
    .X(_01921_));
 sky130_fd_sc_hd__clkbuf_1 _18699_ (.A(_01921_),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _18700_ (.A0(_01639_),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[15].drv.ctrl_en_q_i ),
    .S(_01911_),
    .X(_01922_));
 sky130_fd_sc_hd__and2_1 _18701_ (.A(_01906_),
    .B(_01922_),
    .X(_01923_));
 sky130_fd_sc_hd__clkbuf_1 _18702_ (.A(_01923_),
    .X(_00654_));
 sky130_fd_sc_hd__mux2_1 _18703_ (.A0(net73),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[16].drv.ctrl_en_q_i ),
    .S(_01911_),
    .X(_01924_));
 sky130_fd_sc_hd__and2_1 _18704_ (.A(_01906_),
    .B(_01924_),
    .X(_01925_));
 sky130_fd_sc_hd__clkbuf_1 _18705_ (.A(_01925_),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_1 _18706_ (.A0(net74),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[17].drv.ctrl_en_q_i ),
    .S(_01911_),
    .X(_01926_));
 sky130_fd_sc_hd__and2_1 _18707_ (.A(_01906_),
    .B(_01926_),
    .X(_01927_));
 sky130_fd_sc_hd__clkbuf_1 _18708_ (.A(_01927_),
    .X(_00656_));
 sky130_fd_sc_hd__buf_2 _18709_ (.A(_01599_),
    .X(_01928_));
 sky130_fd_sc_hd__mux2_1 _18710_ (.A0(net75),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[18].drv.ctrl_en_q_i ),
    .S(_01911_),
    .X(_01929_));
 sky130_fd_sc_hd__and2_1 _18711_ (.A(_01928_),
    .B(_01929_),
    .X(_01930_));
 sky130_fd_sc_hd__clkbuf_1 _18712_ (.A(_01930_),
    .X(_00657_));
 sky130_fd_sc_hd__mux2_1 _18713_ (.A0(net76),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[19].drv.ctrl_en_q_i ),
    .S(_01911_),
    .X(_01931_));
 sky130_fd_sc_hd__and2_1 _18714_ (.A(_01928_),
    .B(_01931_),
    .X(_01932_));
 sky130_fd_sc_hd__clkbuf_1 _18715_ (.A(_01932_),
    .X(_00658_));
 sky130_fd_sc_hd__buf_4 _18716_ (.A(_01888_),
    .X(_01933_));
 sky130_fd_sc_hd__mux2_1 _18717_ (.A0(net78),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[20].drv.ctrl_en_q_i ),
    .S(_01933_),
    .X(_01934_));
 sky130_fd_sc_hd__and2_1 _18718_ (.A(_01928_),
    .B(_01934_),
    .X(_01935_));
 sky130_fd_sc_hd__clkbuf_1 _18719_ (.A(_01935_),
    .X(_00659_));
 sky130_fd_sc_hd__mux2_1 _18720_ (.A0(net79),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[21].drv.ctrl_en_q_i ),
    .S(_01933_),
    .X(_01936_));
 sky130_fd_sc_hd__and2_1 _18721_ (.A(_01928_),
    .B(_01936_),
    .X(_01937_));
 sky130_fd_sc_hd__clkbuf_1 _18722_ (.A(_01937_),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_1 _18723_ (.A0(net80),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[22].drv.ctrl_en_q_i ),
    .S(_01933_),
    .X(_01938_));
 sky130_fd_sc_hd__and2_1 _18724_ (.A(_01928_),
    .B(_01938_),
    .X(_01939_));
 sky130_fd_sc_hd__clkbuf_1 _18725_ (.A(_01939_),
    .X(_00661_));
 sky130_fd_sc_hd__mux2_1 _18726_ (.A0(net81),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[23].drv.ctrl_en_q_i ),
    .S(_01933_),
    .X(_01940_));
 sky130_fd_sc_hd__and2_1 _18727_ (.A(_01928_),
    .B(_01940_),
    .X(_01941_));
 sky130_fd_sc_hd__clkbuf_1 _18728_ (.A(_01941_),
    .X(_00662_));
 sky130_fd_sc_hd__mux2_1 _18729_ (.A0(net82),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[24].drv.ctrl_en_q_i ),
    .S(_01933_),
    .X(_01942_));
 sky130_fd_sc_hd__and2_1 _18730_ (.A(_01928_),
    .B(_01942_),
    .X(_01943_));
 sky130_fd_sc_hd__clkbuf_1 _18731_ (.A(_01943_),
    .X(_00663_));
 sky130_fd_sc_hd__mux2_1 _18732_ (.A0(net83),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[25].drv.ctrl_en_q_i ),
    .S(_01933_),
    .X(_01944_));
 sky130_fd_sc_hd__and2_1 _18733_ (.A(_01928_),
    .B(_01944_),
    .X(_01945_));
 sky130_fd_sc_hd__clkbuf_1 _18734_ (.A(_01945_),
    .X(_00664_));
 sky130_fd_sc_hd__mux2_1 _18735_ (.A0(net84),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[26].drv.ctrl_en_q_i ),
    .S(_01933_),
    .X(_01946_));
 sky130_fd_sc_hd__and2_1 _18736_ (.A(_01928_),
    .B(_01946_),
    .X(_01947_));
 sky130_fd_sc_hd__clkbuf_1 _18737_ (.A(_01947_),
    .X(_00665_));
 sky130_fd_sc_hd__mux2_1 _18738_ (.A0(net85),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[27].drv.ctrl_en_q_i ),
    .S(_01933_),
    .X(_01948_));
 sky130_fd_sc_hd__and2_1 _18739_ (.A(_01928_),
    .B(_01948_),
    .X(_01949_));
 sky130_fd_sc_hd__clkbuf_1 _18740_ (.A(_01949_),
    .X(_00666_));
 sky130_fd_sc_hd__buf_4 _18741_ (.A(_01599_),
    .X(_01950_));
 sky130_fd_sc_hd__mux2_1 _18742_ (.A0(net86),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[28].drv.ctrl_en_q_i ),
    .S(_01933_),
    .X(_01951_));
 sky130_fd_sc_hd__and2_1 _18743_ (.A(_01950_),
    .B(_01951_),
    .X(_01952_));
 sky130_fd_sc_hd__clkbuf_1 _18744_ (.A(_01952_),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_1 _18745_ (.A0(net87),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[29].drv.ctrl_en_q_i ),
    .S(_01933_),
    .X(_01953_));
 sky130_fd_sc_hd__and2_1 _18746_ (.A(_01950_),
    .B(_01953_),
    .X(_01954_));
 sky130_fd_sc_hd__clkbuf_1 _18747_ (.A(_01954_),
    .X(_00668_));
 sky130_fd_sc_hd__mux2_1 _18748_ (.A0(net89),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[30].drv.ctrl_en_q_i ),
    .S(_01888_),
    .X(_01955_));
 sky130_fd_sc_hd__and2_1 _18749_ (.A(_01950_),
    .B(_01955_),
    .X(_01956_));
 sky130_fd_sc_hd__clkbuf_1 _18750_ (.A(_01956_),
    .X(_00669_));
 sky130_fd_sc_hd__mux2_1 _18751_ (.A0(net90),
    .A1(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[31].drv.ctrl_en_q_i ),
    .S(_01888_),
    .X(_01957_));
 sky130_fd_sc_hd__and2_1 _18752_ (.A(_01950_),
    .B(_01957_),
    .X(_01958_));
 sky130_fd_sc_hd__clkbuf_1 _18753_ (.A(_01958_),
    .X(_00670_));
 sky130_fd_sc_hd__buf_4 _18754_ (.A(_01604_),
    .X(_01959_));
 sky130_fd_sc_hd__or2_2 _18755_ (.A(_01959_),
    .B(_01887_),
    .X(_01960_));
 sky130_fd_sc_hd__clkbuf_4 _18756_ (.A(_01960_),
    .X(_01961_));
 sky130_fd_sc_hd__mux2_1 _18757_ (.A0(net73),
    .A1(_09782_),
    .S(_01961_),
    .X(_01962_));
 sky130_fd_sc_hd__and2_1 _18758_ (.A(_01950_),
    .B(_01962_),
    .X(_01963_));
 sky130_fd_sc_hd__clkbuf_1 _18759_ (.A(_01963_),
    .X(_00671_));
 sky130_fd_sc_hd__buf_2 _18760_ (.A(_01961_),
    .X(_01964_));
 sky130_fd_sc_hd__nand2_1 _18761_ (.A(_09814_),
    .B(_01964_),
    .Y(_01965_));
 sky130_fd_sc_hd__o211a_1 _18762_ (.A1(_01660_),
    .A2(_01964_),
    .B1(_01965_),
    .C1(_01861_),
    .X(_00672_));
 sky130_fd_sc_hd__mux2_1 _18763_ (.A0(_01663_),
    .A1(\wfg_drive_pat_top.cfg_begin_q[1] ),
    .S(_01961_),
    .X(_01966_));
 sky130_fd_sc_hd__and2_1 _18764_ (.A(_01950_),
    .B(_01966_),
    .X(_01967_));
 sky130_fd_sc_hd__clkbuf_1 _18765_ (.A(_01967_),
    .X(_00673_));
 sky130_fd_sc_hd__mux2_1 _18766_ (.A0(_01666_),
    .A1(\wfg_drive_pat_top.cfg_begin_q[2] ),
    .S(_01961_),
    .X(_01968_));
 sky130_fd_sc_hd__and2_1 _18767_ (.A(_01950_),
    .B(_01968_),
    .X(_01969_));
 sky130_fd_sc_hd__clkbuf_1 _18768_ (.A(_01969_),
    .X(_00674_));
 sky130_fd_sc_hd__mux2_1 _18769_ (.A0(_01669_),
    .A1(\wfg_drive_pat_top.cfg_begin_q[3] ),
    .S(_01961_),
    .X(_01970_));
 sky130_fd_sc_hd__and2_1 _18770_ (.A(_01950_),
    .B(_01970_),
    .X(_01971_));
 sky130_fd_sc_hd__clkbuf_1 _18771_ (.A(_01971_),
    .X(_00675_));
 sky130_fd_sc_hd__mux2_1 _18772_ (.A0(_01672_),
    .A1(\wfg_drive_pat_top.cfg_begin_q[4] ),
    .S(_01961_),
    .X(_01972_));
 sky130_fd_sc_hd__and2_1 _18773_ (.A(_01950_),
    .B(_01972_),
    .X(_01973_));
 sky130_fd_sc_hd__clkbuf_1 _18774_ (.A(_01973_),
    .X(_00676_));
 sky130_fd_sc_hd__mux2_1 _18775_ (.A0(_01675_),
    .A1(\wfg_drive_pat_top.cfg_begin_q[5] ),
    .S(_01961_),
    .X(_01974_));
 sky130_fd_sc_hd__and2_1 _18776_ (.A(_01950_),
    .B(_01974_),
    .X(_01975_));
 sky130_fd_sc_hd__clkbuf_1 _18777_ (.A(_01975_),
    .X(_00677_));
 sky130_fd_sc_hd__nand2_1 _18778_ (.A(_09815_),
    .B(_01964_),
    .Y(_01976_));
 sky130_fd_sc_hd__o211a_1 _18779_ (.A1(_01679_),
    .A2(_01964_),
    .B1(_01976_),
    .C1(_01861_),
    .X(_00678_));
 sky130_fd_sc_hd__nand2_1 _18780_ (.A(_09811_),
    .B(_01964_),
    .Y(_01977_));
 sky130_fd_sc_hd__o211a_1 _18781_ (.A1(_01682_),
    .A2(_01964_),
    .B1(_01977_),
    .C1(_01861_),
    .X(_00679_));
 sky130_fd_sc_hd__nand2_1 _18782_ (.A(_09793_),
    .B(_01964_),
    .Y(_01978_));
 sky130_fd_sc_hd__o211a_1 _18783_ (.A1(_01601_),
    .A2(_01964_),
    .B1(_01978_),
    .C1(_01861_),
    .X(_00680_));
 sky130_fd_sc_hd__buf_2 _18784_ (.A(_01599_),
    .X(_01979_));
 sky130_fd_sc_hd__mux2_1 _18785_ (.A0(_01620_),
    .A1(\wfg_drive_pat_top.cfg_end_q[9] ),
    .S(_01961_),
    .X(_01980_));
 sky130_fd_sc_hd__and2_1 _18786_ (.A(_01979_),
    .B(_01980_),
    .X(_01981_));
 sky130_fd_sc_hd__clkbuf_1 _18787_ (.A(_01981_),
    .X(_00681_));
 sky130_fd_sc_hd__mux2_1 _18788_ (.A0(_01624_),
    .A1(\wfg_drive_pat_top.cfg_end_q[10] ),
    .S(_01960_),
    .X(_01982_));
 sky130_fd_sc_hd__and2_1 _18789_ (.A(_01979_),
    .B(_01982_),
    .X(_01983_));
 sky130_fd_sc_hd__clkbuf_1 _18790_ (.A(_01983_),
    .X(_00682_));
 sky130_fd_sc_hd__mux2_1 _18791_ (.A0(_01627_),
    .A1(\wfg_drive_pat_top.cfg_end_q[11] ),
    .S(_01960_),
    .X(_01984_));
 sky130_fd_sc_hd__and2_1 _18792_ (.A(_01979_),
    .B(_01984_),
    .X(_01985_));
 sky130_fd_sc_hd__clkbuf_1 _18793_ (.A(_01985_),
    .X(_00683_));
 sky130_fd_sc_hd__mux2_1 _18794_ (.A0(_01630_),
    .A1(\wfg_drive_pat_top.cfg_end_q[12] ),
    .S(_01960_),
    .X(_01986_));
 sky130_fd_sc_hd__and2_1 _18795_ (.A(_01979_),
    .B(_01986_),
    .X(_01987_));
 sky130_fd_sc_hd__clkbuf_1 _18796_ (.A(_01987_),
    .X(_00684_));
 sky130_fd_sc_hd__nand2_1 _18797_ (.A(_09775_),
    .B(_01961_),
    .Y(_01988_));
 sky130_fd_sc_hd__o211a_1 _18798_ (.A1(_01633_),
    .A2(_01964_),
    .B1(_01988_),
    .C1(_01861_),
    .X(_00685_));
 sky130_fd_sc_hd__mux2_1 _18799_ (.A0(_01636_),
    .A1(\wfg_drive_pat_top.cfg_end_q[14] ),
    .S(_01960_),
    .X(_01989_));
 sky130_fd_sc_hd__and2_1 _18800_ (.A(_01979_),
    .B(_01989_),
    .X(_01990_));
 sky130_fd_sc_hd__clkbuf_1 _18801_ (.A(_01990_),
    .X(_00686_));
 sky130_fd_sc_hd__nand2_1 _18802_ (.A(_09778_),
    .B(_01961_),
    .Y(_01991_));
 sky130_fd_sc_hd__o211a_1 _18803_ (.A1(_01639_),
    .A2(_01964_),
    .B1(_01991_),
    .C1(_01861_),
    .X(_00687_));
 sky130_fd_sc_hd__or2_4 _18804_ (.A(_01762_),
    .B(_01887_),
    .X(_01992_));
 sky130_fd_sc_hd__buf_4 _18805_ (.A(_01992_),
    .X(_01993_));
 sky130_fd_sc_hd__mux2_1 _18806_ (.A0(_01884_),
    .A1(\wfg_drive_pat_top.patsel0_low_q[0] ),
    .S(_01993_),
    .X(_01994_));
 sky130_fd_sc_hd__and2_1 _18807_ (.A(_01979_),
    .B(_01994_),
    .X(_01995_));
 sky130_fd_sc_hd__clkbuf_1 _18808_ (.A(_01995_),
    .X(_00688_));
 sky130_fd_sc_hd__mux2_1 _18809_ (.A0(_01663_),
    .A1(\wfg_drive_pat_top.patsel0_low_q[1] ),
    .S(_01993_),
    .X(_01996_));
 sky130_fd_sc_hd__and2_1 _18810_ (.A(_01979_),
    .B(_01996_),
    .X(_01997_));
 sky130_fd_sc_hd__clkbuf_1 _18811_ (.A(_01997_),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_1 _18812_ (.A0(_01666_),
    .A1(\wfg_drive_pat_top.patsel0_low_q[2] ),
    .S(_01993_),
    .X(_01998_));
 sky130_fd_sc_hd__and2_1 _18813_ (.A(_01979_),
    .B(_01998_),
    .X(_01999_));
 sky130_fd_sc_hd__clkbuf_1 _18814_ (.A(_01999_),
    .X(_00690_));
 sky130_fd_sc_hd__mux2_1 _18815_ (.A0(_01669_),
    .A1(\wfg_drive_pat_top.patsel0_low_q[3] ),
    .S(_01993_),
    .X(_02000_));
 sky130_fd_sc_hd__and2_1 _18816_ (.A(_01979_),
    .B(_02000_),
    .X(_02001_));
 sky130_fd_sc_hd__clkbuf_1 _18817_ (.A(_02001_),
    .X(_00691_));
 sky130_fd_sc_hd__mux2_1 _18818_ (.A0(_01672_),
    .A1(\wfg_drive_pat_top.patsel0_low_q[4] ),
    .S(_01993_),
    .X(_02002_));
 sky130_fd_sc_hd__and2_1 _18819_ (.A(_01979_),
    .B(_02002_),
    .X(_02003_));
 sky130_fd_sc_hd__clkbuf_1 _18820_ (.A(_02003_),
    .X(_00692_));
 sky130_fd_sc_hd__buf_2 _18821_ (.A(_01599_),
    .X(_02004_));
 sky130_fd_sc_hd__mux2_1 _18822_ (.A0(_01675_),
    .A1(\wfg_drive_pat_top.patsel0_low_q[5] ),
    .S(_01993_),
    .X(_02005_));
 sky130_fd_sc_hd__and2_1 _18823_ (.A(_02004_),
    .B(_02005_),
    .X(_02006_));
 sky130_fd_sc_hd__clkbuf_1 _18824_ (.A(_02006_),
    .X(_00693_));
 sky130_fd_sc_hd__mux2_1 _18825_ (.A0(_01679_),
    .A1(\wfg_drive_pat_top.patsel0_low_q[6] ),
    .S(_01993_),
    .X(_02007_));
 sky130_fd_sc_hd__and2_1 _18826_ (.A(_02004_),
    .B(_02007_),
    .X(_02008_));
 sky130_fd_sc_hd__clkbuf_1 _18827_ (.A(_02008_),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_1 _18828_ (.A0(_01682_),
    .A1(\wfg_drive_pat_top.patsel0_low_q[7] ),
    .S(_01993_),
    .X(_02009_));
 sky130_fd_sc_hd__and2_1 _18829_ (.A(_02004_),
    .B(_02009_),
    .X(_02010_));
 sky130_fd_sc_hd__clkbuf_1 _18830_ (.A(_02010_),
    .X(_00695_));
 sky130_fd_sc_hd__mux2_1 _18831_ (.A0(_01601_),
    .A1(\wfg_drive_pat_top.patsel0_low_q[8] ),
    .S(_01993_),
    .X(_02011_));
 sky130_fd_sc_hd__and2_1 _18832_ (.A(_02004_),
    .B(_02011_),
    .X(_02012_));
 sky130_fd_sc_hd__clkbuf_1 _18833_ (.A(_02012_),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_1 _18834_ (.A0(_01620_),
    .A1(\wfg_drive_pat_top.patsel0_low_q[9] ),
    .S(_01993_),
    .X(_02013_));
 sky130_fd_sc_hd__and2_1 _18835_ (.A(_02004_),
    .B(_02013_),
    .X(_02014_));
 sky130_fd_sc_hd__clkbuf_1 _18836_ (.A(_02014_),
    .X(_00697_));
 sky130_fd_sc_hd__buf_4 _18837_ (.A(_01992_),
    .X(_02015_));
 sky130_fd_sc_hd__mux2_1 _18838_ (.A0(_01624_),
    .A1(\wfg_drive_pat_top.patsel0_low_q[10] ),
    .S(_02015_),
    .X(_02016_));
 sky130_fd_sc_hd__and2_1 _18839_ (.A(_02004_),
    .B(_02016_),
    .X(_02017_));
 sky130_fd_sc_hd__clkbuf_1 _18840_ (.A(_02017_),
    .X(_00698_));
 sky130_fd_sc_hd__mux2_1 _18841_ (.A0(_01627_),
    .A1(\wfg_drive_pat_top.patsel0_low_q[11] ),
    .S(_02015_),
    .X(_02018_));
 sky130_fd_sc_hd__and2_1 _18842_ (.A(_02004_),
    .B(_02018_),
    .X(_02019_));
 sky130_fd_sc_hd__clkbuf_1 _18843_ (.A(_02019_),
    .X(_00699_));
 sky130_fd_sc_hd__mux2_1 _18844_ (.A0(_01630_),
    .A1(\wfg_drive_pat_top.patsel0_low_q[12] ),
    .S(_02015_),
    .X(_02020_));
 sky130_fd_sc_hd__and2_1 _18845_ (.A(_02004_),
    .B(_02020_),
    .X(_02021_));
 sky130_fd_sc_hd__clkbuf_1 _18846_ (.A(_02021_),
    .X(_00700_));
 sky130_fd_sc_hd__mux2_1 _18847_ (.A0(_01633_),
    .A1(\wfg_drive_pat_top.patsel0_low_q[13] ),
    .S(_02015_),
    .X(_02022_));
 sky130_fd_sc_hd__and2_1 _18848_ (.A(_02004_),
    .B(_02022_),
    .X(_02023_));
 sky130_fd_sc_hd__clkbuf_1 _18849_ (.A(_02023_),
    .X(_00701_));
 sky130_fd_sc_hd__mux2_1 _18850_ (.A0(_01636_),
    .A1(\wfg_drive_pat_top.patsel0_low_q[14] ),
    .S(_02015_),
    .X(_02024_));
 sky130_fd_sc_hd__and2_1 _18851_ (.A(_02004_),
    .B(_02024_),
    .X(_02025_));
 sky130_fd_sc_hd__clkbuf_1 _18852_ (.A(_02025_),
    .X(_00702_));
 sky130_fd_sc_hd__buf_2 _18853_ (.A(_01599_),
    .X(_02026_));
 sky130_fd_sc_hd__mux2_1 _18854_ (.A0(_01639_),
    .A1(\wfg_drive_pat_top.patsel0_low_q[15] ),
    .S(_02015_),
    .X(_02027_));
 sky130_fd_sc_hd__and2_1 _18855_ (.A(_02026_),
    .B(_02027_),
    .X(_02028_));
 sky130_fd_sc_hd__clkbuf_1 _18856_ (.A(_02028_),
    .X(_00703_));
 sky130_fd_sc_hd__mux2_1 _18857_ (.A0(net73),
    .A1(\wfg_drive_pat_top.patsel0_low_q[16] ),
    .S(_02015_),
    .X(_02029_));
 sky130_fd_sc_hd__and2_1 _18858_ (.A(_02026_),
    .B(_02029_),
    .X(_02030_));
 sky130_fd_sc_hd__clkbuf_1 _18859_ (.A(_02030_),
    .X(_00704_));
 sky130_fd_sc_hd__mux2_1 _18860_ (.A0(net74),
    .A1(\wfg_drive_pat_top.patsel0_low_q[17] ),
    .S(_02015_),
    .X(_02031_));
 sky130_fd_sc_hd__and2_1 _18861_ (.A(_02026_),
    .B(_02031_),
    .X(_02032_));
 sky130_fd_sc_hd__clkbuf_1 _18862_ (.A(_02032_),
    .X(_00705_));
 sky130_fd_sc_hd__mux2_1 _18863_ (.A0(net75),
    .A1(\wfg_drive_pat_top.patsel0_low_q[18] ),
    .S(_02015_),
    .X(_02033_));
 sky130_fd_sc_hd__and2_1 _18864_ (.A(_02026_),
    .B(_02033_),
    .X(_02034_));
 sky130_fd_sc_hd__clkbuf_1 _18865_ (.A(_02034_),
    .X(_00706_));
 sky130_fd_sc_hd__mux2_1 _18866_ (.A0(net76),
    .A1(\wfg_drive_pat_top.patsel0_low_q[19] ),
    .S(_02015_),
    .X(_02035_));
 sky130_fd_sc_hd__and2_1 _18867_ (.A(_02026_),
    .B(_02035_),
    .X(_02036_));
 sky130_fd_sc_hd__clkbuf_1 _18868_ (.A(_02036_),
    .X(_00707_));
 sky130_fd_sc_hd__buf_4 _18869_ (.A(_01992_),
    .X(_02037_));
 sky130_fd_sc_hd__mux2_1 _18870_ (.A0(net78),
    .A1(\wfg_drive_pat_top.patsel0_low_q[20] ),
    .S(_02037_),
    .X(_02038_));
 sky130_fd_sc_hd__and2_1 _18871_ (.A(_02026_),
    .B(_02038_),
    .X(_02039_));
 sky130_fd_sc_hd__clkbuf_1 _18872_ (.A(_02039_),
    .X(_00708_));
 sky130_fd_sc_hd__mux2_1 _18873_ (.A0(net79),
    .A1(\wfg_drive_pat_top.patsel0_low_q[21] ),
    .S(_02037_),
    .X(_02040_));
 sky130_fd_sc_hd__and2_1 _18874_ (.A(_02026_),
    .B(_02040_),
    .X(_02041_));
 sky130_fd_sc_hd__clkbuf_1 _18875_ (.A(_02041_),
    .X(_00709_));
 sky130_fd_sc_hd__mux2_1 _18876_ (.A0(net80),
    .A1(\wfg_drive_pat_top.patsel0_low_q[22] ),
    .S(_02037_),
    .X(_02042_));
 sky130_fd_sc_hd__and2_1 _18877_ (.A(_02026_),
    .B(_02042_),
    .X(_02043_));
 sky130_fd_sc_hd__clkbuf_1 _18878_ (.A(_02043_),
    .X(_00710_));
 sky130_fd_sc_hd__mux2_1 _18879_ (.A0(net81),
    .A1(\wfg_drive_pat_top.patsel0_low_q[23] ),
    .S(_02037_),
    .X(_02044_));
 sky130_fd_sc_hd__and2_1 _18880_ (.A(_02026_),
    .B(_02044_),
    .X(_02045_));
 sky130_fd_sc_hd__clkbuf_1 _18881_ (.A(_02045_),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_1 _18882_ (.A0(net82),
    .A1(\wfg_drive_pat_top.patsel0_low_q[24] ),
    .S(_02037_),
    .X(_02046_));
 sky130_fd_sc_hd__and2_1 _18883_ (.A(_02026_),
    .B(_02046_),
    .X(_02047_));
 sky130_fd_sc_hd__clkbuf_1 _18884_ (.A(_02047_),
    .X(_00712_));
 sky130_fd_sc_hd__buf_6 _18885_ (.A(_01588_),
    .X(_02048_));
 sky130_fd_sc_hd__clkbuf_4 _18886_ (.A(_02048_),
    .X(_02049_));
 sky130_fd_sc_hd__mux2_1 _18887_ (.A0(net83),
    .A1(\wfg_drive_pat_top.patsel0_low_q[25] ),
    .S(_02037_),
    .X(_02050_));
 sky130_fd_sc_hd__and2_1 _18888_ (.A(_02049_),
    .B(_02050_),
    .X(_02051_));
 sky130_fd_sc_hd__clkbuf_1 _18889_ (.A(_02051_),
    .X(_00713_));
 sky130_fd_sc_hd__mux2_1 _18890_ (.A0(net84),
    .A1(\wfg_drive_pat_top.patsel0_low_q[26] ),
    .S(_02037_),
    .X(_02052_));
 sky130_fd_sc_hd__and2_1 _18891_ (.A(_02049_),
    .B(_02052_),
    .X(_02053_));
 sky130_fd_sc_hd__clkbuf_1 _18892_ (.A(_02053_),
    .X(_00714_));
 sky130_fd_sc_hd__mux2_1 _18893_ (.A0(net85),
    .A1(\wfg_drive_pat_top.patsel0_low_q[27] ),
    .S(_02037_),
    .X(_02054_));
 sky130_fd_sc_hd__and2_1 _18894_ (.A(_02049_),
    .B(_02054_),
    .X(_02055_));
 sky130_fd_sc_hd__clkbuf_1 _18895_ (.A(_02055_),
    .X(_00715_));
 sky130_fd_sc_hd__mux2_1 _18896_ (.A0(net86),
    .A1(\wfg_drive_pat_top.patsel0_low_q[28] ),
    .S(_02037_),
    .X(_02056_));
 sky130_fd_sc_hd__and2_1 _18897_ (.A(_02049_),
    .B(_02056_),
    .X(_02057_));
 sky130_fd_sc_hd__clkbuf_1 _18898_ (.A(_02057_),
    .X(_00716_));
 sky130_fd_sc_hd__mux2_1 _18899_ (.A0(net87),
    .A1(\wfg_drive_pat_top.patsel0_low_q[29] ),
    .S(_02037_),
    .X(_02058_));
 sky130_fd_sc_hd__and2_1 _18900_ (.A(_02049_),
    .B(_02058_),
    .X(_02059_));
 sky130_fd_sc_hd__clkbuf_1 _18901_ (.A(_02059_),
    .X(_00717_));
 sky130_fd_sc_hd__mux2_1 _18902_ (.A0(net89),
    .A1(\wfg_drive_pat_top.patsel0_low_q[30] ),
    .S(_01992_),
    .X(_02060_));
 sky130_fd_sc_hd__and2_1 _18903_ (.A(_02049_),
    .B(_02060_),
    .X(_02061_));
 sky130_fd_sc_hd__clkbuf_1 _18904_ (.A(_02061_),
    .X(_00718_));
 sky130_fd_sc_hd__mux2_1 _18905_ (.A0(net90),
    .A1(\wfg_drive_pat_top.patsel0_low_q[31] ),
    .S(_01992_),
    .X(_02062_));
 sky130_fd_sc_hd__and2_1 _18906_ (.A(_02049_),
    .B(_02062_),
    .X(_02063_));
 sky130_fd_sc_hd__clkbuf_1 _18907_ (.A(_02063_),
    .X(_00719_));
 sky130_fd_sc_hd__or3_4 _18908_ (.A(_01886_),
    .B(_01756_),
    .C(_01887_),
    .X(_02064_));
 sky130_fd_sc_hd__buf_4 _18909_ (.A(_02064_),
    .X(_02065_));
 sky130_fd_sc_hd__mux2_1 _18910_ (.A0(_01884_),
    .A1(\wfg_drive_pat_top.patsel1_high_q[0] ),
    .S(_02065_),
    .X(_02066_));
 sky130_fd_sc_hd__and2_1 _18911_ (.A(_02049_),
    .B(_02066_),
    .X(_02067_));
 sky130_fd_sc_hd__clkbuf_1 _18912_ (.A(_02067_),
    .X(_00720_));
 sky130_fd_sc_hd__mux2_1 _18913_ (.A0(net77),
    .A1(\wfg_drive_pat_top.patsel1_high_q[1] ),
    .S(_02065_),
    .X(_02068_));
 sky130_fd_sc_hd__and2_1 _18914_ (.A(_02049_),
    .B(_02068_),
    .X(_02069_));
 sky130_fd_sc_hd__clkbuf_1 _18915_ (.A(_02069_),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_1 _18916_ (.A0(_01666_),
    .A1(\wfg_drive_pat_top.patsel1_high_q[2] ),
    .S(_02065_),
    .X(_02070_));
 sky130_fd_sc_hd__and2_1 _18917_ (.A(_02049_),
    .B(_02070_),
    .X(_02071_));
 sky130_fd_sc_hd__clkbuf_1 _18918_ (.A(_02071_),
    .X(_00722_));
 sky130_fd_sc_hd__buf_2 _18919_ (.A(_02048_),
    .X(_02072_));
 sky130_fd_sc_hd__mux2_1 _18920_ (.A0(_01669_),
    .A1(\wfg_drive_pat_top.patsel1_high_q[3] ),
    .S(_02065_),
    .X(_02073_));
 sky130_fd_sc_hd__and2_1 _18921_ (.A(_02072_),
    .B(_02073_),
    .X(_02074_));
 sky130_fd_sc_hd__clkbuf_1 _18922_ (.A(_02074_),
    .X(_00723_));
 sky130_fd_sc_hd__mux2_1 _18923_ (.A0(_01672_),
    .A1(\wfg_drive_pat_top.patsel1_high_q[4] ),
    .S(_02065_),
    .X(_02075_));
 sky130_fd_sc_hd__and2_1 _18924_ (.A(_02072_),
    .B(_02075_),
    .X(_02076_));
 sky130_fd_sc_hd__clkbuf_1 _18925_ (.A(_02076_),
    .X(_00724_));
 sky130_fd_sc_hd__mux2_1 _18926_ (.A0(_01675_),
    .A1(\wfg_drive_pat_top.patsel1_high_q[5] ),
    .S(_02065_),
    .X(_02077_));
 sky130_fd_sc_hd__and2_1 _18927_ (.A(_02072_),
    .B(_02077_),
    .X(_02078_));
 sky130_fd_sc_hd__clkbuf_1 _18928_ (.A(_02078_),
    .X(_00725_));
 sky130_fd_sc_hd__mux2_1 _18929_ (.A0(_01679_),
    .A1(\wfg_drive_pat_top.patsel1_high_q[6] ),
    .S(_02065_),
    .X(_02079_));
 sky130_fd_sc_hd__and2_1 _18930_ (.A(_02072_),
    .B(_02079_),
    .X(_02080_));
 sky130_fd_sc_hd__clkbuf_1 _18931_ (.A(_02080_),
    .X(_00726_));
 sky130_fd_sc_hd__mux2_1 _18932_ (.A0(_01682_),
    .A1(\wfg_drive_pat_top.patsel1_high_q[7] ),
    .S(_02065_),
    .X(_02081_));
 sky130_fd_sc_hd__and2_1 _18933_ (.A(_02072_),
    .B(_02081_),
    .X(_02082_));
 sky130_fd_sc_hd__clkbuf_1 _18934_ (.A(_02082_),
    .X(_00727_));
 sky130_fd_sc_hd__mux2_1 _18935_ (.A0(_01601_),
    .A1(\wfg_drive_pat_top.patsel1_high_q[8] ),
    .S(_02065_),
    .X(_02083_));
 sky130_fd_sc_hd__and2_1 _18936_ (.A(_02072_),
    .B(_02083_),
    .X(_02084_));
 sky130_fd_sc_hd__clkbuf_1 _18937_ (.A(_02084_),
    .X(_00728_));
 sky130_fd_sc_hd__mux2_1 _18938_ (.A0(_01620_),
    .A1(\wfg_drive_pat_top.patsel1_high_q[9] ),
    .S(_02065_),
    .X(_02085_));
 sky130_fd_sc_hd__and2_1 _18939_ (.A(_02072_),
    .B(_02085_),
    .X(_02086_));
 sky130_fd_sc_hd__clkbuf_1 _18940_ (.A(_02086_),
    .X(_00729_));
 sky130_fd_sc_hd__buf_4 _18941_ (.A(_02064_),
    .X(_02087_));
 sky130_fd_sc_hd__mux2_1 _18942_ (.A0(_01624_),
    .A1(\wfg_drive_pat_top.patsel1_high_q[10] ),
    .S(_02087_),
    .X(_02088_));
 sky130_fd_sc_hd__and2_1 _18943_ (.A(_02072_),
    .B(_02088_),
    .X(_02089_));
 sky130_fd_sc_hd__clkbuf_1 _18944_ (.A(_02089_),
    .X(_00730_));
 sky130_fd_sc_hd__mux2_1 _18945_ (.A0(_01627_),
    .A1(\wfg_drive_pat_top.patsel1_high_q[11] ),
    .S(_02087_),
    .X(_02090_));
 sky130_fd_sc_hd__and2_1 _18946_ (.A(_02072_),
    .B(_02090_),
    .X(_02091_));
 sky130_fd_sc_hd__clkbuf_1 _18947_ (.A(_02091_),
    .X(_00731_));
 sky130_fd_sc_hd__mux2_1 _18948_ (.A0(_01630_),
    .A1(\wfg_drive_pat_top.patsel1_high_q[12] ),
    .S(_02087_),
    .X(_02092_));
 sky130_fd_sc_hd__and2_1 _18949_ (.A(_02072_),
    .B(_02092_),
    .X(_02093_));
 sky130_fd_sc_hd__clkbuf_1 _18950_ (.A(_02093_),
    .X(_00732_));
 sky130_fd_sc_hd__buf_2 _18951_ (.A(_02048_),
    .X(_02094_));
 sky130_fd_sc_hd__mux2_1 _18952_ (.A0(_01633_),
    .A1(\wfg_drive_pat_top.patsel1_high_q[13] ),
    .S(_02087_),
    .X(_02095_));
 sky130_fd_sc_hd__and2_1 _18953_ (.A(_02094_),
    .B(_02095_),
    .X(_02096_));
 sky130_fd_sc_hd__clkbuf_1 _18954_ (.A(_02096_),
    .X(_00733_));
 sky130_fd_sc_hd__mux2_1 _18955_ (.A0(_01636_),
    .A1(\wfg_drive_pat_top.patsel1_high_q[14] ),
    .S(_02087_),
    .X(_02097_));
 sky130_fd_sc_hd__and2_1 _18956_ (.A(_02094_),
    .B(_02097_),
    .X(_02098_));
 sky130_fd_sc_hd__clkbuf_1 _18957_ (.A(_02098_),
    .X(_00734_));
 sky130_fd_sc_hd__mux2_1 _18958_ (.A0(_01639_),
    .A1(\wfg_drive_pat_top.patsel1_high_q[15] ),
    .S(_02087_),
    .X(_02099_));
 sky130_fd_sc_hd__and2_1 _18959_ (.A(_02094_),
    .B(_02099_),
    .X(_02100_));
 sky130_fd_sc_hd__clkbuf_1 _18960_ (.A(_02100_),
    .X(_00735_));
 sky130_fd_sc_hd__mux2_1 _18961_ (.A0(net73),
    .A1(\wfg_drive_pat_top.patsel1_high_q[16] ),
    .S(_02087_),
    .X(_02101_));
 sky130_fd_sc_hd__and2_1 _18962_ (.A(_02094_),
    .B(_02101_),
    .X(_02102_));
 sky130_fd_sc_hd__clkbuf_1 _18963_ (.A(_02102_),
    .X(_00736_));
 sky130_fd_sc_hd__mux2_1 _18964_ (.A0(net74),
    .A1(\wfg_drive_pat_top.patsel1_high_q[17] ),
    .S(_02087_),
    .X(_02103_));
 sky130_fd_sc_hd__and2_1 _18965_ (.A(_02094_),
    .B(_02103_),
    .X(_02104_));
 sky130_fd_sc_hd__clkbuf_1 _18966_ (.A(_02104_),
    .X(_00737_));
 sky130_fd_sc_hd__mux2_1 _18967_ (.A0(net75),
    .A1(\wfg_drive_pat_top.patsel1_high_q[18] ),
    .S(_02087_),
    .X(_02105_));
 sky130_fd_sc_hd__and2_1 _18968_ (.A(_02094_),
    .B(_02105_),
    .X(_02106_));
 sky130_fd_sc_hd__clkbuf_1 _18969_ (.A(_02106_),
    .X(_00738_));
 sky130_fd_sc_hd__mux2_1 _18970_ (.A0(net76),
    .A1(\wfg_drive_pat_top.patsel1_high_q[19] ),
    .S(_02087_),
    .X(_02107_));
 sky130_fd_sc_hd__and2_1 _18971_ (.A(_02094_),
    .B(_02107_),
    .X(_02108_));
 sky130_fd_sc_hd__clkbuf_1 _18972_ (.A(_02108_),
    .X(_00739_));
 sky130_fd_sc_hd__buf_4 _18973_ (.A(_02064_),
    .X(_02109_));
 sky130_fd_sc_hd__mux2_1 _18974_ (.A0(net78),
    .A1(\wfg_drive_pat_top.patsel1_high_q[20] ),
    .S(_02109_),
    .X(_02110_));
 sky130_fd_sc_hd__and2_1 _18975_ (.A(_02094_),
    .B(_02110_),
    .X(_02111_));
 sky130_fd_sc_hd__clkbuf_1 _18976_ (.A(_02111_),
    .X(_00740_));
 sky130_fd_sc_hd__mux2_1 _18977_ (.A0(net79),
    .A1(\wfg_drive_pat_top.patsel1_high_q[21] ),
    .S(_02109_),
    .X(_02112_));
 sky130_fd_sc_hd__and2_1 _18978_ (.A(_02094_),
    .B(_02112_),
    .X(_02113_));
 sky130_fd_sc_hd__clkbuf_1 _18979_ (.A(_02113_),
    .X(_00741_));
 sky130_fd_sc_hd__mux2_1 _18980_ (.A0(net80),
    .A1(\wfg_drive_pat_top.patsel1_high_q[22] ),
    .S(_02109_),
    .X(_02114_));
 sky130_fd_sc_hd__and2_1 _18981_ (.A(_02094_),
    .B(_02114_),
    .X(_02115_));
 sky130_fd_sc_hd__clkbuf_1 _18982_ (.A(_02115_),
    .X(_00742_));
 sky130_fd_sc_hd__buf_4 _18983_ (.A(_02048_),
    .X(_02116_));
 sky130_fd_sc_hd__mux2_1 _18984_ (.A0(net81),
    .A1(\wfg_drive_pat_top.patsel1_high_q[23] ),
    .S(_02109_),
    .X(_02117_));
 sky130_fd_sc_hd__and2_1 _18985_ (.A(_02116_),
    .B(_02117_),
    .X(_02118_));
 sky130_fd_sc_hd__clkbuf_1 _18986_ (.A(_02118_),
    .X(_00743_));
 sky130_fd_sc_hd__mux2_1 _18987_ (.A0(net82),
    .A1(\wfg_drive_pat_top.patsel1_high_q[24] ),
    .S(_02109_),
    .X(_02119_));
 sky130_fd_sc_hd__and2_1 _18988_ (.A(_02116_),
    .B(_02119_),
    .X(_02120_));
 sky130_fd_sc_hd__clkbuf_1 _18989_ (.A(_02120_),
    .X(_00744_));
 sky130_fd_sc_hd__mux2_1 _18990_ (.A0(net83),
    .A1(\wfg_drive_pat_top.patsel1_high_q[25] ),
    .S(_02109_),
    .X(_02121_));
 sky130_fd_sc_hd__and2_1 _18991_ (.A(_02116_),
    .B(_02121_),
    .X(_02122_));
 sky130_fd_sc_hd__clkbuf_1 _18992_ (.A(_02122_),
    .X(_00745_));
 sky130_fd_sc_hd__mux2_1 _18993_ (.A0(net84),
    .A1(\wfg_drive_pat_top.patsel1_high_q[26] ),
    .S(_02109_),
    .X(_02123_));
 sky130_fd_sc_hd__and2_1 _18994_ (.A(_02116_),
    .B(_02123_),
    .X(_02124_));
 sky130_fd_sc_hd__clkbuf_1 _18995_ (.A(_02124_),
    .X(_00746_));
 sky130_fd_sc_hd__mux2_1 _18996_ (.A0(net85),
    .A1(\wfg_drive_pat_top.patsel1_high_q[27] ),
    .S(_02109_),
    .X(_02125_));
 sky130_fd_sc_hd__and2_1 _18997_ (.A(_02116_),
    .B(_02125_),
    .X(_02126_));
 sky130_fd_sc_hd__clkbuf_1 _18998_ (.A(_02126_),
    .X(_00747_));
 sky130_fd_sc_hd__mux2_1 _18999_ (.A0(net86),
    .A1(\wfg_drive_pat_top.patsel1_high_q[28] ),
    .S(_02109_),
    .X(_02127_));
 sky130_fd_sc_hd__and2_1 _19000_ (.A(_02116_),
    .B(_02127_),
    .X(_02128_));
 sky130_fd_sc_hd__clkbuf_1 _19001_ (.A(_02128_),
    .X(_00748_));
 sky130_fd_sc_hd__mux2_1 _19002_ (.A0(net87),
    .A1(\wfg_drive_pat_top.patsel1_high_q[29] ),
    .S(_02109_),
    .X(_02129_));
 sky130_fd_sc_hd__and2_1 _19003_ (.A(_02116_),
    .B(_02129_),
    .X(_02130_));
 sky130_fd_sc_hd__clkbuf_1 _19004_ (.A(_02130_),
    .X(_00749_));
 sky130_fd_sc_hd__mux2_1 _19005_ (.A0(net89),
    .A1(\wfg_drive_pat_top.patsel1_high_q[30] ),
    .S(_02064_),
    .X(_02131_));
 sky130_fd_sc_hd__and2_1 _19006_ (.A(_02116_),
    .B(_02131_),
    .X(_02132_));
 sky130_fd_sc_hd__clkbuf_1 _19007_ (.A(_02132_),
    .X(_00750_));
 sky130_fd_sc_hd__mux2_1 _19008_ (.A0(net90),
    .A1(\wfg_drive_pat_top.patsel1_high_q[31] ),
    .S(_02064_),
    .X(_02133_));
 sky130_fd_sc_hd__and2_1 _19009_ (.A(_02116_),
    .B(_02133_),
    .X(_02134_));
 sky130_fd_sc_hd__clkbuf_1 _19010_ (.A(_02134_),
    .X(_00751_));
 sky130_fd_sc_hd__inv_2 _19011_ (.A(_01749_),
    .Y(_00143_));
 sky130_fd_sc_hd__inv_2 _19012_ (.A(_01749_),
    .Y(_00144_));
 sky130_fd_sc_hd__inv_2 _19013_ (.A(_01749_),
    .Y(_00145_));
 sky130_fd_sc_hd__inv_2 _19014_ (.A(_01749_),
    .Y(_00146_));
 sky130_fd_sc_hd__inv_2 _19015_ (.A(_01749_),
    .Y(_00147_));
 sky130_fd_sc_hd__inv_2 _19016_ (.A(_01749_),
    .Y(_00148_));
 sky130_fd_sc_hd__inv_2 _19017_ (.A(_01749_),
    .Y(_00149_));
 sky130_fd_sc_hd__inv_2 _19018_ (.A(_01749_),
    .Y(_00150_));
 sky130_fd_sc_hd__buf_4 _19019_ (.A(_01597_),
    .X(_02135_));
 sky130_fd_sc_hd__inv_2 _19020_ (.A(_02135_),
    .Y(_00151_));
 sky130_fd_sc_hd__inv_2 _19021_ (.A(_02135_),
    .Y(_00152_));
 sky130_fd_sc_hd__inv_2 _19022_ (.A(_02135_),
    .Y(_00153_));
 sky130_fd_sc_hd__inv_2 _19023_ (.A(_02135_),
    .Y(_00154_));
 sky130_fd_sc_hd__inv_2 _19024_ (.A(_02135_),
    .Y(_00155_));
 sky130_fd_sc_hd__inv_2 _19025_ (.A(_02135_),
    .Y(_00156_));
 sky130_fd_sc_hd__inv_2 _19026_ (.A(_02135_),
    .Y(_00157_));
 sky130_fd_sc_hd__inv_2 _19027_ (.A(_02135_),
    .Y(_00158_));
 sky130_fd_sc_hd__or3_4 _19028_ (.A(net59),
    .B(_01441_),
    .C(_01424_),
    .X(_02136_));
 sky130_fd_sc_hd__nor2_2 _19029_ (.A(_02136_),
    .B(_01686_),
    .Y(_02137_));
 sky130_fd_sc_hd__and3b_1 _19030_ (.A_N(\wfg_stim_sine_top.wbs_ack_o ),
    .B(_01697_),
    .C(_02137_),
    .X(_02138_));
 sky130_fd_sc_hd__clkbuf_1 _19031_ (.A(_02138_),
    .X(_00752_));
 sky130_fd_sc_hd__inv_2 _19032_ (.A(_02135_),
    .Y(_00159_));
 sky130_fd_sc_hd__inv_2 _19033_ (.A(_02135_),
    .Y(_00160_));
 sky130_fd_sc_hd__clkbuf_8 _19034_ (.A(_01597_),
    .X(_02139_));
 sky130_fd_sc_hd__inv_2 _19035_ (.A(_02139_),
    .Y(_00161_));
 sky130_fd_sc_hd__inv_2 _19036_ (.A(_02139_),
    .Y(_00162_));
 sky130_fd_sc_hd__inv_2 _19037_ (.A(_02139_),
    .Y(_00163_));
 sky130_fd_sc_hd__inv_2 _19038_ (.A(_02139_),
    .Y(_00164_));
 sky130_fd_sc_hd__inv_2 _19039_ (.A(_02139_),
    .Y(_00165_));
 sky130_fd_sc_hd__inv_2 _19040_ (.A(_02139_),
    .Y(_00166_));
 sky130_fd_sc_hd__inv_2 _19041_ (.A(_02139_),
    .Y(_00167_));
 sky130_fd_sc_hd__inv_2 _19042_ (.A(_02139_),
    .Y(_00168_));
 sky130_fd_sc_hd__mux2_1 _19043_ (.A0(\wfg_subcore_top.wfg_subcore.temp_subcycle ),
    .A1(\wfg_subcore_top.wfg_subcore.subcycle_dly ),
    .S(_01590_),
    .X(_02140_));
 sky130_fd_sc_hd__clkbuf_1 _19044_ (.A(_02140_),
    .X(_00763_));
 sky130_fd_sc_hd__mux2_1 _19045_ (.A0(\wfg_subcore_top.wfg_subcore.temp_sync ),
    .A1(\wfg_subcore_top.wfg_subcore.sync_dly ),
    .S(_01590_),
    .X(_02141_));
 sky130_fd_sc_hd__clkbuf_1 _19046_ (.A(_02141_),
    .X(_00764_));
 sky130_fd_sc_hd__inv_2 _19047_ (.A(_02139_),
    .Y(_00169_));
 sky130_fd_sc_hd__inv_2 _19048_ (.A(_02139_),
    .Y(_00170_));
 sky130_fd_sc_hd__buf_6 _19049_ (.A(_01590_),
    .X(_02142_));
 sky130_fd_sc_hd__buf_4 _19050_ (.A(_02142_),
    .X(_02143_));
 sky130_fd_sc_hd__inv_2 _19051_ (.A(_02143_),
    .Y(_00171_));
 sky130_fd_sc_hd__inv_2 _19052_ (.A(_02143_),
    .Y(_00172_));
 sky130_fd_sc_hd__inv_2 _19053_ (.A(_02143_),
    .Y(_00173_));
 sky130_fd_sc_hd__inv_2 _19054_ (.A(_02143_),
    .Y(_00174_));
 sky130_fd_sc_hd__inv_2 _19055_ (.A(_02143_),
    .Y(_00175_));
 sky130_fd_sc_hd__inv_2 _19056_ (.A(_02143_),
    .Y(_00176_));
 sky130_fd_sc_hd__and2_1 _19057_ (.A(_01706_),
    .B(_02137_),
    .X(_02144_));
 sky130_fd_sc_hd__buf_2 _19058_ (.A(_02144_),
    .X(_02145_));
 sky130_fd_sc_hd__buf_2 _19059_ (.A(_02145_),
    .X(_02146_));
 sky130_fd_sc_hd__or3b_1 _19060_ (.A(net59),
    .B(_01424_),
    .C_N(_01885_),
    .X(_02147_));
 sky130_fd_sc_hd__o211a_1 _19061_ (.A1(net55),
    .A2(net58),
    .B1(_01426_),
    .C1(_01755_),
    .X(_02148_));
 sky130_fd_sc_hd__inv_2 _19062_ (.A(_01604_),
    .Y(_02149_));
 sky130_fd_sc_hd__or2_1 _19063_ (.A(_01424_),
    .B(_01425_),
    .X(_02150_));
 sky130_fd_sc_hd__nor2_1 _19064_ (.A(_02150_),
    .B(_01756_),
    .Y(_02151_));
 sky130_fd_sc_hd__a32o_1 _19065_ (.A1(\wfg_stim_sine_top.inc_val_q[0] ),
    .A2(_01427_),
    .A3(_02149_),
    .B1(_02151_),
    .B2(\wfg_stim_sine_top.offset_val_q[0] ),
    .X(_02152_));
 sky130_fd_sc_hd__inv_2 _19066_ (.A(_07043_),
    .Y(_02153_));
 sky130_fd_sc_hd__o31ai_1 _19067_ (.A1(_02153_),
    .A2(_02150_),
    .A3(_01763_),
    .B1(_02148_),
    .Y(_02154_));
 sky130_fd_sc_hd__o22a_1 _19068_ (.A1(\wfg_stim_sine_top.ctrl_en_q ),
    .A2(_02148_),
    .B1(_02152_),
    .B2(_02154_),
    .X(_02155_));
 sky130_fd_sc_hd__or4_1 _19069_ (.A(_02147_),
    .B(_01686_),
    .C(_01713_),
    .D(_02155_),
    .X(_02156_));
 sky130_fd_sc_hd__buf_2 _19070_ (.A(_01730_),
    .X(_02157_));
 sky130_fd_sc_hd__o211a_1 _19071_ (.A1(\wfg_stim_sine_top.wbs_dat_o[0] ),
    .A2(_02146_),
    .B1(_02156_),
    .C1(_02157_),
    .X(_00773_));
 sky130_fd_sc_hd__nor2_4 _19072_ (.A(_02136_),
    .B(_01756_),
    .Y(_02158_));
 sky130_fd_sc_hd__buf_2 _19073_ (.A(_02158_),
    .X(_02159_));
 sky130_fd_sc_hd__nor2_2 _19074_ (.A(_02136_),
    .B(_01763_),
    .Y(_02160_));
 sky130_fd_sc_hd__buf_2 _19075_ (.A(_02160_),
    .X(_02161_));
 sky130_fd_sc_hd__nor2_2 _19076_ (.A(_02136_),
    .B(_01959_),
    .Y(_02162_));
 sky130_fd_sc_hd__buf_2 _19077_ (.A(_02162_),
    .X(_02163_));
 sky130_fd_sc_hd__a22o_1 _19078_ (.A1(_07044_),
    .A2(_02161_),
    .B1(_02163_),
    .B2(\wfg_stim_sine_top.inc_val_q[1] ),
    .X(_02164_));
 sky130_fd_sc_hd__nand2_4 _19079_ (.A(_01706_),
    .B(_02137_),
    .Y(_02165_));
 sky130_fd_sc_hd__buf_2 _19080_ (.A(_02165_),
    .X(_02166_));
 sky130_fd_sc_hd__a211o_1 _19081_ (.A1(\wfg_stim_sine_top.offset_val_q[1] ),
    .A2(_02159_),
    .B1(_02164_),
    .C1(_02166_),
    .X(_02167_));
 sky130_fd_sc_hd__o211a_1 _19082_ (.A1(\wfg_stim_sine_top.wbs_dat_o[1] ),
    .A2(_02146_),
    .B1(_02167_),
    .C1(_02157_),
    .X(_00774_));
 sky130_fd_sc_hd__a22o_1 _19083_ (.A1(\wfg_stim_sine_top.offset_val_q[2] ),
    .A2(_02158_),
    .B1(_02163_),
    .B2(\wfg_stim_sine_top.inc_val_q[2] ),
    .X(_02168_));
 sky130_fd_sc_hd__a211o_1 _19084_ (.A1(_06605_),
    .A2(_02161_),
    .B1(_02165_),
    .C1(_02168_),
    .X(_02169_));
 sky130_fd_sc_hd__o211a_1 _19085_ (.A1(\wfg_stim_sine_top.wbs_dat_o[2] ),
    .A2(_02146_),
    .B1(_02169_),
    .C1(_02157_),
    .X(_00775_));
 sky130_fd_sc_hd__a22o_1 _19086_ (.A1(_07206_),
    .A2(_02161_),
    .B1(_02163_),
    .B2(\wfg_stim_sine_top.inc_val_q[3] ),
    .X(_02170_));
 sky130_fd_sc_hd__a211o_1 _19087_ (.A1(\wfg_stim_sine_top.offset_val_q[3] ),
    .A2(_02159_),
    .B1(_02170_),
    .C1(_02166_),
    .X(_02171_));
 sky130_fd_sc_hd__o211a_1 _19088_ (.A1(\wfg_stim_sine_top.wbs_dat_o[3] ),
    .A2(_02146_),
    .B1(_02171_),
    .C1(_02157_),
    .X(_00776_));
 sky130_fd_sc_hd__a22o_1 _19089_ (.A1(\wfg_stim_sine_top.offset_val_q[4] ),
    .A2(_02158_),
    .B1(_02163_),
    .B2(\wfg_stim_sine_top.inc_val_q[4] ),
    .X(_02172_));
 sky130_fd_sc_hd__a211o_1 _19090_ (.A1(_06551_),
    .A2(_02161_),
    .B1(_02165_),
    .C1(_02172_),
    .X(_02173_));
 sky130_fd_sc_hd__o211a_1 _19091_ (.A1(\wfg_stim_sine_top.wbs_dat_o[4] ),
    .A2(_02146_),
    .B1(_02173_),
    .C1(_02157_),
    .X(_00777_));
 sky130_fd_sc_hd__a22o_1 _19092_ (.A1(\wfg_stim_sine_top.offset_val_q[5] ),
    .A2(_02158_),
    .B1(_02163_),
    .B2(\wfg_stim_sine_top.inc_val_q[5] ),
    .X(_02174_));
 sky130_fd_sc_hd__a211o_1 _19093_ (.A1(_06549_),
    .A2(_02161_),
    .B1(_02165_),
    .C1(_02174_),
    .X(_02175_));
 sky130_fd_sc_hd__o211a_1 _19094_ (.A1(\wfg_stim_sine_top.wbs_dat_o[5] ),
    .A2(_02146_),
    .B1(_02175_),
    .C1(_02157_),
    .X(_00778_));
 sky130_fd_sc_hd__a22o_1 _19095_ (.A1(_06547_),
    .A2(_02161_),
    .B1(_02163_),
    .B2(\wfg_stim_sine_top.inc_val_q[6] ),
    .X(_02176_));
 sky130_fd_sc_hd__a211o_1 _19096_ (.A1(\wfg_stim_sine_top.offset_val_q[6] ),
    .A2(_02159_),
    .B1(_02176_),
    .C1(_02166_),
    .X(_02177_));
 sky130_fd_sc_hd__o211a_1 _19097_ (.A1(\wfg_stim_sine_top.wbs_dat_o[6] ),
    .A2(_02146_),
    .B1(_02177_),
    .C1(_02157_),
    .X(_00779_));
 sky130_fd_sc_hd__a22o_1 _19098_ (.A1(\wfg_stim_sine_top.offset_val_q[7] ),
    .A2(_02158_),
    .B1(_02163_),
    .B2(\wfg_stim_sine_top.inc_val_q[7] ),
    .X(_02178_));
 sky130_fd_sc_hd__a211o_1 _19099_ (.A1(_06486_),
    .A2(_02161_),
    .B1(_02165_),
    .C1(_02178_),
    .X(_02179_));
 sky130_fd_sc_hd__o211a_1 _19100_ (.A1(\wfg_stim_sine_top.wbs_dat_o[7] ),
    .A2(_02146_),
    .B1(_02179_),
    .C1(_02157_),
    .X(_00780_));
 sky130_fd_sc_hd__a22o_1 _19101_ (.A1(_06725_),
    .A2(_02160_),
    .B1(_02162_),
    .B2(\wfg_stim_sine_top.inc_val_q[8] ),
    .X(_02180_));
 sky130_fd_sc_hd__a211o_1 _19102_ (.A1(\wfg_stim_sine_top.offset_val_q[8] ),
    .A2(_02159_),
    .B1(_02180_),
    .C1(_02166_),
    .X(_02181_));
 sky130_fd_sc_hd__o211a_1 _19103_ (.A1(\wfg_stim_sine_top.wbs_dat_o[8] ),
    .A2(_02146_),
    .B1(_02181_),
    .C1(_02157_),
    .X(_00781_));
 sky130_fd_sc_hd__a22o_1 _19104_ (.A1(\wfg_stim_sine_top.offset_val_q[9] ),
    .A2(_02158_),
    .B1(_02163_),
    .B2(\wfg_stim_sine_top.inc_val_q[9] ),
    .X(_02182_));
 sky130_fd_sc_hd__a211o_1 _19105_ (.A1(_06714_),
    .A2(_02161_),
    .B1(_02165_),
    .C1(_02182_),
    .X(_02183_));
 sky130_fd_sc_hd__o211a_1 _19106_ (.A1(\wfg_stim_sine_top.wbs_dat_o[9] ),
    .A2(_02146_),
    .B1(_02183_),
    .C1(_02157_),
    .X(_00782_));
 sky130_fd_sc_hd__a22o_1 _19107_ (.A1(_06451_),
    .A2(_02160_),
    .B1(_02162_),
    .B2(\wfg_stim_sine_top.inc_val_q[10] ),
    .X(_02184_));
 sky130_fd_sc_hd__a211o_1 _19108_ (.A1(\wfg_stim_sine_top.offset_val_q[10] ),
    .A2(_02159_),
    .B1(_02184_),
    .C1(_02166_),
    .X(_02185_));
 sky130_fd_sc_hd__clkbuf_4 _19109_ (.A(_01589_),
    .X(_02186_));
 sky130_fd_sc_hd__o211a_1 _19110_ (.A1(\wfg_stim_sine_top.wbs_dat_o[10] ),
    .A2(_02145_),
    .B1(_02185_),
    .C1(_02186_),
    .X(_00783_));
 sky130_fd_sc_hd__a22o_1 _19111_ (.A1(_06471_),
    .A2(_02160_),
    .B1(_02162_),
    .B2(\wfg_stim_sine_top.inc_val_q[11] ),
    .X(_02187_));
 sky130_fd_sc_hd__a211o_1 _19112_ (.A1(\wfg_stim_sine_top.offset_val_q[11] ),
    .A2(_02159_),
    .B1(_02187_),
    .C1(_02166_),
    .X(_02188_));
 sky130_fd_sc_hd__o211a_1 _19113_ (.A1(\wfg_stim_sine_top.wbs_dat_o[11] ),
    .A2(_02145_),
    .B1(_02188_),
    .C1(_02186_),
    .X(_00784_));
 sky130_fd_sc_hd__a22o_1 _19114_ (.A1(_06474_),
    .A2(_02160_),
    .B1(_02162_),
    .B2(\wfg_stim_sine_top.inc_val_q[12] ),
    .X(_02189_));
 sky130_fd_sc_hd__a211o_1 _19115_ (.A1(\wfg_stim_sine_top.offset_val_q[12] ),
    .A2(_02159_),
    .B1(_02189_),
    .C1(_02166_),
    .X(_02190_));
 sky130_fd_sc_hd__o211a_1 _19116_ (.A1(\wfg_stim_sine_top.wbs_dat_o[12] ),
    .A2(_02145_),
    .B1(_02190_),
    .C1(_02186_),
    .X(_00785_));
 sky130_fd_sc_hd__a22o_1 _19117_ (.A1(\wfg_stim_sine_top.offset_val_q[13] ),
    .A2(_02158_),
    .B1(_02163_),
    .B2(\wfg_stim_sine_top.inc_val_q[13] ),
    .X(_02191_));
 sky130_fd_sc_hd__a211o_1 _19118_ (.A1(_06509_),
    .A2(_02161_),
    .B1(_02165_),
    .C1(_02191_),
    .X(_02192_));
 sky130_fd_sc_hd__o211a_1 _19119_ (.A1(\wfg_stim_sine_top.wbs_dat_o[13] ),
    .A2(_02145_),
    .B1(_02192_),
    .C1(_02186_),
    .X(_00786_));
 sky130_fd_sc_hd__a22o_1 _19120_ (.A1(\wfg_stim_sine_top.offset_val_q[14] ),
    .A2(_02158_),
    .B1(_02163_),
    .B2(\wfg_stim_sine_top.inc_val_q[14] ),
    .X(_02193_));
 sky130_fd_sc_hd__a211o_1 _19121_ (.A1(_06505_),
    .A2(_02161_),
    .B1(_02165_),
    .C1(_02193_),
    .X(_02194_));
 sky130_fd_sc_hd__o211a_1 _19122_ (.A1(\wfg_stim_sine_top.wbs_dat_o[14] ),
    .A2(_02145_),
    .B1(_02194_),
    .C1(_02186_),
    .X(_00787_));
 sky130_fd_sc_hd__a22o_1 _19123_ (.A1(_08081_),
    .A2(_02160_),
    .B1(_02162_),
    .B2(\wfg_stim_sine_top.inc_val_q[15] ),
    .X(_02195_));
 sky130_fd_sc_hd__a211o_1 _19124_ (.A1(\wfg_stim_sine_top.offset_val_q[15] ),
    .A2(_02159_),
    .B1(_02195_),
    .C1(_02166_),
    .X(_02196_));
 sky130_fd_sc_hd__o211a_1 _19125_ (.A1(\wfg_stim_sine_top.wbs_dat_o[15] ),
    .A2(_02145_),
    .B1(_02196_),
    .C1(_02186_),
    .X(_00788_));
 sky130_fd_sc_hd__a21o_1 _19126_ (.A1(\wfg_stim_sine_top.offset_val_q[16] ),
    .A2(_02159_),
    .B1(_02166_),
    .X(_02197_));
 sky130_fd_sc_hd__o211a_1 _19127_ (.A1(\wfg_stim_sine_top.wbs_dat_o[16] ),
    .A2(_02145_),
    .B1(_02197_),
    .C1(_02186_),
    .X(_00789_));
 sky130_fd_sc_hd__a21o_1 _19128_ (.A1(\wfg_stim_sine_top.offset_val_q[17] ),
    .A2(_02159_),
    .B1(_02166_),
    .X(_02198_));
 sky130_fd_sc_hd__o211a_1 _19129_ (.A1(\wfg_stim_sine_top.wbs_dat_o[17] ),
    .A2(_02145_),
    .B1(_02198_),
    .C1(_02186_),
    .X(_00790_));
 sky130_fd_sc_hd__or3_1 _19130_ (.A(_01959_),
    .B(_01605_),
    .C(_01712_),
    .X(_02199_));
 sky130_fd_sc_hd__clkbuf_2 _19131_ (.A(_02199_),
    .X(_02200_));
 sky130_fd_sc_hd__buf_2 _19132_ (.A(_02200_),
    .X(_02201_));
 sky130_fd_sc_hd__and2_1 _19133_ (.A(net100),
    .B(net65),
    .X(_02202_));
 sky130_fd_sc_hd__clkbuf_4 _19134_ (.A(_02202_),
    .X(_02203_));
 sky130_fd_sc_hd__and3_1 _19135_ (.A(_02149_),
    .B(_02203_),
    .C(_01696_),
    .X(_02204_));
 sky130_fd_sc_hd__clkbuf_2 _19136_ (.A(_02204_),
    .X(_02205_));
 sky130_fd_sc_hd__or2_1 _19137_ (.A(\wfg_subcore_top.cfg_subcycle_q[8] ),
    .B(_02205_),
    .X(_02206_));
 sky130_fd_sc_hd__o211a_1 _19138_ (.A1(_01601_),
    .A2(_02201_),
    .B1(_02206_),
    .C1(_02186_),
    .X(_00791_));
 sky130_fd_sc_hd__or2_1 _19139_ (.A(\wfg_subcore_top.cfg_subcycle_q[9] ),
    .B(_02205_),
    .X(_02207_));
 sky130_fd_sc_hd__o211a_1 _19140_ (.A1(_01620_),
    .A2(_02201_),
    .B1(_02207_),
    .C1(_02186_),
    .X(_00792_));
 sky130_fd_sc_hd__or2_1 _19141_ (.A(\wfg_subcore_top.cfg_subcycle_q[10] ),
    .B(_02205_),
    .X(_02208_));
 sky130_fd_sc_hd__buf_2 _19142_ (.A(_01589_),
    .X(_02209_));
 sky130_fd_sc_hd__o211a_1 _19143_ (.A1(_01624_),
    .A2(_02201_),
    .B1(_02208_),
    .C1(_02209_),
    .X(_00793_));
 sky130_fd_sc_hd__or2_1 _19144_ (.A(\wfg_subcore_top.cfg_subcycle_q[11] ),
    .B(_02205_),
    .X(_02210_));
 sky130_fd_sc_hd__o211a_1 _19145_ (.A1(_01627_),
    .A2(_02201_),
    .B1(_02210_),
    .C1(_02209_),
    .X(_00794_));
 sky130_fd_sc_hd__or2_1 _19146_ (.A(\wfg_subcore_top.cfg_subcycle_q[12] ),
    .B(_02205_),
    .X(_02211_));
 sky130_fd_sc_hd__o211a_1 _19147_ (.A1(_01630_),
    .A2(_02201_),
    .B1(_02211_),
    .C1(_02209_),
    .X(_00795_));
 sky130_fd_sc_hd__or2_1 _19148_ (.A(\wfg_subcore_top.cfg_subcycle_q[13] ),
    .B(_02205_),
    .X(_02212_));
 sky130_fd_sc_hd__o211a_1 _19149_ (.A1(_01633_),
    .A2(_02201_),
    .B1(_02212_),
    .C1(_02209_),
    .X(_00796_));
 sky130_fd_sc_hd__or2_1 _19150_ (.A(\wfg_subcore_top.cfg_subcycle_q[14] ),
    .B(_02205_),
    .X(_02213_));
 sky130_fd_sc_hd__o211a_1 _19151_ (.A1(_01636_),
    .A2(_02201_),
    .B1(_02213_),
    .C1(_02209_),
    .X(_00797_));
 sky130_fd_sc_hd__or2_1 _19152_ (.A(\wfg_subcore_top.cfg_subcycle_q[15] ),
    .B(_02205_),
    .X(_02214_));
 sky130_fd_sc_hd__o211a_1 _19153_ (.A1(_01639_),
    .A2(_02201_),
    .B1(_02214_),
    .C1(_02209_),
    .X(_00798_));
 sky130_fd_sc_hd__or2_1 _19154_ (.A(\wfg_subcore_top.cfg_subcycle_q[16] ),
    .B(_02205_),
    .X(_02215_));
 sky130_fd_sc_hd__o211a_1 _19155_ (.A1(net73),
    .A2(_02201_),
    .B1(_02215_),
    .C1(_02209_),
    .X(_00799_));
 sky130_fd_sc_hd__or2_1 _19156_ (.A(\wfg_subcore_top.cfg_subcycle_q[17] ),
    .B(_02205_),
    .X(_02216_));
 sky130_fd_sc_hd__o211a_1 _19157_ (.A1(net74),
    .A2(_02201_),
    .B1(_02216_),
    .C1(_02209_),
    .X(_00800_));
 sky130_fd_sc_hd__clkbuf_4 _19158_ (.A(_02200_),
    .X(_02217_));
 sky130_fd_sc_hd__buf_2 _19159_ (.A(_02204_),
    .X(_02218_));
 sky130_fd_sc_hd__or2_1 _19160_ (.A(\wfg_subcore_top.cfg_subcycle_q[18] ),
    .B(_02218_),
    .X(_02219_));
 sky130_fd_sc_hd__o211a_1 _19161_ (.A1(net75),
    .A2(_02217_),
    .B1(_02219_),
    .C1(_02209_),
    .X(_00801_));
 sky130_fd_sc_hd__or2_1 _19162_ (.A(\wfg_subcore_top.cfg_subcycle_q[19] ),
    .B(_02218_),
    .X(_02220_));
 sky130_fd_sc_hd__o211a_1 _19163_ (.A1(net76),
    .A2(_02217_),
    .B1(_02220_),
    .C1(_02209_),
    .X(_00802_));
 sky130_fd_sc_hd__or2_1 _19164_ (.A(\wfg_subcore_top.cfg_subcycle_q[20] ),
    .B(_02218_),
    .X(_02221_));
 sky130_fd_sc_hd__clkbuf_4 _19165_ (.A(_01589_),
    .X(_02222_));
 sky130_fd_sc_hd__o211a_1 _19166_ (.A1(net78),
    .A2(_02217_),
    .B1(_02221_),
    .C1(_02222_),
    .X(_00803_));
 sky130_fd_sc_hd__or2_1 _19167_ (.A(\wfg_subcore_top.cfg_subcycle_q[21] ),
    .B(_02218_),
    .X(_02223_));
 sky130_fd_sc_hd__o211a_1 _19168_ (.A1(net79),
    .A2(_02217_),
    .B1(_02223_),
    .C1(_02222_),
    .X(_00804_));
 sky130_fd_sc_hd__or2_1 _19169_ (.A(\wfg_subcore_top.cfg_subcycle_q[22] ),
    .B(_02218_),
    .X(_02224_));
 sky130_fd_sc_hd__o211a_1 _19170_ (.A1(net80),
    .A2(_02217_),
    .B1(_02224_),
    .C1(_02222_),
    .X(_00805_));
 sky130_fd_sc_hd__or2_1 _19171_ (.A(\wfg_subcore_top.cfg_subcycle_q[23] ),
    .B(_02218_),
    .X(_02225_));
 sky130_fd_sc_hd__o211a_1 _19172_ (.A1(net81),
    .A2(_02217_),
    .B1(_02225_),
    .C1(_02222_),
    .X(_00806_));
 sky130_fd_sc_hd__or2_1 _19173_ (.A(\wfg_subcore_top.cfg_sync_q[0] ),
    .B(_02218_),
    .X(_02226_));
 sky130_fd_sc_hd__o211a_1 _19174_ (.A1(_01660_),
    .A2(_02217_),
    .B1(_02226_),
    .C1(_02222_),
    .X(_00807_));
 sky130_fd_sc_hd__or2_1 _19175_ (.A(\wfg_subcore_top.cfg_sync_q[1] ),
    .B(_02218_),
    .X(_02227_));
 sky130_fd_sc_hd__o211a_1 _19176_ (.A1(_01663_),
    .A2(_02217_),
    .B1(_02227_),
    .C1(_02222_),
    .X(_00808_));
 sky130_fd_sc_hd__or2_1 _19177_ (.A(\wfg_subcore_top.cfg_sync_q[2] ),
    .B(_02218_),
    .X(_02228_));
 sky130_fd_sc_hd__o211a_1 _19178_ (.A1(_01666_),
    .A2(_02217_),
    .B1(_02228_),
    .C1(_02222_),
    .X(_00809_));
 sky130_fd_sc_hd__or2_1 _19179_ (.A(\wfg_subcore_top.cfg_sync_q[3] ),
    .B(_02218_),
    .X(_02229_));
 sky130_fd_sc_hd__o211a_1 _19180_ (.A1(_01669_),
    .A2(_02217_),
    .B1(_02229_),
    .C1(_02222_),
    .X(_00810_));
 sky130_fd_sc_hd__or2_1 _19181_ (.A(\wfg_subcore_top.cfg_sync_q[4] ),
    .B(_02204_),
    .X(_02230_));
 sky130_fd_sc_hd__o211a_1 _19182_ (.A1(_01672_),
    .A2(_02200_),
    .B1(_02230_),
    .C1(_02222_),
    .X(_00811_));
 sky130_fd_sc_hd__or2_1 _19183_ (.A(\wfg_subcore_top.cfg_sync_q[5] ),
    .B(_02204_),
    .X(_02231_));
 sky130_fd_sc_hd__o211a_1 _19184_ (.A1(_01675_),
    .A2(_02200_),
    .B1(_02231_),
    .C1(_02222_),
    .X(_00812_));
 sky130_fd_sc_hd__or2_1 _19185_ (.A(\wfg_subcore_top.cfg_sync_q[6] ),
    .B(_02204_),
    .X(_02232_));
 sky130_fd_sc_hd__clkbuf_4 _19186_ (.A(_01589_),
    .X(_02233_));
 sky130_fd_sc_hd__o211a_1 _19187_ (.A1(_01679_),
    .A2(_02200_),
    .B1(_02232_),
    .C1(_02233_),
    .X(_00813_));
 sky130_fd_sc_hd__nand2_1 _19188_ (.A(_09758_),
    .B(_02200_),
    .Y(_02234_));
 sky130_fd_sc_hd__o211a_1 _19189_ (.A1(_01682_),
    .A2(_02200_),
    .B1(_02234_),
    .C1(_02233_),
    .X(_00814_));
 sky130_fd_sc_hd__a31o_1 _19190_ (.A1(_02203_),
    .A2(_01709_),
    .A3(_01696_),
    .B1(\wfg_subcore_top.active_o ),
    .X(_02235_));
 sky130_fd_sc_hd__or4_1 _19191_ (.A(net66),
    .B(_01605_),
    .C(_01691_),
    .D(_01712_),
    .X(_02236_));
 sky130_fd_sc_hd__and3_1 _19192_ (.A(_01685_),
    .B(_02235_),
    .C(_02236_),
    .X(_02237_));
 sky130_fd_sc_hd__clkbuf_1 _19193_ (.A(_02237_),
    .X(_00815_));
 sky130_fd_sc_hd__or3_4 _19194_ (.A(net59),
    .B(_01431_),
    .C(_01441_),
    .X(_02238_));
 sky130_fd_sc_hd__nor2_2 _19195_ (.A(_02238_),
    .B(_01686_),
    .Y(_02239_));
 sky130_fd_sc_hd__and3b_1 _19196_ (.A_N(\wfg_drive_spi_top.wbs_ack_o ),
    .B(_01697_),
    .C(_02239_),
    .X(_02240_));
 sky130_fd_sc_hd__clkbuf_1 _19197_ (.A(_02240_),
    .X(_00816_));
 sky130_fd_sc_hd__and2_1 _19198_ (.A(_01706_),
    .B(_02239_),
    .X(_02241_));
 sky130_fd_sc_hd__clkbuf_2 _19199_ (.A(_02241_),
    .X(_02242_));
 sky130_fd_sc_hd__nor2_2 _19200_ (.A(_02238_),
    .B(_01761_),
    .Y(_02243_));
 sky130_fd_sc_hd__nand2_2 _19201_ (.A(_01706_),
    .B(_02239_),
    .Y(_02244_));
 sky130_fd_sc_hd__nor2_2 _19202_ (.A(_02238_),
    .B(_01763_),
    .Y(_02245_));
 sky130_fd_sc_hd__o21a_1 _19203_ (.A1(_02238_),
    .A2(_01709_),
    .B1(\wfg_drive_spi_top.ctrl_en_q ),
    .X(_02246_));
 sky130_fd_sc_hd__a21o_1 _19204_ (.A1(\wfg_drive_spi_top.clkcfg_div_q[0] ),
    .A2(_02245_),
    .B1(_02246_),
    .X(_02247_));
 sky130_fd_sc_hd__a211o_1 _19205_ (.A1(\wfg_drive_spi_top.cfg_cpol_q ),
    .A2(_02243_),
    .B1(_02244_),
    .C1(_02247_),
    .X(_02248_));
 sky130_fd_sc_hd__o211a_1 _19206_ (.A1(\wfg_drive_spi_top.wbs_dat_o[0] ),
    .A2(_02242_),
    .B1(_02248_),
    .C1(_02233_),
    .X(_00817_));
 sky130_fd_sc_hd__a221o_1 _19207_ (.A1(\wfg_drive_spi_top.clkcfg_div_q[1] ),
    .A2(_02245_),
    .B1(_02243_),
    .B2(\wfg_drive_spi_top.cfg_lsbfirst_q ),
    .C1(_02244_),
    .X(_02249_));
 sky130_fd_sc_hd__o211a_1 _19208_ (.A1(\wfg_drive_spi_top.wbs_dat_o[1] ),
    .A2(_02242_),
    .B1(_02249_),
    .C1(_02233_),
    .X(_00818_));
 sky130_fd_sc_hd__a221o_1 _19209_ (.A1(\wfg_drive_spi_top.clkcfg_div_q[2] ),
    .A2(_02245_),
    .B1(_02243_),
    .B2(\wfg_drive_spi_top.cfg_dff_q[2] ),
    .C1(_02244_),
    .X(_02250_));
 sky130_fd_sc_hd__o211a_1 _19210_ (.A1(\wfg_drive_spi_top.wbs_dat_o[2] ),
    .A2(_02242_),
    .B1(_02250_),
    .C1(_02233_),
    .X(_00819_));
 sky130_fd_sc_hd__a221o_1 _19211_ (.A1(\wfg_drive_spi_top.clkcfg_div_q[3] ),
    .A2(_02245_),
    .B1(_02243_),
    .B2(\wfg_drive_spi_top.cfg_dff_q[3] ),
    .C1(_02244_),
    .X(_02251_));
 sky130_fd_sc_hd__o211a_1 _19212_ (.A1(\wfg_drive_spi_top.wbs_dat_o[3] ),
    .A2(_02242_),
    .B1(_02251_),
    .C1(_02233_),
    .X(_00820_));
 sky130_fd_sc_hd__a221o_1 _19213_ (.A1(\wfg_drive_spi_top.clkcfg_div_q[4] ),
    .A2(_02245_),
    .B1(_02243_),
    .B2(\wfg_drive_spi_top.cfg_sspol_q ),
    .C1(_02244_),
    .X(_02252_));
 sky130_fd_sc_hd__o211a_1 _19214_ (.A1(\wfg_drive_spi_top.wbs_dat_o[4] ),
    .A2(_02242_),
    .B1(_02252_),
    .C1(_02233_),
    .X(_00821_));
 sky130_fd_sc_hd__a221o_1 _19215_ (.A1(\wfg_drive_spi_top.clkcfg_div_q[5] ),
    .A2(_02245_),
    .B1(_02243_),
    .B2(\wfg_drive_spi_top.cfg_core_sel_q ),
    .C1(_02244_),
    .X(_02253_));
 sky130_fd_sc_hd__o211a_1 _19216_ (.A1(\wfg_drive_spi_top.wbs_dat_o[5] ),
    .A2(_02242_),
    .B1(_02253_),
    .C1(_02233_),
    .X(_00822_));
 sky130_fd_sc_hd__nand2_1 _19217_ (.A(\wfg_drive_spi_top.wbs_dat_o[6] ),
    .B(_02244_),
    .Y(_02254_));
 sky130_fd_sc_hd__and4b_1 _19218_ (.A_N(_02238_),
    .B(_01959_),
    .C(_01691_),
    .D(_02242_),
    .X(_02255_));
 sky130_fd_sc_hd__nand2_1 _19219_ (.A(\wfg_drive_spi_top.clkcfg_div_q[6] ),
    .B(_02255_),
    .Y(_02256_));
 sky130_fd_sc_hd__a21oi_1 _19220_ (.A1(_02254_),
    .A2(_02256_),
    .B1(_01591_),
    .Y(_00823_));
 sky130_fd_sc_hd__nand2_1 _19221_ (.A(\wfg_drive_spi_top.wbs_dat_o[7] ),
    .B(_02244_),
    .Y(_02257_));
 sky130_fd_sc_hd__nand2_1 _19222_ (.A(\wfg_drive_spi_top.clkcfg_div_q[7] ),
    .B(_02255_),
    .Y(_02258_));
 sky130_fd_sc_hd__a21oi_1 _19223_ (.A1(_02257_),
    .A2(_02258_),
    .B1(_01591_),
    .Y(_00824_));
 sky130_fd_sc_hd__or2_2 _19224_ (.A(_01412_),
    .B(_01443_),
    .X(_02259_));
 sky130_fd_sc_hd__nor2_2 _19225_ (.A(_02259_),
    .B(_01686_),
    .Y(_02260_));
 sky130_fd_sc_hd__nand2_1 _19226_ (.A(_02203_),
    .B(_02260_),
    .Y(_02261_));
 sky130_fd_sc_hd__a31o_1 _19227_ (.A1(_02203_),
    .A2(_01709_),
    .A3(_02260_),
    .B1(\wfg_interconnect_top.ctrl_en_q ),
    .X(_02262_));
 sky130_fd_sc_hd__o311a_1 _19228_ (.A1(_01660_),
    .A2(_01691_),
    .A3(_02261_),
    .B1(_02262_),
    .C1(_01600_),
    .X(_00825_));
 sky130_fd_sc_hd__or2_1 _19229_ (.A(_01959_),
    .B(_02261_),
    .X(_02263_));
 sky130_fd_sc_hd__a21oi_1 _19230_ (.A1(_02743_),
    .A2(_02263_),
    .B1(_01591_),
    .Y(_02264_));
 sky130_fd_sc_hd__o21a_1 _19231_ (.A1(_01660_),
    .A2(_02263_),
    .B1(_02264_),
    .X(_00826_));
 sky130_fd_sc_hd__a21oi_1 _19232_ (.A1(_02706_),
    .A2(_02263_),
    .B1(_01591_),
    .Y(_02265_));
 sky130_fd_sc_hd__o21a_1 _19233_ (.A1(_01663_),
    .A2(_02263_),
    .B1(_02265_),
    .X(_00827_));
 sky130_fd_sc_hd__or2_1 _19234_ (.A(_01763_),
    .B(_02261_),
    .X(_02266_));
 sky130_fd_sc_hd__nor2_1 _19235_ (.A(_01763_),
    .B(_02261_),
    .Y(_02267_));
 sky130_fd_sc_hd__or2_1 _19236_ (.A(\wfg_interconnect_top.driver1_select_q[0] ),
    .B(_02267_),
    .X(_02268_));
 sky130_fd_sc_hd__o211a_1 _19237_ (.A1(_01660_),
    .A2(_02266_),
    .B1(_02268_),
    .C1(_02233_),
    .X(_00828_));
 sky130_fd_sc_hd__or2_1 _19238_ (.A(\wfg_interconnect_top.driver1_select_q[1] ),
    .B(_02267_),
    .X(_02269_));
 sky130_fd_sc_hd__o211a_1 _19239_ (.A1(_01663_),
    .A2(_02266_),
    .B1(_02269_),
    .C1(_02233_),
    .X(_00829_));
 sky130_fd_sc_hd__inv_2 _19240_ (.A(_02143_),
    .Y(_00177_));
 sky130_fd_sc_hd__inv_2 _19241_ (.A(_02143_),
    .Y(_00178_));
 sky130_fd_sc_hd__inv_2 _19242_ (.A(_02143_),
    .Y(_00179_));
 sky130_fd_sc_hd__inv_2 _19243_ (.A(_02143_),
    .Y(_00180_));
 sky130_fd_sc_hd__buf_4 _19244_ (.A(_02142_),
    .X(_02270_));
 sky130_fd_sc_hd__inv_2 _19245_ (.A(_02270_),
    .Y(_00181_));
 sky130_fd_sc_hd__inv_2 _19246_ (.A(_02270_),
    .Y(_00182_));
 sky130_fd_sc_hd__inv_2 _19247_ (.A(_02270_),
    .Y(_00183_));
 sky130_fd_sc_hd__inv_2 _19248_ (.A(_02270_),
    .Y(_00184_));
 sky130_fd_sc_hd__inv_2 _19249_ (.A(_02270_),
    .Y(_00185_));
 sky130_fd_sc_hd__inv_2 _19250_ (.A(_02270_),
    .Y(_00186_));
 sky130_fd_sc_hd__inv_2 _19251_ (.A(_02270_),
    .Y(_00187_));
 sky130_fd_sc_hd__inv_2 _19252_ (.A(_02270_),
    .Y(_00188_));
 sky130_fd_sc_hd__inv_2 _19253_ (.A(_02270_),
    .Y(_00189_));
 sky130_fd_sc_hd__inv_2 _19254_ (.A(_02270_),
    .Y(_00190_));
 sky130_fd_sc_hd__buf_6 _19255_ (.A(_02142_),
    .X(_02271_));
 sky130_fd_sc_hd__inv_2 _19256_ (.A(_02271_),
    .Y(_00191_));
 sky130_fd_sc_hd__inv_2 _19257_ (.A(_02271_),
    .Y(_00192_));
 sky130_fd_sc_hd__inv_2 _19258_ (.A(_02271_),
    .Y(_00193_));
 sky130_fd_sc_hd__inv_2 _19259_ (.A(_02271_),
    .Y(_00194_));
 sky130_fd_sc_hd__inv_2 _19260_ (.A(_02271_),
    .Y(_00195_));
 sky130_fd_sc_hd__inv_2 _19261_ (.A(_02271_),
    .Y(_00196_));
 sky130_fd_sc_hd__inv_2 _19262_ (.A(_02271_),
    .Y(_00197_));
 sky130_fd_sc_hd__and3_1 _19263_ (.A(_01513_),
    .B(_01608_),
    .C(_01750_),
    .X(_02272_));
 sky130_fd_sc_hd__and3b_1 _19264_ (.A_N(\wfg_stim_mem_top.wbs_ack_o ),
    .B(_01697_),
    .C(_02272_),
    .X(_02273_));
 sky130_fd_sc_hd__clkbuf_1 _19265_ (.A(_02273_),
    .X(_00851_));
 sky130_fd_sc_hd__inv_2 _19266_ (.A(_02271_),
    .Y(_00198_));
 sky130_fd_sc_hd__inv_2 _19267_ (.A(_02271_),
    .Y(_00199_));
 sky130_fd_sc_hd__inv_2 _19268_ (.A(_02271_),
    .Y(_00200_));
 sky130_fd_sc_hd__buf_4 _19269_ (.A(_02142_),
    .X(_02274_));
 sky130_fd_sc_hd__inv_2 _19270_ (.A(_02274_),
    .Y(_00201_));
 sky130_fd_sc_hd__inv_2 _19271_ (.A(_02274_),
    .Y(_00202_));
 sky130_fd_sc_hd__inv_2 _19272_ (.A(_02274_),
    .Y(_00203_));
 sky130_fd_sc_hd__inv_2 _19273_ (.A(_02274_),
    .Y(_00204_));
 sky130_fd_sc_hd__inv_2 _19274_ (.A(_02274_),
    .Y(_00205_));
 sky130_fd_sc_hd__inv_2 _19275_ (.A(_02274_),
    .Y(_00206_));
 sky130_fd_sc_hd__inv_2 _19276_ (.A(_02274_),
    .Y(_00207_));
 sky130_fd_sc_hd__inv_2 _19277_ (.A(_02274_),
    .Y(_00208_));
 sky130_fd_sc_hd__inv_2 _19278_ (.A(_02274_),
    .Y(_00209_));
 sky130_fd_sc_hd__inv_2 _19279_ (.A(_02274_),
    .Y(_00210_));
 sky130_fd_sc_hd__buf_4 _19280_ (.A(_02142_),
    .X(_02275_));
 sky130_fd_sc_hd__inv_2 _19281_ (.A(_02275_),
    .Y(_00211_));
 sky130_fd_sc_hd__inv_2 _19282_ (.A(_02275_),
    .Y(_00212_));
 sky130_fd_sc_hd__inv_2 _19283_ (.A(_02275_),
    .Y(_00213_));
 sky130_fd_sc_hd__inv_2 _19284_ (.A(_02275_),
    .Y(_00214_));
 sky130_fd_sc_hd__inv_2 _19285_ (.A(_02275_),
    .Y(_00215_));
 sky130_fd_sc_hd__inv_2 _19286_ (.A(_02275_),
    .Y(_00216_));
 sky130_fd_sc_hd__inv_2 _19287_ (.A(_02275_),
    .Y(_00217_));
 sky130_fd_sc_hd__inv_2 _19288_ (.A(_02275_),
    .Y(_00218_));
 sky130_fd_sc_hd__inv_2 _19289_ (.A(_02275_),
    .Y(_00219_));
 sky130_fd_sc_hd__inv_2 _19290_ (.A(_02275_),
    .Y(_00220_));
 sky130_fd_sc_hd__buf_4 _19291_ (.A(_02142_),
    .X(_02276_));
 sky130_fd_sc_hd__inv_2 _19292_ (.A(_02276_),
    .Y(_00221_));
 sky130_fd_sc_hd__inv_2 _19293_ (.A(_02276_),
    .Y(_00222_));
 sky130_fd_sc_hd__inv_2 _19294_ (.A(_02276_),
    .Y(_00223_));
 sky130_fd_sc_hd__inv_2 _19295_ (.A(_02276_),
    .Y(_00224_));
 sky130_fd_sc_hd__inv_2 _19296_ (.A(_02276_),
    .Y(_00225_));
 sky130_fd_sc_hd__inv_2 _19297_ (.A(_02276_),
    .Y(_00226_));
 sky130_fd_sc_hd__inv_2 _19298_ (.A(_02276_),
    .Y(_00227_));
 sky130_fd_sc_hd__inv_2 _19299_ (.A(_02276_),
    .Y(_00228_));
 sky130_fd_sc_hd__inv_2 _19300_ (.A(_02276_),
    .Y(_00229_));
 sky130_fd_sc_hd__inv_2 _19301_ (.A(_02276_),
    .Y(_00230_));
 sky130_fd_sc_hd__buf_6 _19302_ (.A(_02142_),
    .X(_02277_));
 sky130_fd_sc_hd__inv_2 _19303_ (.A(_02277_),
    .Y(_00231_));
 sky130_fd_sc_hd__inv_2 _19304_ (.A(_02277_),
    .Y(_00232_));
 sky130_fd_sc_hd__inv_2 _19305_ (.A(_02277_),
    .Y(_00233_));
 sky130_fd_sc_hd__inv_2 _19306_ (.A(_02277_),
    .Y(_00234_));
 sky130_fd_sc_hd__inv_2 _19307_ (.A(_02277_),
    .Y(_00235_));
 sky130_fd_sc_hd__inv_2 _19308_ (.A(_02277_),
    .Y(_00236_));
 sky130_fd_sc_hd__inv_2 _19309_ (.A(_02277_),
    .Y(_00237_));
 sky130_fd_sc_hd__inv_2 _19310_ (.A(_02277_),
    .Y(_00238_));
 sky130_fd_sc_hd__inv_2 _19311_ (.A(_02277_),
    .Y(_00239_));
 sky130_fd_sc_hd__inv_2 _19312_ (.A(_02277_),
    .Y(_00240_));
 sky130_fd_sc_hd__buf_6 _19313_ (.A(_02142_),
    .X(_02278_));
 sky130_fd_sc_hd__inv_2 _19314_ (.A(_02278_),
    .Y(_00241_));
 sky130_fd_sc_hd__inv_2 _19315_ (.A(_02278_),
    .Y(_00242_));
 sky130_fd_sc_hd__inv_2 _19316_ (.A(_02278_),
    .Y(_00243_));
 sky130_fd_sc_hd__inv_2 _19317_ (.A(_02278_),
    .Y(_00244_));
 sky130_fd_sc_hd__inv_2 _19318_ (.A(_02278_),
    .Y(_00245_));
 sky130_fd_sc_hd__inv_2 _19319_ (.A(_02278_),
    .Y(_00246_));
 sky130_fd_sc_hd__inv_2 _19320_ (.A(_02278_),
    .Y(_00247_));
 sky130_fd_sc_hd__inv_2 _19321_ (.A(_02278_),
    .Y(_00248_));
 sky130_fd_sc_hd__inv_2 _19322_ (.A(_02278_),
    .Y(_00249_));
 sky130_fd_sc_hd__inv_2 _19323_ (.A(_02278_),
    .Y(_00250_));
 sky130_fd_sc_hd__buf_4 _19324_ (.A(_02142_),
    .X(_02279_));
 sky130_fd_sc_hd__inv_2 _19325_ (.A(_02279_),
    .Y(_00251_));
 sky130_fd_sc_hd__inv_2 _19326_ (.A(_02279_),
    .Y(_00252_));
 sky130_fd_sc_hd__inv_2 _19327_ (.A(_02279_),
    .Y(_00253_));
 sky130_fd_sc_hd__inv_2 _19328_ (.A(_02279_),
    .Y(_00254_));
 sky130_fd_sc_hd__inv_2 _19329_ (.A(_02279_),
    .Y(_00255_));
 sky130_fd_sc_hd__inv_2 _19330_ (.A(_02279_),
    .Y(_00256_));
 sky130_fd_sc_hd__inv_2 _19331_ (.A(_02279_),
    .Y(_00257_));
 sky130_fd_sc_hd__inv_2 _19332_ (.A(_02279_),
    .Y(_00258_));
 sky130_fd_sc_hd__inv_2 _19333_ (.A(_02279_),
    .Y(_00259_));
 sky130_fd_sc_hd__inv_2 _19334_ (.A(_02279_),
    .Y(_00260_));
 sky130_fd_sc_hd__buf_6 _19335_ (.A(_02142_),
    .X(_02280_));
 sky130_fd_sc_hd__inv_2 _19336_ (.A(_02280_),
    .Y(_00261_));
 sky130_fd_sc_hd__inv_2 _19337_ (.A(_02280_),
    .Y(_00262_));
 sky130_fd_sc_hd__inv_2 _19338_ (.A(_02280_),
    .Y(_00263_));
 sky130_fd_sc_hd__inv_2 _19339_ (.A(_02280_),
    .Y(_00264_));
 sky130_fd_sc_hd__inv_2 _19340_ (.A(_02280_),
    .Y(_00265_));
 sky130_fd_sc_hd__inv_2 _19341_ (.A(_02280_),
    .Y(_00266_));
 sky130_fd_sc_hd__inv_2 _19342_ (.A(_02280_),
    .Y(_00267_));
 sky130_fd_sc_hd__inv_2 _19343_ (.A(_02280_),
    .Y(_00268_));
 sky130_fd_sc_hd__inv_2 _19344_ (.A(_02280_),
    .Y(_00269_));
 sky130_fd_sc_hd__inv_2 _19345_ (.A(_02280_),
    .Y(_00270_));
 sky130_fd_sc_hd__buf_12 _19346_ (.A(net98),
    .X(_02281_));
 sky130_fd_sc_hd__buf_4 _19347_ (.A(_02281_),
    .X(_02282_));
 sky130_fd_sc_hd__inv_2 _19348_ (.A(_02282_),
    .Y(_00271_));
 sky130_fd_sc_hd__inv_2 _19349_ (.A(_02282_),
    .Y(_00272_));
 sky130_fd_sc_hd__inv_2 _19350_ (.A(_02282_),
    .Y(_00273_));
 sky130_fd_sc_hd__inv_2 _19351_ (.A(_02282_),
    .Y(_00274_));
 sky130_fd_sc_hd__inv_2 _19352_ (.A(_02282_),
    .Y(_00275_));
 sky130_fd_sc_hd__inv_2 _19353_ (.A(_02282_),
    .Y(_00276_));
 sky130_fd_sc_hd__inv_2 _19354_ (.A(_02282_),
    .Y(_00277_));
 sky130_fd_sc_hd__inv_2 _19355_ (.A(_02282_),
    .Y(_00278_));
 sky130_fd_sc_hd__inv_2 _19356_ (.A(_02282_),
    .Y(_00279_));
 sky130_fd_sc_hd__inv_2 _19357_ (.A(_02282_),
    .Y(_00280_));
 sky130_fd_sc_hd__buf_6 _19358_ (.A(_02281_),
    .X(_02283_));
 sky130_fd_sc_hd__inv_2 _19359_ (.A(_02283_),
    .Y(_00281_));
 sky130_fd_sc_hd__inv_2 _19360_ (.A(_02283_),
    .Y(_00282_));
 sky130_fd_sc_hd__inv_2 _19361_ (.A(_02283_),
    .Y(_00283_));
 sky130_fd_sc_hd__inv_2 _19362_ (.A(_02283_),
    .Y(_00284_));
 sky130_fd_sc_hd__inv_2 _19363_ (.A(_02283_),
    .Y(_00285_));
 sky130_fd_sc_hd__inv_2 _19364_ (.A(_02283_),
    .Y(_00286_));
 sky130_fd_sc_hd__inv_2 _19365_ (.A(_02283_),
    .Y(_00287_));
 sky130_fd_sc_hd__inv_2 _19366_ (.A(_02283_),
    .Y(_00288_));
 sky130_fd_sc_hd__inv_2 _19367_ (.A(_02283_),
    .Y(_00289_));
 sky130_fd_sc_hd__inv_2 _19368_ (.A(_02283_),
    .Y(_00290_));
 sky130_fd_sc_hd__buf_4 _19369_ (.A(_02281_),
    .X(_02284_));
 sky130_fd_sc_hd__inv_2 _19370_ (.A(_02284_),
    .Y(_00291_));
 sky130_fd_sc_hd__inv_2 _19371_ (.A(_02284_),
    .Y(_00292_));
 sky130_fd_sc_hd__inv_2 _19372_ (.A(_02284_),
    .Y(_00293_));
 sky130_fd_sc_hd__inv_2 _19373_ (.A(_02284_),
    .Y(_00294_));
 sky130_fd_sc_hd__inv_2 _19374_ (.A(_02284_),
    .Y(_00295_));
 sky130_fd_sc_hd__inv_2 _19375_ (.A(_02284_),
    .Y(_00296_));
 sky130_fd_sc_hd__inv_2 _19376_ (.A(_02284_),
    .Y(_00297_));
 sky130_fd_sc_hd__inv_2 _19377_ (.A(_02284_),
    .Y(_00298_));
 sky130_fd_sc_hd__inv_2 _19378_ (.A(_02284_),
    .Y(_00299_));
 sky130_fd_sc_hd__inv_2 _19379_ (.A(_02284_),
    .Y(_00300_));
 sky130_fd_sc_hd__buf_6 _19380_ (.A(_02281_),
    .X(_02285_));
 sky130_fd_sc_hd__inv_2 _19381_ (.A(_02285_),
    .Y(_00301_));
 sky130_fd_sc_hd__inv_2 _19382_ (.A(_02285_),
    .Y(_00302_));
 sky130_fd_sc_hd__inv_2 _19383_ (.A(_02285_),
    .Y(_00303_));
 sky130_fd_sc_hd__inv_2 _19384_ (.A(_02285_),
    .Y(_00304_));
 sky130_fd_sc_hd__inv_2 _19385_ (.A(_02285_),
    .Y(_00305_));
 sky130_fd_sc_hd__inv_2 _19386_ (.A(_02285_),
    .Y(_00306_));
 sky130_fd_sc_hd__inv_2 _19387_ (.A(_02285_),
    .Y(_00307_));
 sky130_fd_sc_hd__inv_2 _19388_ (.A(_02285_),
    .Y(_00308_));
 sky130_fd_sc_hd__inv_2 _19389_ (.A(_02285_),
    .Y(_00309_));
 sky130_fd_sc_hd__inv_2 _19390_ (.A(_02285_),
    .Y(_00310_));
 sky130_fd_sc_hd__buf_4 _19391_ (.A(_02281_),
    .X(_02286_));
 sky130_fd_sc_hd__inv_2 _19392_ (.A(_02286_),
    .Y(_00311_));
 sky130_fd_sc_hd__inv_2 _19393_ (.A(_02286_),
    .Y(_00312_));
 sky130_fd_sc_hd__inv_2 _19394_ (.A(_02286_),
    .Y(_00313_));
 sky130_fd_sc_hd__inv_2 _19395_ (.A(_02286_),
    .Y(_00314_));
 sky130_fd_sc_hd__inv_2 _19396_ (.A(_02286_),
    .Y(_00315_));
 sky130_fd_sc_hd__inv_2 _19397_ (.A(_02286_),
    .Y(_00316_));
 sky130_fd_sc_hd__inv_2 _19398_ (.A(_02286_),
    .Y(_00317_));
 sky130_fd_sc_hd__inv_2 _19399_ (.A(_02286_),
    .Y(_00318_));
 sky130_fd_sc_hd__inv_2 _19400_ (.A(_02286_),
    .Y(_00319_));
 sky130_fd_sc_hd__inv_2 _19401_ (.A(_02286_),
    .Y(_00320_));
 sky130_fd_sc_hd__buf_6 _19402_ (.A(_02281_),
    .X(_02287_));
 sky130_fd_sc_hd__inv_2 _19403_ (.A(_02287_),
    .Y(_00321_));
 sky130_fd_sc_hd__inv_2 _19404_ (.A(_02287_),
    .Y(_00322_));
 sky130_fd_sc_hd__inv_2 _19405_ (.A(_02287_),
    .Y(_00323_));
 sky130_fd_sc_hd__inv_2 _19406_ (.A(_02287_),
    .Y(_00324_));
 sky130_fd_sc_hd__and3_1 _19407_ (.A(_01429_),
    .B(_01750_),
    .C(_01706_),
    .X(_02288_));
 sky130_fd_sc_hd__clkbuf_4 _19408_ (.A(_02288_),
    .X(_02289_));
 sky130_fd_sc_hd__or2_1 _19409_ (.A(\wfg_stim_mem_top.wbs_dat_o[0] ),
    .B(_02289_),
    .X(_02290_));
 sky130_fd_sc_hd__or2_2 _19410_ (.A(_01424_),
    .B(_01428_),
    .X(_02291_));
 sky130_fd_sc_hd__nor2_4 _19411_ (.A(_02291_),
    .B(_01959_),
    .Y(_02292_));
 sky130_fd_sc_hd__and3_2 _19412_ (.A(_01429_),
    .B(_01959_),
    .C(_01689_),
    .X(_02293_));
 sky130_fd_sc_hd__buf_4 _19413_ (.A(_02293_),
    .X(_02294_));
 sky130_fd_sc_hd__nand2_1 _19414_ (.A(_01429_),
    .B(_01690_),
    .Y(_02295_));
 sky130_fd_sc_hd__nor2_2 _19415_ (.A(_02291_),
    .B(_01763_),
    .Y(_02296_));
 sky130_fd_sc_hd__or3_2 _19416_ (.A(_02291_),
    .B(_01686_),
    .C(_01713_),
    .X(_02297_));
 sky130_fd_sc_hd__a221o_1 _19417_ (.A1(\wfg_stim_mem_top.ctrl_en_q ),
    .A2(_02295_),
    .B1(_02296_),
    .B2(\wfg_stim_mem_top.end_val_q[0] ),
    .C1(_02297_),
    .X(_02298_));
 sky130_fd_sc_hd__a221o_1 _19418_ (.A1(\wfg_stim_mem_top.start_val_q[0] ),
    .A2(_02292_),
    .B1(_02294_),
    .B2(\wfg_stim_mem_top.cfg_inc_q[0] ),
    .C1(_02298_),
    .X(_02299_));
 sky130_fd_sc_hd__and3_1 _19419_ (.A(_01685_),
    .B(_02290_),
    .C(_02299_),
    .X(_02300_));
 sky130_fd_sc_hd__clkbuf_1 _19420_ (.A(_02300_),
    .X(_00978_));
 sky130_fd_sc_hd__buf_2 _19421_ (.A(_02289_),
    .X(_02301_));
 sky130_fd_sc_hd__clkbuf_4 _19422_ (.A(_02292_),
    .X(_02302_));
 sky130_fd_sc_hd__clkbuf_4 _19423_ (.A(_02296_),
    .X(_02303_));
 sky130_fd_sc_hd__buf_4 _19424_ (.A(_02297_),
    .X(_02304_));
 sky130_fd_sc_hd__a221o_1 _19425_ (.A1(\wfg_stim_mem_top.cfg_inc_q[1] ),
    .A2(_02294_),
    .B1(_02303_),
    .B2(\wfg_stim_mem_top.end_val_q[1] ),
    .C1(_02304_),
    .X(_02305_));
 sky130_fd_sc_hd__a21o_1 _19426_ (.A1(\wfg_stim_mem_top.start_val_q[1] ),
    .A2(_02302_),
    .B1(_02305_),
    .X(_02306_));
 sky130_fd_sc_hd__buf_2 _19427_ (.A(_01589_),
    .X(_02307_));
 sky130_fd_sc_hd__o211a_1 _19428_ (.A1(\wfg_stim_mem_top.wbs_dat_o[1] ),
    .A2(_02301_),
    .B1(_02306_),
    .C1(_02307_),
    .X(_00979_));
 sky130_fd_sc_hd__a221o_1 _19429_ (.A1(\wfg_stim_mem_top.cfg_inc_q[2] ),
    .A2(_02294_),
    .B1(_02303_),
    .B2(\wfg_stim_mem_top.end_val_q[2] ),
    .C1(_02304_),
    .X(_02308_));
 sky130_fd_sc_hd__a21o_1 _19430_ (.A1(\wfg_stim_mem_top.start_val_q[2] ),
    .A2(_02302_),
    .B1(_02308_),
    .X(_02309_));
 sky130_fd_sc_hd__o211a_1 _19431_ (.A1(\wfg_stim_mem_top.wbs_dat_o[2] ),
    .A2(_02301_),
    .B1(_02309_),
    .C1(_02307_),
    .X(_00980_));
 sky130_fd_sc_hd__clkbuf_4 _19432_ (.A(_02293_),
    .X(_02310_));
 sky130_fd_sc_hd__clkbuf_4 _19433_ (.A(_02297_),
    .X(_02311_));
 sky130_fd_sc_hd__a221o_1 _19434_ (.A1(\wfg_stim_mem_top.start_val_q[3] ),
    .A2(_02292_),
    .B1(_02303_),
    .B2(\wfg_stim_mem_top.end_val_q[3] ),
    .C1(_02311_),
    .X(_02312_));
 sky130_fd_sc_hd__a21o_1 _19435_ (.A1(\wfg_stim_mem_top.cfg_inc_q[3] ),
    .A2(_02310_),
    .B1(_02312_),
    .X(_02313_));
 sky130_fd_sc_hd__o211a_1 _19436_ (.A1(\wfg_stim_mem_top.wbs_dat_o[3] ),
    .A2(_02301_),
    .B1(_02313_),
    .C1(_02307_),
    .X(_00981_));
 sky130_fd_sc_hd__a221o_1 _19437_ (.A1(\wfg_stim_mem_top.cfg_inc_q[4] ),
    .A2(_02294_),
    .B1(_02303_),
    .B2(\wfg_stim_mem_top.end_val_q[4] ),
    .C1(_02311_),
    .X(_02314_));
 sky130_fd_sc_hd__a21o_1 _19438_ (.A1(\wfg_stim_mem_top.start_val_q[4] ),
    .A2(_02302_),
    .B1(_02314_),
    .X(_02315_));
 sky130_fd_sc_hd__o211a_1 _19439_ (.A1(\wfg_stim_mem_top.wbs_dat_o[4] ),
    .A2(_02301_),
    .B1(_02315_),
    .C1(_02307_),
    .X(_00982_));
 sky130_fd_sc_hd__a221o_1 _19440_ (.A1(\wfg_stim_mem_top.cfg_inc_q[5] ),
    .A2(_02294_),
    .B1(_02303_),
    .B2(\wfg_stim_mem_top.end_val_q[5] ),
    .C1(_02311_),
    .X(_02316_));
 sky130_fd_sc_hd__a21o_1 _19441_ (.A1(\wfg_stim_mem_top.start_val_q[5] ),
    .A2(_02302_),
    .B1(_02316_),
    .X(_02317_));
 sky130_fd_sc_hd__o211a_1 _19442_ (.A1(\wfg_stim_mem_top.wbs_dat_o[5] ),
    .A2(_02301_),
    .B1(_02317_),
    .C1(_02307_),
    .X(_00983_));
 sky130_fd_sc_hd__a221o_1 _19443_ (.A1(\wfg_stim_mem_top.cfg_inc_q[6] ),
    .A2(_02294_),
    .B1(_02303_),
    .B2(\wfg_stim_mem_top.end_val_q[6] ),
    .C1(_02311_),
    .X(_02318_));
 sky130_fd_sc_hd__a21o_1 _19444_ (.A1(\wfg_stim_mem_top.start_val_q[6] ),
    .A2(_02302_),
    .B1(_02318_),
    .X(_02319_));
 sky130_fd_sc_hd__o211a_1 _19445_ (.A1(\wfg_stim_mem_top.wbs_dat_o[6] ),
    .A2(_02301_),
    .B1(_02319_),
    .C1(_02307_),
    .X(_00984_));
 sky130_fd_sc_hd__a221o_1 _19446_ (.A1(\wfg_stim_mem_top.cfg_inc_q[7] ),
    .A2(_02294_),
    .B1(_02303_),
    .B2(\wfg_stim_mem_top.end_val_q[7] ),
    .C1(_02311_),
    .X(_02320_));
 sky130_fd_sc_hd__a21o_1 _19447_ (.A1(\wfg_stim_mem_top.start_val_q[7] ),
    .A2(_02302_),
    .B1(_02320_),
    .X(_02321_));
 sky130_fd_sc_hd__o211a_1 _19448_ (.A1(\wfg_stim_mem_top.wbs_dat_o[7] ),
    .A2(_02301_),
    .B1(_02321_),
    .C1(_02307_),
    .X(_00985_));
 sky130_fd_sc_hd__a221o_1 _19449_ (.A1(\wfg_stim_mem_top.start_val_q[8] ),
    .A2(_02292_),
    .B1(_02303_),
    .B2(\wfg_stim_mem_top.end_val_q[8] ),
    .C1(_02311_),
    .X(_02322_));
 sky130_fd_sc_hd__a21o_1 _19450_ (.A1(_04081_),
    .A2(_02310_),
    .B1(_02322_),
    .X(_02323_));
 sky130_fd_sc_hd__o211a_1 _19451_ (.A1(\wfg_stim_mem_top.wbs_dat_o[8] ),
    .A2(_02301_),
    .B1(_02323_),
    .C1(_02307_),
    .X(_00986_));
 sky130_fd_sc_hd__a221o_1 _19452_ (.A1(_03492_),
    .A2(_02293_),
    .B1(_02303_),
    .B2(\wfg_stim_mem_top.end_val_q[9] ),
    .C1(_02311_),
    .X(_02324_));
 sky130_fd_sc_hd__a21o_1 _19453_ (.A1(\wfg_stim_mem_top.start_val_q[9] ),
    .A2(_02302_),
    .B1(_02324_),
    .X(_02325_));
 sky130_fd_sc_hd__o211a_1 _19454_ (.A1(\wfg_stim_mem_top.wbs_dat_o[9] ),
    .A2(_02301_),
    .B1(_02325_),
    .C1(_02307_),
    .X(_00987_));
 sky130_fd_sc_hd__a221o_1 _19455_ (.A1(_03435_),
    .A2(_02293_),
    .B1(_02303_),
    .B2(\wfg_stim_mem_top.end_val_q[10] ),
    .C1(_02311_),
    .X(_02326_));
 sky130_fd_sc_hd__a21o_1 _19456_ (.A1(\wfg_stim_mem_top.start_val_q[10] ),
    .A2(_02302_),
    .B1(_02326_),
    .X(_02327_));
 sky130_fd_sc_hd__o211a_1 _19457_ (.A1(\wfg_stim_mem_top.wbs_dat_o[10] ),
    .A2(_02301_),
    .B1(_02327_),
    .C1(_02307_),
    .X(_00988_));
 sky130_fd_sc_hd__a221o_1 _19458_ (.A1(_02909_),
    .A2(_02293_),
    .B1(_02296_),
    .B2(\wfg_stim_mem_top.end_val_q[11] ),
    .C1(_02311_),
    .X(_02328_));
 sky130_fd_sc_hd__a21o_1 _19459_ (.A1(\wfg_stim_mem_top.start_val_q[11] ),
    .A2(_02302_),
    .B1(_02328_),
    .X(_02329_));
 sky130_fd_sc_hd__clkbuf_4 _19460_ (.A(_01589_),
    .X(_02330_));
 sky130_fd_sc_hd__o211a_1 _19461_ (.A1(\wfg_stim_mem_top.wbs_dat_o[11] ),
    .A2(_02289_),
    .B1(_02329_),
    .C1(_02330_),
    .X(_00989_));
 sky130_fd_sc_hd__a221o_1 _19462_ (.A1(\wfg_stim_mem_top.start_val_q[12] ),
    .A2(_02292_),
    .B1(_02296_),
    .B2(\wfg_stim_mem_top.end_val_q[12] ),
    .C1(_02311_),
    .X(_02331_));
 sky130_fd_sc_hd__a21o_1 _19463_ (.A1(_02897_),
    .A2(_02310_),
    .B1(_02331_),
    .X(_02332_));
 sky130_fd_sc_hd__o211a_1 _19464_ (.A1(\wfg_stim_mem_top.wbs_dat_o[12] ),
    .A2(_02289_),
    .B1(_02332_),
    .C1(_02330_),
    .X(_00990_));
 sky130_fd_sc_hd__a221o_1 _19465_ (.A1(_02895_),
    .A2(_02293_),
    .B1(_02296_),
    .B2(\wfg_stim_mem_top.end_val_q[13] ),
    .C1(_02297_),
    .X(_02333_));
 sky130_fd_sc_hd__a21o_1 _19466_ (.A1(\wfg_stim_mem_top.start_val_q[13] ),
    .A2(_02302_),
    .B1(_02333_),
    .X(_02334_));
 sky130_fd_sc_hd__o211a_1 _19467_ (.A1(\wfg_stim_mem_top.wbs_dat_o[13] ),
    .A2(_02289_),
    .B1(_02334_),
    .C1(_02330_),
    .X(_00991_));
 sky130_fd_sc_hd__a221o_1 _19468_ (.A1(\wfg_stim_mem_top.start_val_q[14] ),
    .A2(_02292_),
    .B1(_02296_),
    .B2(\wfg_stim_mem_top.end_val_q[14] ),
    .C1(_02297_),
    .X(_02335_));
 sky130_fd_sc_hd__a21o_1 _19469_ (.A1(_02918_),
    .A2(_02310_),
    .B1(_02335_),
    .X(_02336_));
 sky130_fd_sc_hd__o211a_1 _19470_ (.A1(\wfg_stim_mem_top.wbs_dat_o[14] ),
    .A2(_02289_),
    .B1(_02336_),
    .C1(_02330_),
    .X(_00992_));
 sky130_fd_sc_hd__a221o_1 _19471_ (.A1(\wfg_stim_mem_top.start_val_q[15] ),
    .A2(_02292_),
    .B1(_02296_),
    .B2(\wfg_stim_mem_top.end_val_q[15] ),
    .C1(_02297_),
    .X(_02337_));
 sky130_fd_sc_hd__a21o_1 _19472_ (.A1(_02923_),
    .A2(_02310_),
    .B1(_02337_),
    .X(_02338_));
 sky130_fd_sc_hd__o211a_1 _19473_ (.A1(\wfg_stim_mem_top.wbs_dat_o[15] ),
    .A2(_02289_),
    .B1(_02338_),
    .C1(_02330_),
    .X(_00993_));
 sky130_fd_sc_hd__or2_1 _19474_ (.A(\wfg_stim_mem_top.wbs_dat_o[16] ),
    .B(_02289_),
    .X(_02339_));
 sky130_fd_sc_hd__a21o_1 _19475_ (.A1(_02921_),
    .A2(_02310_),
    .B1(_02304_),
    .X(_02340_));
 sky130_fd_sc_hd__and3_1 _19476_ (.A(_01685_),
    .B(_02339_),
    .C(_02340_),
    .X(_02341_));
 sky130_fd_sc_hd__clkbuf_1 _19477_ (.A(_02341_),
    .X(_00994_));
 sky130_fd_sc_hd__or2_1 _19478_ (.A(\wfg_stim_mem_top.wbs_dat_o[17] ),
    .B(_02289_),
    .X(_02342_));
 sky130_fd_sc_hd__a21o_1 _19479_ (.A1(_03142_),
    .A2(_02310_),
    .B1(_02304_),
    .X(_02343_));
 sky130_fd_sc_hd__and3_1 _19480_ (.A(_01685_),
    .B(_02342_),
    .C(_02343_),
    .X(_02344_));
 sky130_fd_sc_hd__clkbuf_1 _19481_ (.A(_02344_),
    .X(_00995_));
 sky130_fd_sc_hd__or2_1 _19482_ (.A(\wfg_stim_mem_top.wbs_dat_o[18] ),
    .B(_02289_),
    .X(_02345_));
 sky130_fd_sc_hd__a21o_1 _19483_ (.A1(_03302_),
    .A2(_02310_),
    .B1(_02304_),
    .X(_02346_));
 sky130_fd_sc_hd__and3_1 _19484_ (.A(_01685_),
    .B(_02345_),
    .C(_02346_),
    .X(_02347_));
 sky130_fd_sc_hd__clkbuf_1 _19485_ (.A(_02347_),
    .X(_00996_));
 sky130_fd_sc_hd__or2_1 _19486_ (.A(\wfg_stim_mem_top.wbs_dat_o[19] ),
    .B(_02288_),
    .X(_02348_));
 sky130_fd_sc_hd__a21o_1 _19487_ (.A1(_02969_),
    .A2(_02310_),
    .B1(_02304_),
    .X(_02349_));
 sky130_fd_sc_hd__and3_1 _19488_ (.A(_01685_),
    .B(_02348_),
    .C(_02349_),
    .X(_02350_));
 sky130_fd_sc_hd__clkbuf_1 _19489_ (.A(_02350_),
    .X(_00997_));
 sky130_fd_sc_hd__or2_1 _19490_ (.A(\wfg_stim_mem_top.wbs_dat_o[20] ),
    .B(_02288_),
    .X(_02351_));
 sky130_fd_sc_hd__a21o_1 _19491_ (.A1(_02950_),
    .A2(_02310_),
    .B1(_02304_),
    .X(_02352_));
 sky130_fd_sc_hd__and3_1 _19492_ (.A(_01730_),
    .B(_02351_),
    .C(_02352_),
    .X(_02353_));
 sky130_fd_sc_hd__clkbuf_1 _19493_ (.A(_02353_),
    .X(_00998_));
 sky130_fd_sc_hd__or2_1 _19494_ (.A(\wfg_stim_mem_top.wbs_dat_o[21] ),
    .B(_02288_),
    .X(_02354_));
 sky130_fd_sc_hd__a21o_1 _19495_ (.A1(_02986_),
    .A2(_02294_),
    .B1(_02304_),
    .X(_02355_));
 sky130_fd_sc_hd__and3_1 _19496_ (.A(_01730_),
    .B(_02354_),
    .C(_02355_),
    .X(_02356_));
 sky130_fd_sc_hd__clkbuf_1 _19497_ (.A(_02356_),
    .X(_00999_));
 sky130_fd_sc_hd__or2_1 _19498_ (.A(\wfg_stim_mem_top.wbs_dat_o[22] ),
    .B(_02288_),
    .X(_02357_));
 sky130_fd_sc_hd__a21o_1 _19499_ (.A1(_02988_),
    .A2(_02294_),
    .B1(_02304_),
    .X(_02358_));
 sky130_fd_sc_hd__and3_1 _19500_ (.A(_01730_),
    .B(_02357_),
    .C(_02358_),
    .X(_02359_));
 sky130_fd_sc_hd__clkbuf_1 _19501_ (.A(_02359_),
    .X(_01000_));
 sky130_fd_sc_hd__or2_1 _19502_ (.A(\wfg_stim_mem_top.wbs_dat_o[23] ),
    .B(_02288_),
    .X(_02360_));
 sky130_fd_sc_hd__a21o_1 _19503_ (.A1(_03016_),
    .A2(_02294_),
    .B1(_02304_),
    .X(_02361_));
 sky130_fd_sc_hd__and3_1 _19504_ (.A(_01730_),
    .B(_02360_),
    .C(_02361_),
    .X(_02362_));
 sky130_fd_sc_hd__clkbuf_1 _19505_ (.A(_02362_),
    .X(_01001_));
 sky130_fd_sc_hd__or3_2 _19506_ (.A(_02147_),
    .B(_01605_),
    .C(_01607_),
    .X(_02363_));
 sky130_fd_sc_hd__o21ai_1 _19507_ (.A1(_01691_),
    .A2(_02363_),
    .B1(_09610_),
    .Y(_02364_));
 sky130_fd_sc_hd__or3_1 _19508_ (.A(_01884_),
    .B(_01691_),
    .C(_02363_),
    .X(_02365_));
 sky130_fd_sc_hd__and3_1 _19509_ (.A(_01730_),
    .B(_02364_),
    .C(_02365_),
    .X(_02366_));
 sky130_fd_sc_hd__clkbuf_1 _19510_ (.A(_02366_),
    .X(_01002_));
 sky130_fd_sc_hd__or3_1 _19511_ (.A(_02147_),
    .B(_01762_),
    .C(_02363_),
    .X(_02367_));
 sky130_fd_sc_hd__buf_2 _19512_ (.A(_02367_),
    .X(_02368_));
 sky130_fd_sc_hd__clkbuf_4 _19513_ (.A(_02368_),
    .X(_02369_));
 sky130_fd_sc_hd__mux2_1 _19514_ (.A0(_01884_),
    .A1(_07043_),
    .S(_02369_),
    .X(_02370_));
 sky130_fd_sc_hd__and2_1 _19515_ (.A(_02116_),
    .B(_02370_),
    .X(_02371_));
 sky130_fd_sc_hd__clkbuf_1 _19516_ (.A(_02371_),
    .X(_01003_));
 sky130_fd_sc_hd__clkbuf_2 _19517_ (.A(_02048_),
    .X(_02372_));
 sky130_fd_sc_hd__mux2_1 _19518_ (.A0(net77),
    .A1(_07044_),
    .S(_02369_),
    .X(_02373_));
 sky130_fd_sc_hd__and2_1 _19519_ (.A(_02372_),
    .B(_02373_),
    .X(_02374_));
 sky130_fd_sc_hd__clkbuf_1 _19520_ (.A(_02374_),
    .X(_01004_));
 sky130_fd_sc_hd__mux2_1 _19521_ (.A0(_01666_),
    .A1(_06605_),
    .S(_02369_),
    .X(_02375_));
 sky130_fd_sc_hd__and2_1 _19522_ (.A(_02372_),
    .B(_02375_),
    .X(_02376_));
 sky130_fd_sc_hd__clkbuf_1 _19523_ (.A(_02376_),
    .X(_01005_));
 sky130_fd_sc_hd__mux2_1 _19524_ (.A0(_01669_),
    .A1(_07206_),
    .S(_02369_),
    .X(_02377_));
 sky130_fd_sc_hd__and2_1 _19525_ (.A(_02372_),
    .B(_02377_),
    .X(_02378_));
 sky130_fd_sc_hd__clkbuf_1 _19526_ (.A(_02378_),
    .X(_01006_));
 sky130_fd_sc_hd__mux2_1 _19527_ (.A0(_01672_),
    .A1(_06551_),
    .S(_02369_),
    .X(_02379_));
 sky130_fd_sc_hd__and2_1 _19528_ (.A(_02372_),
    .B(_02379_),
    .X(_02380_));
 sky130_fd_sc_hd__clkbuf_1 _19529_ (.A(_02380_),
    .X(_01007_));
 sky130_fd_sc_hd__mux2_1 _19530_ (.A0(_01675_),
    .A1(_06549_),
    .S(_02369_),
    .X(_02381_));
 sky130_fd_sc_hd__and2_1 _19531_ (.A(_02372_),
    .B(_02381_),
    .X(_02382_));
 sky130_fd_sc_hd__clkbuf_1 _19532_ (.A(_02382_),
    .X(_01008_));
 sky130_fd_sc_hd__mux2_1 _19533_ (.A0(_01679_),
    .A1(_06547_),
    .S(_02369_),
    .X(_02383_));
 sky130_fd_sc_hd__and2_1 _19534_ (.A(_02372_),
    .B(_02383_),
    .X(_02384_));
 sky130_fd_sc_hd__clkbuf_1 _19535_ (.A(_02384_),
    .X(_01009_));
 sky130_fd_sc_hd__mux2_1 _19536_ (.A0(_01682_),
    .A1(_06486_),
    .S(_02369_),
    .X(_02385_));
 sky130_fd_sc_hd__and2_1 _19537_ (.A(_02372_),
    .B(_02385_),
    .X(_02386_));
 sky130_fd_sc_hd__clkbuf_1 _19538_ (.A(_02386_),
    .X(_01010_));
 sky130_fd_sc_hd__mux2_1 _19539_ (.A0(_01601_),
    .A1(_06725_),
    .S(_02369_),
    .X(_02387_));
 sky130_fd_sc_hd__and2_1 _19540_ (.A(_02372_),
    .B(_02387_),
    .X(_02388_));
 sky130_fd_sc_hd__clkbuf_1 _19541_ (.A(_02388_),
    .X(_01011_));
 sky130_fd_sc_hd__mux2_1 _19542_ (.A0(_01620_),
    .A1(_06714_),
    .S(_02369_),
    .X(_02389_));
 sky130_fd_sc_hd__and2_1 _19543_ (.A(_02372_),
    .B(_02389_),
    .X(_02390_));
 sky130_fd_sc_hd__clkbuf_1 _19544_ (.A(_02390_),
    .X(_01012_));
 sky130_fd_sc_hd__mux2_1 _19545_ (.A0(_01624_),
    .A1(_06451_),
    .S(_02368_),
    .X(_02391_));
 sky130_fd_sc_hd__and2_1 _19546_ (.A(_02372_),
    .B(_02391_),
    .X(_02392_));
 sky130_fd_sc_hd__clkbuf_1 _19547_ (.A(_02392_),
    .X(_01013_));
 sky130_fd_sc_hd__buf_2 _19548_ (.A(_02048_),
    .X(_02393_));
 sky130_fd_sc_hd__mux2_1 _19549_ (.A0(_01627_),
    .A1(_06471_),
    .S(_02368_),
    .X(_02394_));
 sky130_fd_sc_hd__and2_1 _19550_ (.A(_02393_),
    .B(_02394_),
    .X(_02395_));
 sky130_fd_sc_hd__clkbuf_1 _19551_ (.A(_02395_),
    .X(_01014_));
 sky130_fd_sc_hd__mux2_1 _19552_ (.A0(_01630_),
    .A1(_06474_),
    .S(_02368_),
    .X(_02396_));
 sky130_fd_sc_hd__and2_1 _19553_ (.A(_02393_),
    .B(_02396_),
    .X(_02397_));
 sky130_fd_sc_hd__clkbuf_1 _19554_ (.A(_02397_),
    .X(_01015_));
 sky130_fd_sc_hd__mux2_1 _19555_ (.A0(_01633_),
    .A1(_06509_),
    .S(_02368_),
    .X(_02398_));
 sky130_fd_sc_hd__and2_1 _19556_ (.A(_02393_),
    .B(_02398_),
    .X(_02399_));
 sky130_fd_sc_hd__clkbuf_1 _19557_ (.A(_02399_),
    .X(_01016_));
 sky130_fd_sc_hd__mux2_1 _19558_ (.A0(net71),
    .A1(_06505_),
    .S(_02368_),
    .X(_02400_));
 sky130_fd_sc_hd__or2_1 _19559_ (.A(_01837_),
    .B(_02400_),
    .X(_02401_));
 sky130_fd_sc_hd__clkbuf_1 _19560_ (.A(_02401_),
    .X(_01017_));
 sky130_fd_sc_hd__mux2_1 _19561_ (.A0(_01639_),
    .A1(_08082_),
    .S(_02368_),
    .X(_02402_));
 sky130_fd_sc_hd__and2_1 _19562_ (.A(_02393_),
    .B(_02402_),
    .X(_02403_));
 sky130_fd_sc_hd__clkbuf_1 _19563_ (.A(_02403_),
    .X(_01018_));
 sky130_fd_sc_hd__or2_1 _19564_ (.A(_01604_),
    .B(_02363_),
    .X(_02404_));
 sky130_fd_sc_hd__clkbuf_4 _19565_ (.A(_02404_),
    .X(_02405_));
 sky130_fd_sc_hd__buf_4 _19566_ (.A(_02405_),
    .X(_02406_));
 sky130_fd_sc_hd__mux2_1 _19567_ (.A0(_01884_),
    .A1(\wfg_stim_sine_top.inc_val_q[0] ),
    .S(_02406_),
    .X(_02407_));
 sky130_fd_sc_hd__and2_1 _19568_ (.A(_02393_),
    .B(_02407_),
    .X(_02408_));
 sky130_fd_sc_hd__clkbuf_1 _19569_ (.A(_02408_),
    .X(_01019_));
 sky130_fd_sc_hd__mux2_1 _19570_ (.A0(net77),
    .A1(\wfg_stim_sine_top.inc_val_q[1] ),
    .S(_02406_),
    .X(_02409_));
 sky130_fd_sc_hd__and2_1 _19571_ (.A(_02393_),
    .B(_02409_),
    .X(_02410_));
 sky130_fd_sc_hd__clkbuf_1 _19572_ (.A(_02410_),
    .X(_01020_));
 sky130_fd_sc_hd__mux2_1 _19573_ (.A0(_01666_),
    .A1(\wfg_stim_sine_top.inc_val_q[2] ),
    .S(_02406_),
    .X(_02411_));
 sky130_fd_sc_hd__and2_1 _19574_ (.A(_02393_),
    .B(_02411_),
    .X(_02412_));
 sky130_fd_sc_hd__clkbuf_1 _19575_ (.A(_02412_),
    .X(_01021_));
 sky130_fd_sc_hd__mux2_1 _19576_ (.A0(_01669_),
    .A1(\wfg_stim_sine_top.inc_val_q[3] ),
    .S(_02406_),
    .X(_02413_));
 sky130_fd_sc_hd__and2_1 _19577_ (.A(_02393_),
    .B(_02413_),
    .X(_02414_));
 sky130_fd_sc_hd__clkbuf_1 _19578_ (.A(_02414_),
    .X(_01022_));
 sky130_fd_sc_hd__mux2_1 _19579_ (.A0(_01672_),
    .A1(\wfg_stim_sine_top.inc_val_q[4] ),
    .S(_02406_),
    .X(_02415_));
 sky130_fd_sc_hd__and2_1 _19580_ (.A(_02393_),
    .B(_02415_),
    .X(_02416_));
 sky130_fd_sc_hd__clkbuf_1 _19581_ (.A(_02416_),
    .X(_01023_));
 sky130_fd_sc_hd__mux2_1 _19582_ (.A0(_01675_),
    .A1(\wfg_stim_sine_top.inc_val_q[5] ),
    .S(_02406_),
    .X(_02417_));
 sky130_fd_sc_hd__and2_1 _19583_ (.A(_02393_),
    .B(_02417_),
    .X(_02418_));
 sky130_fd_sc_hd__clkbuf_1 _19584_ (.A(_02418_),
    .X(_01024_));
 sky130_fd_sc_hd__buf_2 _19585_ (.A(_02048_),
    .X(_02419_));
 sky130_fd_sc_hd__mux2_1 _19586_ (.A0(_01679_),
    .A1(\wfg_stim_sine_top.inc_val_q[6] ),
    .S(_02406_),
    .X(_02420_));
 sky130_fd_sc_hd__and2_1 _19587_ (.A(_02419_),
    .B(_02420_),
    .X(_02421_));
 sky130_fd_sc_hd__clkbuf_1 _19588_ (.A(_02421_),
    .X(_01025_));
 sky130_fd_sc_hd__mux2_1 _19589_ (.A0(_01682_),
    .A1(\wfg_stim_sine_top.inc_val_q[7] ),
    .S(_02406_),
    .X(_02422_));
 sky130_fd_sc_hd__and2_1 _19590_ (.A(_02419_),
    .B(_02422_),
    .X(_02423_));
 sky130_fd_sc_hd__clkbuf_1 _19591_ (.A(_02423_),
    .X(_01026_));
 sky130_fd_sc_hd__mux2_1 _19592_ (.A0(_01601_),
    .A1(\wfg_stim_sine_top.inc_val_q[8] ),
    .S(_02406_),
    .X(_02424_));
 sky130_fd_sc_hd__and2_1 _19593_ (.A(_02419_),
    .B(_02424_),
    .X(_02425_));
 sky130_fd_sc_hd__clkbuf_1 _19594_ (.A(_02425_),
    .X(_01027_));
 sky130_fd_sc_hd__mux2_1 _19595_ (.A0(_01620_),
    .A1(\wfg_stim_sine_top.inc_val_q[9] ),
    .S(_02406_),
    .X(_02426_));
 sky130_fd_sc_hd__and2_1 _19596_ (.A(_02419_),
    .B(_02426_),
    .X(_02427_));
 sky130_fd_sc_hd__clkbuf_1 _19597_ (.A(_02427_),
    .X(_01028_));
 sky130_fd_sc_hd__mux2_1 _19598_ (.A0(_01624_),
    .A1(\wfg_stim_sine_top.inc_val_q[10] ),
    .S(_02405_),
    .X(_02428_));
 sky130_fd_sc_hd__and2_1 _19599_ (.A(_02419_),
    .B(_02428_),
    .X(_02429_));
 sky130_fd_sc_hd__clkbuf_1 _19600_ (.A(_02429_),
    .X(_01029_));
 sky130_fd_sc_hd__mux2_1 _19601_ (.A0(_01627_),
    .A1(\wfg_stim_sine_top.inc_val_q[11] ),
    .S(_02405_),
    .X(_02430_));
 sky130_fd_sc_hd__and2_1 _19602_ (.A(_02419_),
    .B(_02430_),
    .X(_02431_));
 sky130_fd_sc_hd__clkbuf_1 _19603_ (.A(_02431_),
    .X(_01030_));
 sky130_fd_sc_hd__mux2_1 _19604_ (.A0(net69),
    .A1(\wfg_stim_sine_top.inc_val_q[12] ),
    .S(_02405_),
    .X(_02432_));
 sky130_fd_sc_hd__or2_1 _19605_ (.A(_01837_),
    .B(_02432_),
    .X(_02433_));
 sky130_fd_sc_hd__clkbuf_1 _19606_ (.A(_02433_),
    .X(_01031_));
 sky130_fd_sc_hd__mux2_1 _19607_ (.A0(_01633_),
    .A1(\wfg_stim_sine_top.inc_val_q[13] ),
    .S(_02405_),
    .X(_02434_));
 sky130_fd_sc_hd__and2_1 _19608_ (.A(_02419_),
    .B(_02434_),
    .X(_02435_));
 sky130_fd_sc_hd__clkbuf_1 _19609_ (.A(_02435_),
    .X(_01032_));
 sky130_fd_sc_hd__mux2_1 _19610_ (.A0(_01636_),
    .A1(\wfg_stim_sine_top.inc_val_q[14] ),
    .S(_02405_),
    .X(_02436_));
 sky130_fd_sc_hd__and2_1 _19611_ (.A(_02419_),
    .B(_02436_),
    .X(_02437_));
 sky130_fd_sc_hd__clkbuf_1 _19612_ (.A(_02437_),
    .X(_01033_));
 sky130_fd_sc_hd__mux2_1 _19613_ (.A0(_01639_),
    .A1(\wfg_stim_sine_top.inc_val_q[15] ),
    .S(_02405_),
    .X(_02438_));
 sky130_fd_sc_hd__and2_1 _19614_ (.A(_02419_),
    .B(_02438_),
    .X(_02439_));
 sky130_fd_sc_hd__clkbuf_1 _19615_ (.A(_02439_),
    .X(_01034_));
 sky130_fd_sc_hd__or3_1 _19616_ (.A(_02147_),
    .B(_01756_),
    .C(_02363_),
    .X(_02440_));
 sky130_fd_sc_hd__clkbuf_4 _19617_ (.A(_02440_),
    .X(_02441_));
 sky130_fd_sc_hd__buf_4 _19618_ (.A(_02441_),
    .X(_02442_));
 sky130_fd_sc_hd__mux2_1 _19619_ (.A0(_01884_),
    .A1(\wfg_stim_sine_top.offset_val_q[0] ),
    .S(_02442_),
    .X(_02443_));
 sky130_fd_sc_hd__and2_1 _19620_ (.A(_02419_),
    .B(_02443_),
    .X(_02444_));
 sky130_fd_sc_hd__clkbuf_1 _19621_ (.A(_02444_),
    .X(_01035_));
 sky130_fd_sc_hd__buf_2 _19622_ (.A(_02048_),
    .X(_02445_));
 sky130_fd_sc_hd__mux2_1 _19623_ (.A0(net77),
    .A1(\wfg_stim_sine_top.offset_val_q[1] ),
    .S(_02442_),
    .X(_02446_));
 sky130_fd_sc_hd__and2_1 _19624_ (.A(_02445_),
    .B(_02446_),
    .X(_02447_));
 sky130_fd_sc_hd__clkbuf_1 _19625_ (.A(_02447_),
    .X(_01036_));
 sky130_fd_sc_hd__mux2_1 _19626_ (.A0(net88),
    .A1(\wfg_stim_sine_top.offset_val_q[2] ),
    .S(_02442_),
    .X(_02448_));
 sky130_fd_sc_hd__and2_1 _19627_ (.A(_02445_),
    .B(_02448_),
    .X(_02449_));
 sky130_fd_sc_hd__clkbuf_1 _19628_ (.A(_02449_),
    .X(_01037_));
 sky130_fd_sc_hd__mux2_1 _19629_ (.A0(net91),
    .A1(\wfg_stim_sine_top.offset_val_q[3] ),
    .S(_02442_),
    .X(_02450_));
 sky130_fd_sc_hd__and2_1 _19630_ (.A(_02445_),
    .B(_02450_),
    .X(_02451_));
 sky130_fd_sc_hd__clkbuf_1 _19631_ (.A(_02451_),
    .X(_01038_));
 sky130_fd_sc_hd__mux2_1 _19632_ (.A0(net92),
    .A1(\wfg_stim_sine_top.offset_val_q[4] ),
    .S(_02442_),
    .X(_02452_));
 sky130_fd_sc_hd__and2_1 _19633_ (.A(_02445_),
    .B(_02452_),
    .X(_02453_));
 sky130_fd_sc_hd__clkbuf_1 _19634_ (.A(_02453_),
    .X(_01039_));
 sky130_fd_sc_hd__mux2_1 _19635_ (.A0(net93),
    .A1(\wfg_stim_sine_top.offset_val_q[5] ),
    .S(_02442_),
    .X(_02454_));
 sky130_fd_sc_hd__and2_1 _19636_ (.A(_02445_),
    .B(_02454_),
    .X(_02455_));
 sky130_fd_sc_hd__clkbuf_1 _19637_ (.A(_02455_),
    .X(_01040_));
 sky130_fd_sc_hd__mux2_1 _19638_ (.A0(_01679_),
    .A1(\wfg_stim_sine_top.offset_val_q[6] ),
    .S(_02442_),
    .X(_02456_));
 sky130_fd_sc_hd__and2_1 _19639_ (.A(_02445_),
    .B(_02456_),
    .X(_02457_));
 sky130_fd_sc_hd__clkbuf_1 _19640_ (.A(_02457_),
    .X(_01041_));
 sky130_fd_sc_hd__mux2_1 _19641_ (.A0(_01682_),
    .A1(\wfg_stim_sine_top.offset_val_q[7] ),
    .S(_02442_),
    .X(_02458_));
 sky130_fd_sc_hd__and2_1 _19642_ (.A(_02445_),
    .B(_02458_),
    .X(_02459_));
 sky130_fd_sc_hd__clkbuf_1 _19643_ (.A(_02459_),
    .X(_01042_));
 sky130_fd_sc_hd__mux2_1 _19644_ (.A0(_01601_),
    .A1(\wfg_stim_sine_top.offset_val_q[8] ),
    .S(_02442_),
    .X(_02460_));
 sky130_fd_sc_hd__and2_1 _19645_ (.A(_02445_),
    .B(_02460_),
    .X(_02461_));
 sky130_fd_sc_hd__clkbuf_1 _19646_ (.A(_02461_),
    .X(_01043_));
 sky130_fd_sc_hd__mux2_1 _19647_ (.A0(_01620_),
    .A1(\wfg_stim_sine_top.offset_val_q[9] ),
    .S(_02442_),
    .X(_02462_));
 sky130_fd_sc_hd__and2_1 _19648_ (.A(_02445_),
    .B(_02462_),
    .X(_02463_));
 sky130_fd_sc_hd__clkbuf_1 _19649_ (.A(_02463_),
    .X(_01044_));
 sky130_fd_sc_hd__mux2_1 _19650_ (.A0(_01624_),
    .A1(\wfg_stim_sine_top.offset_val_q[10] ),
    .S(_02441_),
    .X(_02464_));
 sky130_fd_sc_hd__and2_1 _19651_ (.A(_02445_),
    .B(_02464_),
    .X(_02465_));
 sky130_fd_sc_hd__clkbuf_1 _19652_ (.A(_02465_),
    .X(_01045_));
 sky130_fd_sc_hd__buf_4 _19653_ (.A(_02048_),
    .X(_02466_));
 sky130_fd_sc_hd__mux2_1 _19654_ (.A0(_01627_),
    .A1(\wfg_stim_sine_top.offset_val_q[11] ),
    .S(_02441_),
    .X(_02467_));
 sky130_fd_sc_hd__and2_1 _19655_ (.A(_02466_),
    .B(_02467_),
    .X(_02468_));
 sky130_fd_sc_hd__clkbuf_1 _19656_ (.A(_02468_),
    .X(_01046_));
 sky130_fd_sc_hd__mux2_1 _19657_ (.A0(_01630_),
    .A1(\wfg_stim_sine_top.offset_val_q[12] ),
    .S(_02441_),
    .X(_02469_));
 sky130_fd_sc_hd__and2_1 _19658_ (.A(_02466_),
    .B(_02469_),
    .X(_02470_));
 sky130_fd_sc_hd__clkbuf_1 _19659_ (.A(_02470_),
    .X(_01047_));
 sky130_fd_sc_hd__mux2_1 _19660_ (.A0(_01633_),
    .A1(\wfg_stim_sine_top.offset_val_q[13] ),
    .S(_02441_),
    .X(_02471_));
 sky130_fd_sc_hd__and2_1 _19661_ (.A(_02466_),
    .B(_02471_),
    .X(_02472_));
 sky130_fd_sc_hd__clkbuf_1 _19662_ (.A(_02472_),
    .X(_01048_));
 sky130_fd_sc_hd__mux2_1 _19663_ (.A0(_01636_),
    .A1(\wfg_stim_sine_top.offset_val_q[14] ),
    .S(_02441_),
    .X(_02473_));
 sky130_fd_sc_hd__and2_1 _19664_ (.A(_02466_),
    .B(_02473_),
    .X(_02474_));
 sky130_fd_sc_hd__clkbuf_1 _19665_ (.A(_02474_),
    .X(_01049_));
 sky130_fd_sc_hd__mux2_1 _19666_ (.A0(_01639_),
    .A1(\wfg_stim_sine_top.offset_val_q[15] ),
    .S(_02441_),
    .X(_02475_));
 sky130_fd_sc_hd__and2_1 _19667_ (.A(_02466_),
    .B(_02475_),
    .X(_02476_));
 sky130_fd_sc_hd__clkbuf_1 _19668_ (.A(_02476_),
    .X(_01050_));
 sky130_fd_sc_hd__mux2_1 _19669_ (.A0(net73),
    .A1(\wfg_stim_sine_top.offset_val_q[16] ),
    .S(_02441_),
    .X(_02477_));
 sky130_fd_sc_hd__and2_1 _19670_ (.A(_02466_),
    .B(_02477_),
    .X(_02478_));
 sky130_fd_sc_hd__clkbuf_1 _19671_ (.A(_02478_),
    .X(_01051_));
 sky130_fd_sc_hd__mux2_1 _19672_ (.A0(net74),
    .A1(\wfg_stim_sine_top.offset_val_q[17] ),
    .S(_02441_),
    .X(_02479_));
 sky130_fd_sc_hd__and2_1 _19673_ (.A(_02466_),
    .B(_02479_),
    .X(_02480_));
 sky130_fd_sc_hd__clkbuf_1 _19674_ (.A(_02480_),
    .X(_01052_));
 sky130_fd_sc_hd__inv_2 _19675_ (.A(_02287_),
    .Y(_00325_));
 sky130_fd_sc_hd__and3b_1 _19676_ (.A_N(\wfg_interconnect_top.wbs_ack_o ),
    .B(_01697_),
    .C(_02260_),
    .X(_02481_));
 sky130_fd_sc_hd__clkbuf_1 _19677_ (.A(_02481_),
    .X(_01053_));
 sky130_fd_sc_hd__inv_2 _19678_ (.A(_02287_),
    .Y(_00326_));
 sky130_fd_sc_hd__inv_2 _19679_ (.A(_02287_),
    .Y(_00327_));
 sky130_fd_sc_hd__inv_2 _19680_ (.A(_02287_),
    .Y(_00328_));
 sky130_fd_sc_hd__inv_2 _19681_ (.A(_02287_),
    .Y(_00329_));
 sky130_fd_sc_hd__inv_2 _19682_ (.A(_02287_),
    .Y(_00330_));
 sky130_fd_sc_hd__buf_6 _19683_ (.A(_02281_),
    .X(_02482_));
 sky130_fd_sc_hd__inv_2 _19684_ (.A(_02482_),
    .Y(_00331_));
 sky130_fd_sc_hd__inv_2 _19685_ (.A(_02482_),
    .Y(_00332_));
 sky130_fd_sc_hd__inv_2 _19686_ (.A(_02482_),
    .Y(_00333_));
 sky130_fd_sc_hd__inv_2 _19687_ (.A(_02482_),
    .Y(_00334_));
 sky130_fd_sc_hd__inv_2 _19688_ (.A(_02482_),
    .Y(_00335_));
 sky130_fd_sc_hd__inv_2 _19689_ (.A(_02482_),
    .Y(_00336_));
 sky130_fd_sc_hd__inv_2 _19690_ (.A(_02482_),
    .Y(_00337_));
 sky130_fd_sc_hd__inv_2 _19691_ (.A(_02482_),
    .Y(_00338_));
 sky130_fd_sc_hd__inv_2 _19692_ (.A(_02482_),
    .Y(_00339_));
 sky130_fd_sc_hd__inv_2 _19693_ (.A(_02482_),
    .Y(_00340_));
 sky130_fd_sc_hd__buf_4 _19694_ (.A(_02281_),
    .X(_02483_));
 sky130_fd_sc_hd__clkinv_4 _19695_ (.A(_02483_),
    .Y(_00341_));
 sky130_fd_sc_hd__inv_2 _19696_ (.A(_02483_),
    .Y(_00342_));
 sky130_fd_sc_hd__inv_2 _19697_ (.A(_02483_),
    .Y(_00343_));
 sky130_fd_sc_hd__inv_2 _19698_ (.A(_02483_),
    .Y(_00344_));
 sky130_fd_sc_hd__inv_2 _19699_ (.A(_02483_),
    .Y(_00345_));
 sky130_fd_sc_hd__inv_2 _19700_ (.A(_02483_),
    .Y(_00346_));
 sky130_fd_sc_hd__inv_2 _19701_ (.A(_02483_),
    .Y(_00347_));
 sky130_fd_sc_hd__inv_2 _19702_ (.A(_02483_),
    .Y(_00348_));
 sky130_fd_sc_hd__inv_2 _19703_ (.A(_02483_),
    .Y(_00349_));
 sky130_fd_sc_hd__inv_2 _19704_ (.A(_02483_),
    .Y(_00350_));
 sky130_fd_sc_hd__buf_4 _19705_ (.A(_02281_),
    .X(_02484_));
 sky130_fd_sc_hd__inv_2 _19706_ (.A(_02484_),
    .Y(_00351_));
 sky130_fd_sc_hd__inv_2 _19707_ (.A(_02484_),
    .Y(_00352_));
 sky130_fd_sc_hd__inv_2 _19708_ (.A(_02484_),
    .Y(_00353_));
 sky130_fd_sc_hd__inv_2 _19709_ (.A(_02484_),
    .Y(_00354_));
 sky130_fd_sc_hd__inv_2 _19710_ (.A(_02484_),
    .Y(_00355_));
 sky130_fd_sc_hd__inv_2 _19711_ (.A(_02484_),
    .Y(_00356_));
 sky130_fd_sc_hd__inv_2 _19712_ (.A(_02484_),
    .Y(_00357_));
 sky130_fd_sc_hd__inv_2 _19713_ (.A(_02484_),
    .Y(_00358_));
 sky130_fd_sc_hd__inv_2 _19714_ (.A(_02484_),
    .Y(_00359_));
 sky130_fd_sc_hd__inv_2 _19715_ (.A(_02484_),
    .Y(_00360_));
 sky130_fd_sc_hd__buf_4 _19716_ (.A(_02281_),
    .X(_02485_));
 sky130_fd_sc_hd__inv_2 _19717_ (.A(_02485_),
    .Y(_00361_));
 sky130_fd_sc_hd__inv_2 _19718_ (.A(_02485_),
    .Y(_00362_));
 sky130_fd_sc_hd__inv_2 _19719_ (.A(_02485_),
    .Y(_00363_));
 sky130_fd_sc_hd__inv_2 _19720_ (.A(_02485_),
    .Y(_00364_));
 sky130_fd_sc_hd__inv_2 _19721_ (.A(_02485_),
    .Y(_00365_));
 sky130_fd_sc_hd__inv_2 _19722_ (.A(_02485_),
    .Y(_00366_));
 sky130_fd_sc_hd__inv_2 _19723_ (.A(_02485_),
    .Y(_00367_));
 sky130_fd_sc_hd__inv_2 _19724_ (.A(_02485_),
    .Y(_00368_));
 sky130_fd_sc_hd__inv_2 _19725_ (.A(_02485_),
    .Y(_00369_));
 sky130_fd_sc_hd__inv_2 _19726_ (.A(_02485_),
    .Y(_00370_));
 sky130_fd_sc_hd__buf_6 _19727_ (.A(net98),
    .X(_02486_));
 sky130_fd_sc_hd__buf_6 _19728_ (.A(_02486_),
    .X(_02487_));
 sky130_fd_sc_hd__inv_2 _19729_ (.A(_02487_),
    .Y(_00371_));
 sky130_fd_sc_hd__inv_2 _19730_ (.A(_02487_),
    .Y(_00372_));
 sky130_fd_sc_hd__inv_2 _19731_ (.A(_02487_),
    .Y(_00373_));
 sky130_fd_sc_hd__inv_2 _19732_ (.A(_02487_),
    .Y(_00374_));
 sky130_fd_sc_hd__inv_2 _19733_ (.A(_02487_),
    .Y(_00375_));
 sky130_fd_sc_hd__inv_2 _19734_ (.A(_02487_),
    .Y(_00376_));
 sky130_fd_sc_hd__inv_2 _19735_ (.A(_02487_),
    .Y(_00377_));
 sky130_fd_sc_hd__inv_2 _19736_ (.A(_02487_),
    .Y(_00378_));
 sky130_fd_sc_hd__inv_2 _19737_ (.A(_02487_),
    .Y(_00379_));
 sky130_fd_sc_hd__inv_2 _19738_ (.A(_02487_),
    .Y(_00380_));
 sky130_fd_sc_hd__buf_4 _19739_ (.A(_02486_),
    .X(_02488_));
 sky130_fd_sc_hd__inv_2 _19740_ (.A(_02488_),
    .Y(_00381_));
 sky130_fd_sc_hd__inv_2 _19741_ (.A(_02488_),
    .Y(_00382_));
 sky130_fd_sc_hd__inv_2 _19742_ (.A(_02488_),
    .Y(_00383_));
 sky130_fd_sc_hd__inv_2 _19743_ (.A(_02488_),
    .Y(_00384_));
 sky130_fd_sc_hd__inv_2 _19744_ (.A(_02488_),
    .Y(_00385_));
 sky130_fd_sc_hd__inv_2 _19745_ (.A(_02488_),
    .Y(_00386_));
 sky130_fd_sc_hd__inv_2 _19746_ (.A(_02488_),
    .Y(_00387_));
 sky130_fd_sc_hd__inv_2 _19747_ (.A(_02488_),
    .Y(_00388_));
 sky130_fd_sc_hd__inv_2 _19748_ (.A(_02488_),
    .Y(_00389_));
 sky130_fd_sc_hd__inv_2 _19749_ (.A(_02488_),
    .Y(_00390_));
 sky130_fd_sc_hd__buf_4 _19750_ (.A(_02486_),
    .X(_02489_));
 sky130_fd_sc_hd__inv_2 _19751_ (.A(_02489_),
    .Y(_00391_));
 sky130_fd_sc_hd__inv_2 _19752_ (.A(_02489_),
    .Y(_00392_));
 sky130_fd_sc_hd__inv_2 _19753_ (.A(_02489_),
    .Y(_00393_));
 sky130_fd_sc_hd__inv_2 _19754_ (.A(_02489_),
    .Y(_00394_));
 sky130_fd_sc_hd__inv_2 _19755_ (.A(_02489_),
    .Y(_00395_));
 sky130_fd_sc_hd__inv_2 _19756_ (.A(_02489_),
    .Y(_00396_));
 sky130_fd_sc_hd__inv_2 _19757_ (.A(_02489_),
    .Y(_00397_));
 sky130_fd_sc_hd__inv_2 _19758_ (.A(_02489_),
    .Y(_00398_));
 sky130_fd_sc_hd__inv_2 _19759_ (.A(_02489_),
    .Y(_00399_));
 sky130_fd_sc_hd__inv_2 _19760_ (.A(_02489_),
    .Y(_00400_));
 sky130_fd_sc_hd__buf_6 _19761_ (.A(_02486_),
    .X(_02490_));
 sky130_fd_sc_hd__inv_2 _19762_ (.A(_02490_),
    .Y(_00401_));
 sky130_fd_sc_hd__inv_2 _19763_ (.A(_02490_),
    .Y(_00402_));
 sky130_fd_sc_hd__inv_2 _19764_ (.A(_02490_),
    .Y(_00403_));
 sky130_fd_sc_hd__inv_2 _19765_ (.A(_02490_),
    .Y(_00404_));
 sky130_fd_sc_hd__inv_2 _19766_ (.A(_02490_),
    .Y(_00405_));
 sky130_fd_sc_hd__and2_1 _19767_ (.A(_01706_),
    .B(_02260_),
    .X(_02491_));
 sky130_fd_sc_hd__nor2_1 _19768_ (.A(_02259_),
    .B(_01763_),
    .Y(_02492_));
 sky130_fd_sc_hd__inv_2 _19769_ (.A(_02492_),
    .Y(_02493_));
 sky130_fd_sc_hd__nor2_1 _19770_ (.A(_02259_),
    .B(_01959_),
    .Y(_02494_));
 sky130_fd_sc_hd__inv_2 _19771_ (.A(_02494_),
    .Y(_02495_));
 sky130_fd_sc_hd__nand2_1 _19772_ (.A(_01706_),
    .B(_02260_),
    .Y(_02496_));
 sky130_fd_sc_hd__a221o_1 _19773_ (.A1(\wfg_interconnect_top.driver1_select_q[0] ),
    .A2(_02492_),
    .B1(_02494_),
    .B2(\wfg_interconnect_top.driver0_select_q[0] ),
    .C1(_02496_),
    .X(_02497_));
 sky130_fd_sc_hd__a31o_1 _19774_ (.A1(\wfg_interconnect_top.ctrl_en_q ),
    .A2(_02493_),
    .A3(_02495_),
    .B1(_02497_),
    .X(_02498_));
 sky130_fd_sc_hd__o211a_1 _19775_ (.A1(\wfg_interconnect_top.wbs_dat_o[0] ),
    .A2(_02491_),
    .B1(_02498_),
    .C1(_02330_),
    .X(_01134_));
 sky130_fd_sc_hd__a221o_1 _19776_ (.A1(\wfg_interconnect_top.driver1_select_q[1] ),
    .A2(_02492_),
    .B1(_02494_),
    .B2(\wfg_interconnect_top.driver0_select_q[1] ),
    .C1(_02496_),
    .X(_02499_));
 sky130_fd_sc_hd__o211a_1 _19777_ (.A1(\wfg_interconnect_top.wbs_dat_o[1] ),
    .A2(_02491_),
    .B1(_02499_),
    .C1(_02330_),
    .X(_01135_));
 sky130_fd_sc_hd__nand4_4 _19778_ (.A(_01608_),
    .B(_01885_),
    .C(_02203_),
    .D(_01750_),
    .Y(_02500_));
 sky130_fd_sc_hd__o21ai_1 _19779_ (.A1(_01691_),
    .A2(_02500_),
    .B1(net111),
    .Y(_02501_));
 sky130_fd_sc_hd__o311a_1 _19780_ (.A1(_01660_),
    .A2(_01691_),
    .A3(_02500_),
    .B1(_02501_),
    .C1(_01600_),
    .X(_01136_));
 sky130_fd_sc_hd__or2_1 _19781_ (.A(_01756_),
    .B(_02500_),
    .X(_02502_));
 sky130_fd_sc_hd__buf_4 _19782_ (.A(_02502_),
    .X(_02503_));
 sky130_fd_sc_hd__mux2_1 _19783_ (.A0(net96),
    .A1(_04081_),
    .S(_02503_),
    .X(_02504_));
 sky130_fd_sc_hd__or2_1 _19784_ (.A(_01837_),
    .B(_02504_),
    .X(_02505_));
 sky130_fd_sc_hd__clkbuf_1 _19785_ (.A(_02505_),
    .X(_01137_));
 sky130_fd_sc_hd__buf_4 _19786_ (.A(_02503_),
    .X(_02506_));
 sky130_fd_sc_hd__mux2_1 _19787_ (.A0(_01620_),
    .A1(_03492_),
    .S(_02506_),
    .X(_02507_));
 sky130_fd_sc_hd__and2_1 _19788_ (.A(_02466_),
    .B(_02507_),
    .X(_02508_));
 sky130_fd_sc_hd__clkbuf_1 _19789_ (.A(_02508_),
    .X(_01138_));
 sky130_fd_sc_hd__mux2_1 _19790_ (.A0(_01624_),
    .A1(_03435_),
    .S(_02506_),
    .X(_02509_));
 sky130_fd_sc_hd__and2_1 _19791_ (.A(_02466_),
    .B(_02509_),
    .X(_02510_));
 sky130_fd_sc_hd__clkbuf_1 _19792_ (.A(_02510_),
    .X(_01139_));
 sky130_fd_sc_hd__mux2_1 _19793_ (.A0(_01627_),
    .A1(_02909_),
    .S(_02506_),
    .X(_02511_));
 sky130_fd_sc_hd__and2_1 _19794_ (.A(_02466_),
    .B(_02511_),
    .X(_02512_));
 sky130_fd_sc_hd__clkbuf_1 _19795_ (.A(_02512_),
    .X(_01140_));
 sky130_fd_sc_hd__clkbuf_2 _19796_ (.A(_02048_),
    .X(_02513_));
 sky130_fd_sc_hd__mux2_1 _19797_ (.A0(_01630_),
    .A1(_02897_),
    .S(_02506_),
    .X(_02514_));
 sky130_fd_sc_hd__and2_1 _19798_ (.A(_02513_),
    .B(_02514_),
    .X(_02515_));
 sky130_fd_sc_hd__clkbuf_1 _19799_ (.A(_02515_),
    .X(_01141_));
 sky130_fd_sc_hd__mux2_1 _19800_ (.A0(_01633_),
    .A1(_02895_),
    .S(_02506_),
    .X(_02516_));
 sky130_fd_sc_hd__and2_1 _19801_ (.A(_02513_),
    .B(_02516_),
    .X(_02517_));
 sky130_fd_sc_hd__clkbuf_1 _19802_ (.A(_02517_),
    .X(_01142_));
 sky130_fd_sc_hd__mux2_1 _19803_ (.A0(_01636_),
    .A1(_02918_),
    .S(_02506_),
    .X(_02518_));
 sky130_fd_sc_hd__and2_1 _19804_ (.A(_02513_),
    .B(_02518_),
    .X(_02519_));
 sky130_fd_sc_hd__clkbuf_1 _19805_ (.A(_02519_),
    .X(_01143_));
 sky130_fd_sc_hd__mux2_1 _19806_ (.A0(_01639_),
    .A1(_02923_),
    .S(_02506_),
    .X(_02520_));
 sky130_fd_sc_hd__and2_1 _19807_ (.A(_02513_),
    .B(_02520_),
    .X(_02521_));
 sky130_fd_sc_hd__clkbuf_1 _19808_ (.A(_02521_),
    .X(_01144_));
 sky130_fd_sc_hd__mux2_1 _19809_ (.A0(net73),
    .A1(_02921_),
    .S(_02506_),
    .X(_02522_));
 sky130_fd_sc_hd__and2_1 _19810_ (.A(_02513_),
    .B(_02522_),
    .X(_02523_));
 sky130_fd_sc_hd__clkbuf_1 _19811_ (.A(_02523_),
    .X(_01145_));
 sky130_fd_sc_hd__mux2_1 _19812_ (.A0(net74),
    .A1(_03142_),
    .S(_02506_),
    .X(_02524_));
 sky130_fd_sc_hd__and2_1 _19813_ (.A(_02513_),
    .B(_02524_),
    .X(_02525_));
 sky130_fd_sc_hd__clkbuf_1 _19814_ (.A(_02525_),
    .X(_01146_));
 sky130_fd_sc_hd__mux2_1 _19815_ (.A0(net75),
    .A1(_03302_),
    .S(_02506_),
    .X(_02526_));
 sky130_fd_sc_hd__and2_1 _19816_ (.A(_02513_),
    .B(_02526_),
    .X(_02527_));
 sky130_fd_sc_hd__clkbuf_1 _19817_ (.A(_02527_),
    .X(_01147_));
 sky130_fd_sc_hd__buf_6 _19818_ (.A(_02503_),
    .X(_02528_));
 sky130_fd_sc_hd__mux2_1 _19819_ (.A0(net76),
    .A1(_02969_),
    .S(_02528_),
    .X(_02529_));
 sky130_fd_sc_hd__and2_1 _19820_ (.A(_02513_),
    .B(_02529_),
    .X(_02530_));
 sky130_fd_sc_hd__clkbuf_1 _19821_ (.A(_02530_),
    .X(_01148_));
 sky130_fd_sc_hd__mux2_1 _19822_ (.A0(net78),
    .A1(_02950_),
    .S(_02528_),
    .X(_02531_));
 sky130_fd_sc_hd__and2_1 _19823_ (.A(_02513_),
    .B(_02531_),
    .X(_02532_));
 sky130_fd_sc_hd__clkbuf_1 _19824_ (.A(_02532_),
    .X(_01149_));
 sky130_fd_sc_hd__mux2_1 _19825_ (.A0(net79),
    .A1(_02986_),
    .S(_02528_),
    .X(_02533_));
 sky130_fd_sc_hd__and2_1 _19826_ (.A(_02513_),
    .B(_02533_),
    .X(_02534_));
 sky130_fd_sc_hd__clkbuf_1 _19827_ (.A(_02534_),
    .X(_01150_));
 sky130_fd_sc_hd__clkbuf_4 _19828_ (.A(_01588_),
    .X(_02535_));
 sky130_fd_sc_hd__mux2_2 _19829_ (.A0(net80),
    .A1(_02988_),
    .S(_02528_),
    .X(_02536_));
 sky130_fd_sc_hd__and2_1 _19830_ (.A(_02535_),
    .B(_02536_),
    .X(_02537_));
 sky130_fd_sc_hd__clkbuf_1 _19831_ (.A(_02537_),
    .X(_01151_));
 sky130_fd_sc_hd__mux2_2 _19832_ (.A0(net81),
    .A1(_03016_),
    .S(_02528_),
    .X(_02538_));
 sky130_fd_sc_hd__and2_1 _19833_ (.A(_02535_),
    .B(_02538_),
    .X(_02539_));
 sky130_fd_sc_hd__clkbuf_1 _19834_ (.A(_02539_),
    .X(_01152_));
 sky130_fd_sc_hd__mux2_1 _19835_ (.A0(_01884_),
    .A1(\wfg_stim_mem_top.cfg_inc_q[0] ),
    .S(_02503_),
    .X(_02540_));
 sky130_fd_sc_hd__or2_1 _19836_ (.A(_01837_),
    .B(_02540_),
    .X(_02541_));
 sky130_fd_sc_hd__clkbuf_1 _19837_ (.A(_02541_),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_1 _19838_ (.A0(net77),
    .A1(\wfg_stim_mem_top.cfg_inc_q[1] ),
    .S(_02528_),
    .X(_02542_));
 sky130_fd_sc_hd__and2_1 _19839_ (.A(_02535_),
    .B(_02542_),
    .X(_02543_));
 sky130_fd_sc_hd__clkbuf_1 _19840_ (.A(_02543_),
    .X(_01154_));
 sky130_fd_sc_hd__mux2_1 _19841_ (.A0(net88),
    .A1(\wfg_stim_mem_top.cfg_inc_q[2] ),
    .S(_02528_),
    .X(_02544_));
 sky130_fd_sc_hd__and2_1 _19842_ (.A(_02535_),
    .B(_02544_),
    .X(_02545_));
 sky130_fd_sc_hd__clkbuf_1 _19843_ (.A(_02545_),
    .X(_01155_));
 sky130_fd_sc_hd__mux2_1 _19844_ (.A0(net91),
    .A1(\wfg_stim_mem_top.cfg_inc_q[3] ),
    .S(_02528_),
    .X(_02546_));
 sky130_fd_sc_hd__and2_1 _19845_ (.A(_02535_),
    .B(_02546_),
    .X(_02547_));
 sky130_fd_sc_hd__clkbuf_1 _19846_ (.A(_02547_),
    .X(_01156_));
 sky130_fd_sc_hd__mux2_1 _19847_ (.A0(net92),
    .A1(\wfg_stim_mem_top.cfg_inc_q[4] ),
    .S(_02528_),
    .X(_02548_));
 sky130_fd_sc_hd__and2_1 _19848_ (.A(_02535_),
    .B(_02548_),
    .X(_02549_));
 sky130_fd_sc_hd__clkbuf_1 _19849_ (.A(_02549_),
    .X(_01157_));
 sky130_fd_sc_hd__mux2_1 _19850_ (.A0(net93),
    .A1(\wfg_stim_mem_top.cfg_inc_q[5] ),
    .S(_02528_),
    .X(_02550_));
 sky130_fd_sc_hd__and2_1 _19851_ (.A(_02535_),
    .B(_02550_),
    .X(_02551_));
 sky130_fd_sc_hd__clkbuf_1 _19852_ (.A(_02551_),
    .X(_01158_));
 sky130_fd_sc_hd__mux2_1 _19853_ (.A0(net94),
    .A1(\wfg_stim_mem_top.cfg_inc_q[6] ),
    .S(_02503_),
    .X(_02552_));
 sky130_fd_sc_hd__and2_1 _19854_ (.A(_02535_),
    .B(_02552_),
    .X(_02553_));
 sky130_fd_sc_hd__clkbuf_1 _19855_ (.A(_02553_),
    .X(_01159_));
 sky130_fd_sc_hd__mux2_1 _19856_ (.A0(net95),
    .A1(\wfg_stim_mem_top.cfg_inc_q[7] ),
    .S(_02503_),
    .X(_02554_));
 sky130_fd_sc_hd__and2_1 _19857_ (.A(_02535_),
    .B(_02554_),
    .X(_02555_));
 sky130_fd_sc_hd__clkbuf_1 _19858_ (.A(_02555_),
    .X(_01160_));
 sky130_fd_sc_hd__or2_1 _19859_ (.A(_01762_),
    .B(_02500_),
    .X(_02556_));
 sky130_fd_sc_hd__buf_2 _19860_ (.A(_02556_),
    .X(_02557_));
 sky130_fd_sc_hd__buf_4 _19861_ (.A(_02557_),
    .X(_02558_));
 sky130_fd_sc_hd__mux2_1 _19862_ (.A0(_01884_),
    .A1(\wfg_stim_mem_top.end_val_q[0] ),
    .S(_02558_),
    .X(_02559_));
 sky130_fd_sc_hd__and2_1 _19863_ (.A(_02535_),
    .B(_02559_),
    .X(_02560_));
 sky130_fd_sc_hd__clkbuf_1 _19864_ (.A(_02560_),
    .X(_01161_));
 sky130_fd_sc_hd__buf_2 _19865_ (.A(_01588_),
    .X(_02561_));
 sky130_fd_sc_hd__mux2_1 _19866_ (.A0(net77),
    .A1(\wfg_stim_mem_top.end_val_q[1] ),
    .S(_02558_),
    .X(_02562_));
 sky130_fd_sc_hd__and2_1 _19867_ (.A(_02561_),
    .B(_02562_),
    .X(_02563_));
 sky130_fd_sc_hd__clkbuf_1 _19868_ (.A(_02563_),
    .X(_01162_));
 sky130_fd_sc_hd__mux2_1 _19869_ (.A0(net88),
    .A1(\wfg_stim_mem_top.end_val_q[2] ),
    .S(_02558_),
    .X(_02564_));
 sky130_fd_sc_hd__and2_1 _19870_ (.A(_02561_),
    .B(_02564_),
    .X(_02565_));
 sky130_fd_sc_hd__clkbuf_1 _19871_ (.A(_02565_),
    .X(_01163_));
 sky130_fd_sc_hd__mux2_1 _19872_ (.A0(net91),
    .A1(\wfg_stim_mem_top.end_val_q[3] ),
    .S(_02558_),
    .X(_02566_));
 sky130_fd_sc_hd__and2_1 _19873_ (.A(_02561_),
    .B(_02566_),
    .X(_02567_));
 sky130_fd_sc_hd__clkbuf_1 _19874_ (.A(_02567_),
    .X(_01164_));
 sky130_fd_sc_hd__mux2_1 _19875_ (.A0(net92),
    .A1(\wfg_stim_mem_top.end_val_q[4] ),
    .S(_02558_),
    .X(_02568_));
 sky130_fd_sc_hd__and2_1 _19876_ (.A(_02561_),
    .B(_02568_),
    .X(_02569_));
 sky130_fd_sc_hd__clkbuf_1 _19877_ (.A(_02569_),
    .X(_01165_));
 sky130_fd_sc_hd__mux2_1 _19878_ (.A0(net93),
    .A1(\wfg_stim_mem_top.end_val_q[5] ),
    .S(_02558_),
    .X(_02570_));
 sky130_fd_sc_hd__and2_1 _19879_ (.A(_02561_),
    .B(_02570_),
    .X(_02571_));
 sky130_fd_sc_hd__clkbuf_1 _19880_ (.A(_02571_),
    .X(_01166_));
 sky130_fd_sc_hd__mux2_1 _19881_ (.A0(net94),
    .A1(\wfg_stim_mem_top.end_val_q[6] ),
    .S(_02558_),
    .X(_02572_));
 sky130_fd_sc_hd__and2_1 _19882_ (.A(_02561_),
    .B(_02572_),
    .X(_02573_));
 sky130_fd_sc_hd__clkbuf_1 _19883_ (.A(_02573_),
    .X(_01167_));
 sky130_fd_sc_hd__mux2_1 _19884_ (.A0(net95),
    .A1(\wfg_stim_mem_top.end_val_q[7] ),
    .S(_02558_),
    .X(_02574_));
 sky130_fd_sc_hd__and2_1 _19885_ (.A(_02561_),
    .B(_02574_),
    .X(_02575_));
 sky130_fd_sc_hd__clkbuf_1 _19886_ (.A(_02575_),
    .X(_01168_));
 sky130_fd_sc_hd__mux2_1 _19887_ (.A0(_01601_),
    .A1(\wfg_stim_mem_top.end_val_q[8] ),
    .S(_02558_),
    .X(_02576_));
 sky130_fd_sc_hd__and2_1 _19888_ (.A(_02561_),
    .B(_02576_),
    .X(_02577_));
 sky130_fd_sc_hd__clkbuf_1 _19889_ (.A(_02577_),
    .X(_01169_));
 sky130_fd_sc_hd__mux2_1 _19890_ (.A0(net97),
    .A1(\wfg_stim_mem_top.end_val_q[9] ),
    .S(_02558_),
    .X(_02578_));
 sky130_fd_sc_hd__and2_1 _19891_ (.A(_02561_),
    .B(_02578_),
    .X(_02579_));
 sky130_fd_sc_hd__clkbuf_1 _19892_ (.A(_02579_),
    .X(_01170_));
 sky130_fd_sc_hd__mux2_1 _19893_ (.A0(net67),
    .A1(\wfg_stim_mem_top.end_val_q[10] ),
    .S(_02557_),
    .X(_02580_));
 sky130_fd_sc_hd__and2_1 _19894_ (.A(_02561_),
    .B(_02580_),
    .X(_02581_));
 sky130_fd_sc_hd__clkbuf_1 _19895_ (.A(_02581_),
    .X(_01171_));
 sky130_fd_sc_hd__clkbuf_4 _19896_ (.A(_01588_),
    .X(_02582_));
 sky130_fd_sc_hd__mux2_1 _19897_ (.A0(net68),
    .A1(\wfg_stim_mem_top.end_val_q[11] ),
    .S(_02557_),
    .X(_02583_));
 sky130_fd_sc_hd__and2_1 _19898_ (.A(_02582_),
    .B(_02583_),
    .X(_02584_));
 sky130_fd_sc_hd__clkbuf_1 _19899_ (.A(_02584_),
    .X(_01172_));
 sky130_fd_sc_hd__mux2_1 _19900_ (.A0(_01630_),
    .A1(\wfg_stim_mem_top.end_val_q[12] ),
    .S(_02557_),
    .X(_02585_));
 sky130_fd_sc_hd__and2_1 _19901_ (.A(_02582_),
    .B(_02585_),
    .X(_02586_));
 sky130_fd_sc_hd__clkbuf_1 _19902_ (.A(_02586_),
    .X(_01173_));
 sky130_fd_sc_hd__mux2_1 _19903_ (.A0(net70),
    .A1(\wfg_stim_mem_top.end_val_q[13] ),
    .S(_02557_),
    .X(_02587_));
 sky130_fd_sc_hd__and2_1 _19904_ (.A(_02582_),
    .B(_02587_),
    .X(_02588_));
 sky130_fd_sc_hd__clkbuf_1 _19905_ (.A(_02588_),
    .X(_01174_));
 sky130_fd_sc_hd__mux2_1 _19906_ (.A0(_01636_),
    .A1(\wfg_stim_mem_top.end_val_q[14] ),
    .S(_02557_),
    .X(_02589_));
 sky130_fd_sc_hd__and2_1 _19907_ (.A(_02582_),
    .B(_02589_),
    .X(_02590_));
 sky130_fd_sc_hd__clkbuf_1 _19908_ (.A(_02590_),
    .X(_01175_));
 sky130_fd_sc_hd__mux2_1 _19909_ (.A0(net72),
    .A1(\wfg_stim_mem_top.end_val_q[15] ),
    .S(_02557_),
    .X(_02591_));
 sky130_fd_sc_hd__and2_1 _19910_ (.A(_02582_),
    .B(_02591_),
    .X(_02592_));
 sky130_fd_sc_hd__clkbuf_1 _19911_ (.A(_02592_),
    .X(_01176_));
 sky130_fd_sc_hd__or2_1 _19912_ (.A(_01604_),
    .B(_02500_),
    .X(_02593_));
 sky130_fd_sc_hd__clkbuf_4 _19913_ (.A(_02593_),
    .X(_02594_));
 sky130_fd_sc_hd__clkbuf_4 _19914_ (.A(_02594_),
    .X(_02595_));
 sky130_fd_sc_hd__mux2_1 _19915_ (.A0(_01884_),
    .A1(\wfg_stim_mem_top.start_val_q[0] ),
    .S(_02595_),
    .X(_02596_));
 sky130_fd_sc_hd__and2_1 _19916_ (.A(_02582_),
    .B(_02596_),
    .X(_02597_));
 sky130_fd_sc_hd__clkbuf_1 _19917_ (.A(_02597_),
    .X(_01177_));
 sky130_fd_sc_hd__nand2_1 _19918_ (.A(_06300_),
    .B(_02595_),
    .Y(_02598_));
 sky130_fd_sc_hd__o211a_1 _19919_ (.A1(_01663_),
    .A2(_02595_),
    .B1(_02598_),
    .C1(_02330_),
    .X(_01178_));
 sky130_fd_sc_hd__mux2_1 _19920_ (.A0(net88),
    .A1(\wfg_stim_mem_top.start_val_q[2] ),
    .S(_02595_),
    .X(_02599_));
 sky130_fd_sc_hd__and2_1 _19921_ (.A(_02582_),
    .B(_02599_),
    .X(_02600_));
 sky130_fd_sc_hd__clkbuf_1 _19922_ (.A(_02600_),
    .X(_01179_));
 sky130_fd_sc_hd__mux2_1 _19923_ (.A0(net91),
    .A1(\wfg_stim_mem_top.start_val_q[3] ),
    .S(_02595_),
    .X(_02601_));
 sky130_fd_sc_hd__and2_1 _19924_ (.A(_02582_),
    .B(_02601_),
    .X(_02602_));
 sky130_fd_sc_hd__clkbuf_1 _19925_ (.A(_02602_),
    .X(_01180_));
 sky130_fd_sc_hd__mux2_1 _19926_ (.A0(net92),
    .A1(\wfg_stim_mem_top.start_val_q[4] ),
    .S(_02595_),
    .X(_02603_));
 sky130_fd_sc_hd__and2_1 _19927_ (.A(_02582_),
    .B(_02603_),
    .X(_02604_));
 sky130_fd_sc_hd__clkbuf_1 _19928_ (.A(_02604_),
    .X(_01181_));
 sky130_fd_sc_hd__mux2_1 _19929_ (.A0(net93),
    .A1(\wfg_stim_mem_top.start_val_q[5] ),
    .S(_02595_),
    .X(_02605_));
 sky130_fd_sc_hd__and2_1 _19930_ (.A(_02582_),
    .B(_02605_),
    .X(_02606_));
 sky130_fd_sc_hd__clkbuf_1 _19931_ (.A(_02606_),
    .X(_01182_));
 sky130_fd_sc_hd__buf_2 _19932_ (.A(_01588_),
    .X(_02607_));
 sky130_fd_sc_hd__mux2_1 _19933_ (.A0(net94),
    .A1(\wfg_stim_mem_top.start_val_q[6] ),
    .S(_02595_),
    .X(_02608_));
 sky130_fd_sc_hd__and2_1 _19934_ (.A(_02607_),
    .B(_02608_),
    .X(_02609_));
 sky130_fd_sc_hd__clkbuf_1 _19935_ (.A(_02609_),
    .X(_01183_));
 sky130_fd_sc_hd__mux2_1 _19936_ (.A0(net95),
    .A1(\wfg_stim_mem_top.start_val_q[7] ),
    .S(_02595_),
    .X(_02610_));
 sky130_fd_sc_hd__and2_1 _19937_ (.A(_02607_),
    .B(_02610_),
    .X(_02611_));
 sky130_fd_sc_hd__clkbuf_1 _19938_ (.A(_02611_),
    .X(_01184_));
 sky130_fd_sc_hd__mux2_1 _19939_ (.A0(net96),
    .A1(\wfg_stim_mem_top.start_val_q[8] ),
    .S(_02595_),
    .X(_02612_));
 sky130_fd_sc_hd__and2_1 _19940_ (.A(_02607_),
    .B(_02612_),
    .X(_02613_));
 sky130_fd_sc_hd__clkbuf_1 _19941_ (.A(_02613_),
    .X(_01185_));
 sky130_fd_sc_hd__mux2_1 _19942_ (.A0(net97),
    .A1(\wfg_stim_mem_top.start_val_q[9] ),
    .S(_02594_),
    .X(_02614_));
 sky130_fd_sc_hd__and2_1 _19943_ (.A(_02607_),
    .B(_02614_),
    .X(_02615_));
 sky130_fd_sc_hd__clkbuf_1 _19944_ (.A(_02615_),
    .X(_01186_));
 sky130_fd_sc_hd__mux2_1 _19945_ (.A0(net67),
    .A1(\wfg_stim_mem_top.start_val_q[10] ),
    .S(_02594_),
    .X(_02616_));
 sky130_fd_sc_hd__and2_1 _19946_ (.A(_02607_),
    .B(_02616_),
    .X(_02617_));
 sky130_fd_sc_hd__clkbuf_1 _19947_ (.A(_02617_),
    .X(_01187_));
 sky130_fd_sc_hd__mux2_1 _19948_ (.A0(net68),
    .A1(\wfg_stim_mem_top.start_val_q[11] ),
    .S(_02594_),
    .X(_02618_));
 sky130_fd_sc_hd__and2_1 _19949_ (.A(_02607_),
    .B(_02618_),
    .X(_02619_));
 sky130_fd_sc_hd__clkbuf_1 _19950_ (.A(_02619_),
    .X(_01188_));
 sky130_fd_sc_hd__mux2_1 _19951_ (.A0(net69),
    .A1(\wfg_stim_mem_top.start_val_q[12] ),
    .S(_02594_),
    .X(_02620_));
 sky130_fd_sc_hd__and2_1 _19952_ (.A(_02607_),
    .B(_02620_),
    .X(_02621_));
 sky130_fd_sc_hd__clkbuf_1 _19953_ (.A(_02621_),
    .X(_01189_));
 sky130_fd_sc_hd__mux2_1 _19954_ (.A0(net70),
    .A1(\wfg_stim_mem_top.start_val_q[13] ),
    .S(_02594_),
    .X(_02622_));
 sky130_fd_sc_hd__and2_1 _19955_ (.A(_02607_),
    .B(_02622_),
    .X(_02623_));
 sky130_fd_sc_hd__clkbuf_1 _19956_ (.A(_02623_),
    .X(_01190_));
 sky130_fd_sc_hd__mux2_1 _19957_ (.A0(net71),
    .A1(\wfg_stim_mem_top.start_val_q[14] ),
    .S(_02594_),
    .X(_02624_));
 sky130_fd_sc_hd__and2_1 _19958_ (.A(_02607_),
    .B(_02624_),
    .X(_02625_));
 sky130_fd_sc_hd__clkbuf_1 _19959_ (.A(_02625_),
    .X(_01191_));
 sky130_fd_sc_hd__mux2_1 _19960_ (.A0(net72),
    .A1(\wfg_stim_mem_top.start_val_q[15] ),
    .S(_02594_),
    .X(_02626_));
 sky130_fd_sc_hd__and2_1 _19961_ (.A(_02607_),
    .B(_02626_),
    .X(_02627_));
 sky130_fd_sc_hd__clkbuf_1 _19962_ (.A(_02627_),
    .X(_01192_));
 sky130_fd_sc_hd__inv_2 _19963_ (.A(_02490_),
    .Y(_00406_));
 sky130_fd_sc_hd__inv_2 _19964_ (.A(_02490_),
    .Y(_00407_));
 sky130_fd_sc_hd__inv_2 _19965_ (.A(_02490_),
    .Y(_00408_));
 sky130_fd_sc_hd__inv_2 _19966_ (.A(_02490_),
    .Y(_00409_));
 sky130_fd_sc_hd__inv_2 _19967_ (.A(_02490_),
    .Y(_00410_));
 sky130_fd_sc_hd__and4b_1 _19968_ (.A_N(\wfg_drive_pat_top.wbs_ack_o ),
    .B(_01453_),
    .C(_01750_),
    .D(_01697_),
    .X(_02628_));
 sky130_fd_sc_hd__clkbuf_1 _19969_ (.A(_02628_),
    .X(_01193_));
 sky130_fd_sc_hd__buf_4 _19970_ (.A(_02486_),
    .X(_02629_));
 sky130_fd_sc_hd__inv_2 _19971_ (.A(_02629_),
    .Y(_00411_));
 sky130_fd_sc_hd__inv_2 _19972_ (.A(_02629_),
    .Y(_00412_));
 sky130_fd_sc_hd__inv_2 _19973_ (.A(_02629_),
    .Y(_00413_));
 sky130_fd_sc_hd__inv_2 _19974_ (.A(_02629_),
    .Y(_00414_));
 sky130_fd_sc_hd__inv_2 _19975_ (.A(_02629_),
    .Y(_00415_));
 sky130_fd_sc_hd__inv_2 _19976_ (.A(_02629_),
    .Y(_00416_));
 sky130_fd_sc_hd__inv_2 _19977_ (.A(_02629_),
    .Y(_00417_));
 sky130_fd_sc_hd__inv_2 _19978_ (.A(_02629_),
    .Y(_00418_));
 sky130_fd_sc_hd__inv_2 _19979_ (.A(_02629_),
    .Y(_00419_));
 sky130_fd_sc_hd__inv_2 _19980_ (.A(_02629_),
    .Y(_00420_));
 sky130_fd_sc_hd__buf_6 _19981_ (.A(_02486_),
    .X(_02630_));
 sky130_fd_sc_hd__inv_2 _19982_ (.A(_02630_),
    .Y(_00421_));
 sky130_fd_sc_hd__inv_2 _19983_ (.A(_02630_),
    .Y(_00422_));
 sky130_fd_sc_hd__inv_2 _19984_ (.A(_02630_),
    .Y(_00423_));
 sky130_fd_sc_hd__inv_2 _19985_ (.A(_02630_),
    .Y(_00424_));
 sky130_fd_sc_hd__inv_2 _19986_ (.A(_02630_),
    .Y(_00425_));
 sky130_fd_sc_hd__inv_2 _19987_ (.A(_02630_),
    .Y(_00426_));
 sky130_fd_sc_hd__inv_2 _19988_ (.A(_02630_),
    .Y(_00427_));
 sky130_fd_sc_hd__inv_2 _19989_ (.A(_02630_),
    .Y(_00428_));
 sky130_fd_sc_hd__inv_2 _19990_ (.A(_02630_),
    .Y(_00429_));
 sky130_fd_sc_hd__inv_2 _19991_ (.A(_02630_),
    .Y(_00430_));
 sky130_fd_sc_hd__clkbuf_8 _19992_ (.A(_02486_),
    .X(_02631_));
 sky130_fd_sc_hd__inv_2 _19993_ (.A(_02631_),
    .Y(_00431_));
 sky130_fd_sc_hd__inv_2 _19994_ (.A(_02631_),
    .Y(_00432_));
 sky130_fd_sc_hd__inv_2 _19995_ (.A(_02631_),
    .Y(_00433_));
 sky130_fd_sc_hd__inv_2 _19996_ (.A(_02631_),
    .Y(_00434_));
 sky130_fd_sc_hd__inv_2 _19997_ (.A(_02631_),
    .Y(_00435_));
 sky130_fd_sc_hd__inv_2 _19998_ (.A(_02631_),
    .Y(_00436_));
 sky130_fd_sc_hd__inv_2 _19999_ (.A(_02631_),
    .Y(_00437_));
 sky130_fd_sc_hd__inv_2 _20000_ (.A(_02631_),
    .Y(_00438_));
 sky130_fd_sc_hd__inv_2 _20001_ (.A(_02631_),
    .Y(_00439_));
 sky130_fd_sc_hd__inv_2 _20002_ (.A(_02631_),
    .Y(_00440_));
 sky130_fd_sc_hd__buf_4 _20003_ (.A(_02486_),
    .X(_02632_));
 sky130_fd_sc_hd__inv_2 _20004_ (.A(_02632_),
    .Y(_00441_));
 sky130_fd_sc_hd__inv_2 _20005_ (.A(_02632_),
    .Y(_00442_));
 sky130_fd_sc_hd__inv_2 _20006_ (.A(_02632_),
    .Y(_00443_));
 sky130_fd_sc_hd__inv_2 _20007_ (.A(_02632_),
    .Y(_00444_));
 sky130_fd_sc_hd__inv_2 _20008_ (.A(_02632_),
    .Y(_00445_));
 sky130_fd_sc_hd__inv_2 _20009_ (.A(_02632_),
    .Y(_00446_));
 sky130_fd_sc_hd__inv_2 _20010_ (.A(_02632_),
    .Y(_00447_));
 sky130_fd_sc_hd__inv_2 _20011_ (.A(_02632_),
    .Y(_00448_));
 sky130_fd_sc_hd__inv_2 _20012_ (.A(_02632_),
    .Y(_00449_));
 sky130_fd_sc_hd__inv_2 _20013_ (.A(_02632_),
    .Y(_00450_));
 sky130_fd_sc_hd__buf_4 _20014_ (.A(_02486_),
    .X(_02633_));
 sky130_fd_sc_hd__inv_2 _20015_ (.A(_02633_),
    .Y(_00451_));
 sky130_fd_sc_hd__inv_2 _20016_ (.A(_02633_),
    .Y(_00452_));
 sky130_fd_sc_hd__inv_2 _20017_ (.A(_02633_),
    .Y(_00453_));
 sky130_fd_sc_hd__inv_2 _20018_ (.A(_02633_),
    .Y(_00454_));
 sky130_fd_sc_hd__inv_2 _20019_ (.A(_02633_),
    .Y(_00455_));
 sky130_fd_sc_hd__inv_2 _20020_ (.A(_02633_),
    .Y(_00456_));
 sky130_fd_sc_hd__inv_2 _20021_ (.A(_02633_),
    .Y(_00457_));
 sky130_fd_sc_hd__inv_2 _20022_ (.A(_02633_),
    .Y(_00458_));
 sky130_fd_sc_hd__inv_2 _20023_ (.A(_02633_),
    .Y(_00459_));
 sky130_fd_sc_hd__inv_2 _20024_ (.A(_02633_),
    .Y(_00460_));
 sky130_fd_sc_hd__buf_6 _20025_ (.A(_02486_),
    .X(_02634_));
 sky130_fd_sc_hd__inv_2 _20026_ (.A(_02634_),
    .Y(_00461_));
 sky130_fd_sc_hd__inv_2 _20027_ (.A(_02634_),
    .Y(_00462_));
 sky130_fd_sc_hd__inv_2 _20028_ (.A(_02634_),
    .Y(_00463_));
 sky130_fd_sc_hd__inv_2 _20029_ (.A(_02634_),
    .Y(_00464_));
 sky130_fd_sc_hd__inv_2 _20030_ (.A(_02634_),
    .Y(_00465_));
 sky130_fd_sc_hd__inv_2 _20031_ (.A(_02634_),
    .Y(_00466_));
 sky130_fd_sc_hd__inv_2 _20032_ (.A(_02634_),
    .Y(_00467_));
 sky130_fd_sc_hd__inv_2 _20033_ (.A(_02634_),
    .Y(_00468_));
 sky130_fd_sc_hd__inv_2 _20034_ (.A(_02634_),
    .Y(_00469_));
 sky130_fd_sc_hd__inv_2 _20035_ (.A(_02634_),
    .Y(_00470_));
 sky130_fd_sc_hd__inv_2 _20036_ (.A(_01591_),
    .Y(_00471_));
 sky130_fd_sc_hd__or2_2 _20037_ (.A(_01688_),
    .B(_01713_),
    .X(_02635_));
 sky130_fd_sc_hd__buf_2 _20038_ (.A(_02635_),
    .X(_02636_));
 sky130_fd_sc_hd__nor2_2 _20039_ (.A(_01687_),
    .B(_01709_),
    .Y(_02637_));
 sky130_fd_sc_hd__or3_1 _20040_ (.A(\wfg_core_top.cfg_sync_q[0] ),
    .B(_01687_),
    .C(_01709_),
    .X(_02638_));
 sky130_fd_sc_hd__nor2_2 _20041_ (.A(_01688_),
    .B(_01713_),
    .Y(_02639_));
 sky130_fd_sc_hd__o211a_1 _20042_ (.A1(\wfg_core_top.active_o ),
    .A2(_02637_),
    .B1(_02638_),
    .C1(_02639_),
    .X(_02640_));
 sky130_fd_sc_hd__a21oi_1 _20043_ (.A1(\wfg_core_top.wbs_dat_o[0] ),
    .A2(_02636_),
    .B1(_02640_),
    .Y(_02641_));
 sky130_fd_sc_hd__nor2_1 _20044_ (.A(_01591_),
    .B(_02641_),
    .Y(_01254_));
 sky130_fd_sc_hd__buf_2 _20045_ (.A(_02639_),
    .X(_02642_));
 sky130_fd_sc_hd__buf_2 _20046_ (.A(_02637_),
    .X(_02643_));
 sky130_fd_sc_hd__a21o_1 _20047_ (.A1(\wfg_core_top.cfg_sync_q[1] ),
    .A2(_02643_),
    .B1(_02636_),
    .X(_02644_));
 sky130_fd_sc_hd__o211a_1 _20048_ (.A1(\wfg_core_top.wbs_dat_o[1] ),
    .A2(_02642_),
    .B1(_02644_),
    .C1(_02330_),
    .X(_01255_));
 sky130_fd_sc_hd__a21o_1 _20049_ (.A1(\wfg_core_top.cfg_sync_q[2] ),
    .A2(_02643_),
    .B1(_02636_),
    .X(_02645_));
 sky130_fd_sc_hd__o211a_1 _20050_ (.A1(\wfg_core_top.wbs_dat_o[2] ),
    .A2(_02642_),
    .B1(_02645_),
    .C1(_02330_),
    .X(_01256_));
 sky130_fd_sc_hd__a21o_1 _20051_ (.A1(\wfg_core_top.cfg_sync_q[3] ),
    .A2(_02643_),
    .B1(_02636_),
    .X(_02646_));
 sky130_fd_sc_hd__buf_2 _20052_ (.A(_01589_),
    .X(_02647_));
 sky130_fd_sc_hd__o211a_1 _20053_ (.A1(\wfg_core_top.wbs_dat_o[3] ),
    .A2(_02642_),
    .B1(_02646_),
    .C1(_02647_),
    .X(_01257_));
 sky130_fd_sc_hd__a21o_1 _20054_ (.A1(\wfg_core_top.cfg_sync_q[4] ),
    .A2(_02643_),
    .B1(_02636_),
    .X(_02648_));
 sky130_fd_sc_hd__o211a_1 _20055_ (.A1(\wfg_core_top.wbs_dat_o[4] ),
    .A2(_02642_),
    .B1(_02648_),
    .C1(_02647_),
    .X(_01258_));
 sky130_fd_sc_hd__a21o_1 _20056_ (.A1(\wfg_core_top.cfg_sync_q[5] ),
    .A2(_02643_),
    .B1(_02636_),
    .X(_02649_));
 sky130_fd_sc_hd__o211a_1 _20057_ (.A1(\wfg_core_top.wbs_dat_o[5] ),
    .A2(_02642_),
    .B1(_02649_),
    .C1(_02647_),
    .X(_01259_));
 sky130_fd_sc_hd__a21o_1 _20058_ (.A1(\wfg_core_top.cfg_sync_q[6] ),
    .A2(_02643_),
    .B1(_02636_),
    .X(_02650_));
 sky130_fd_sc_hd__o211a_1 _20059_ (.A1(\wfg_core_top.wbs_dat_o[6] ),
    .A2(_02642_),
    .B1(_02650_),
    .C1(_02647_),
    .X(_01260_));
 sky130_fd_sc_hd__a21o_1 _20060_ (.A1(\wfg_core_top.cfg_sync_q[7] ),
    .A2(_02643_),
    .B1(_02636_),
    .X(_02651_));
 sky130_fd_sc_hd__o211a_1 _20061_ (.A1(\wfg_core_top.wbs_dat_o[7] ),
    .A2(_02642_),
    .B1(_02651_),
    .C1(_02647_),
    .X(_01261_));
 sky130_fd_sc_hd__a21o_1 _20062_ (.A1(\wfg_core_top.cfg_subcycle_q[8] ),
    .A2(_02643_),
    .B1(_02636_),
    .X(_02652_));
 sky130_fd_sc_hd__o211a_1 _20063_ (.A1(\wfg_core_top.wbs_dat_o[8] ),
    .A2(_02642_),
    .B1(_02652_),
    .C1(_02647_),
    .X(_01262_));
 sky130_fd_sc_hd__a21o_1 _20064_ (.A1(\wfg_core_top.cfg_subcycle_q[9] ),
    .A2(_02643_),
    .B1(_02636_),
    .X(_02653_));
 sky130_fd_sc_hd__o211a_1 _20065_ (.A1(\wfg_core_top.wbs_dat_o[9] ),
    .A2(_02642_),
    .B1(_02653_),
    .C1(_02647_),
    .X(_01263_));
 sky130_fd_sc_hd__buf_2 _20066_ (.A(_02635_),
    .X(_02654_));
 sky130_fd_sc_hd__a21o_1 _20067_ (.A1(\wfg_core_top.cfg_subcycle_q[10] ),
    .A2(_02643_),
    .B1(_02654_),
    .X(_02655_));
 sky130_fd_sc_hd__o211a_1 _20068_ (.A1(\wfg_core_top.wbs_dat_o[10] ),
    .A2(_02642_),
    .B1(_02655_),
    .C1(_02647_),
    .X(_01264_));
 sky130_fd_sc_hd__buf_2 _20069_ (.A(_02639_),
    .X(_02656_));
 sky130_fd_sc_hd__buf_2 _20070_ (.A(_02637_),
    .X(_02657_));
 sky130_fd_sc_hd__a21o_1 _20071_ (.A1(\wfg_core_top.cfg_subcycle_q[11] ),
    .A2(_02657_),
    .B1(_02654_),
    .X(_02658_));
 sky130_fd_sc_hd__o211a_1 _20072_ (.A1(\wfg_core_top.wbs_dat_o[11] ),
    .A2(_02656_),
    .B1(_02658_),
    .C1(_02647_),
    .X(_01265_));
 sky130_fd_sc_hd__a21o_1 _20073_ (.A1(\wfg_core_top.cfg_subcycle_q[12] ),
    .A2(_02657_),
    .B1(_02654_),
    .X(_02659_));
 sky130_fd_sc_hd__o211a_1 _20074_ (.A1(\wfg_core_top.wbs_dat_o[12] ),
    .A2(_02656_),
    .B1(_02659_),
    .C1(_02647_),
    .X(_01266_));
 sky130_fd_sc_hd__a21o_1 _20075_ (.A1(\wfg_core_top.cfg_subcycle_q[13] ),
    .A2(_02657_),
    .B1(_02654_),
    .X(_02660_));
 sky130_fd_sc_hd__buf_2 _20076_ (.A(_01589_),
    .X(_02661_));
 sky130_fd_sc_hd__o211a_1 _20077_ (.A1(\wfg_core_top.wbs_dat_o[13] ),
    .A2(_02656_),
    .B1(_02660_),
    .C1(_02661_),
    .X(_01267_));
 sky130_fd_sc_hd__a21o_1 _20078_ (.A1(\wfg_core_top.cfg_subcycle_q[14] ),
    .A2(_02657_),
    .B1(_02654_),
    .X(_02662_));
 sky130_fd_sc_hd__o211a_1 _20079_ (.A1(\wfg_core_top.wbs_dat_o[14] ),
    .A2(_02656_),
    .B1(_02662_),
    .C1(_02661_),
    .X(_01268_));
 sky130_fd_sc_hd__a21o_1 _20080_ (.A1(\wfg_core_top.cfg_subcycle_q[15] ),
    .A2(_02657_),
    .B1(_02654_),
    .X(_02663_));
 sky130_fd_sc_hd__o211a_1 _20081_ (.A1(\wfg_core_top.wbs_dat_o[15] ),
    .A2(_02656_),
    .B1(_02663_),
    .C1(_02661_),
    .X(_01269_));
 sky130_fd_sc_hd__a21o_1 _20082_ (.A1(\wfg_core_top.cfg_subcycle_q[16] ),
    .A2(_02657_),
    .B1(_02654_),
    .X(_02664_));
 sky130_fd_sc_hd__o211a_1 _20083_ (.A1(\wfg_core_top.wbs_dat_o[16] ),
    .A2(_02656_),
    .B1(_02664_),
    .C1(_02661_),
    .X(_01270_));
 sky130_fd_sc_hd__a21o_1 _20084_ (.A1(\wfg_core_top.cfg_subcycle_q[17] ),
    .A2(_02657_),
    .B1(_02654_),
    .X(_02665_));
 sky130_fd_sc_hd__o211a_1 _20085_ (.A1(\wfg_core_top.wbs_dat_o[17] ),
    .A2(_02656_),
    .B1(_02665_),
    .C1(_02661_),
    .X(_01271_));
 sky130_fd_sc_hd__a21o_1 _20086_ (.A1(\wfg_core_top.cfg_subcycle_q[18] ),
    .A2(_02657_),
    .B1(_02654_),
    .X(_02666_));
 sky130_fd_sc_hd__o211a_1 _20087_ (.A1(\wfg_core_top.wbs_dat_o[18] ),
    .A2(_02656_),
    .B1(_02666_),
    .C1(_02661_),
    .X(_01272_));
 sky130_fd_sc_hd__a21o_1 _20088_ (.A1(\wfg_core_top.cfg_subcycle_q[19] ),
    .A2(_02657_),
    .B1(_02654_),
    .X(_02667_));
 sky130_fd_sc_hd__o211a_1 _20089_ (.A1(\wfg_core_top.wbs_dat_o[19] ),
    .A2(_02656_),
    .B1(_02667_),
    .C1(_02661_),
    .X(_01273_));
 sky130_fd_sc_hd__a21o_1 _20090_ (.A1(\wfg_core_top.cfg_subcycle_q[20] ),
    .A2(_02657_),
    .B1(_02635_),
    .X(_02668_));
 sky130_fd_sc_hd__o211a_1 _20091_ (.A1(\wfg_core_top.wbs_dat_o[20] ),
    .A2(_02656_),
    .B1(_02668_),
    .C1(_02661_),
    .X(_01274_));
 sky130_fd_sc_hd__a21o_1 _20092_ (.A1(\wfg_core_top.cfg_subcycle_q[21] ),
    .A2(_02637_),
    .B1(_02635_),
    .X(_02669_));
 sky130_fd_sc_hd__o211a_1 _20093_ (.A1(\wfg_core_top.wbs_dat_o[21] ),
    .A2(_02639_),
    .B1(_02669_),
    .C1(_02661_),
    .X(_01275_));
 sky130_fd_sc_hd__a21o_1 _20094_ (.A1(\wfg_core_top.cfg_subcycle_q[22] ),
    .A2(_02637_),
    .B1(_02635_),
    .X(_02670_));
 sky130_fd_sc_hd__o211a_1 _20095_ (.A1(\wfg_core_top.wbs_dat_o[22] ),
    .A2(_02639_),
    .B1(_02670_),
    .C1(_02661_),
    .X(_01276_));
 sky130_fd_sc_hd__a21o_1 _20096_ (.A1(\wfg_core_top.cfg_subcycle_q[23] ),
    .A2(_02637_),
    .B1(_02635_),
    .X(_02671_));
 sky130_fd_sc_hd__buf_4 _20097_ (.A(_01589_),
    .X(_02672_));
 sky130_fd_sc_hd__o211a_1 _20098_ (.A1(\wfg_core_top.wbs_dat_o[23] ),
    .A2(_02639_),
    .B1(_02671_),
    .C1(_02672_),
    .X(_01277_));
 sky130_fd_sc_hd__nand2_1 _20099_ (.A(_02203_),
    .B(_02239_),
    .Y(_02673_));
 sky130_fd_sc_hd__a31o_1 _20100_ (.A1(_02203_),
    .A2(_01709_),
    .A3(_02239_),
    .B1(\wfg_drive_spi_top.ctrl_en_q ),
    .X(_02674_));
 sky130_fd_sc_hd__o311a_1 _20101_ (.A1(_01660_),
    .A2(_01691_),
    .A3(_02673_),
    .B1(_02674_),
    .C1(_01600_),
    .X(_01278_));
 sky130_fd_sc_hd__or4_2 _20102_ (.A(_01431_),
    .B(_01425_),
    .C(_01605_),
    .D(_01686_),
    .X(_02675_));
 sky130_fd_sc_hd__or2_1 _20103_ (.A(_01959_),
    .B(_02675_),
    .X(_02676_));
 sky130_fd_sc_hd__clkbuf_2 _20104_ (.A(_02676_),
    .X(_02677_));
 sky130_fd_sc_hd__nor2_1 _20105_ (.A(_01959_),
    .B(_02673_),
    .Y(_02678_));
 sky130_fd_sc_hd__or2_1 _20106_ (.A(\wfg_drive_spi_top.cfg_core_sel_q ),
    .B(_02678_),
    .X(_02679_));
 sky130_fd_sc_hd__o211a_1 _20107_ (.A1(_01675_),
    .A2(_02677_),
    .B1(_02679_),
    .C1(_02672_),
    .X(_01279_));
 sky130_fd_sc_hd__or2_1 _20108_ (.A(\wfg_drive_spi_top.cfg_cpol_q ),
    .B(_02678_),
    .X(_02680_));
 sky130_fd_sc_hd__o211a_1 _20109_ (.A1(_01660_),
    .A2(_02677_),
    .B1(_02680_),
    .C1(_02672_),
    .X(_01280_));
 sky130_fd_sc_hd__or2_1 _20110_ (.A(\wfg_drive_spi_top.cfg_dff_q[2] ),
    .B(_02678_),
    .X(_02681_));
 sky130_fd_sc_hd__o211a_1 _20111_ (.A1(_01666_),
    .A2(_02677_),
    .B1(_02681_),
    .C1(_02672_),
    .X(_01281_));
 sky130_fd_sc_hd__or2_1 _20112_ (.A(\wfg_drive_spi_top.cfg_dff_q[3] ),
    .B(_02678_),
    .X(_02682_));
 sky130_fd_sc_hd__o211a_1 _20113_ (.A1(_01669_),
    .A2(_02677_),
    .B1(_02682_),
    .C1(_02672_),
    .X(_01282_));
 sky130_fd_sc_hd__or2_1 _20114_ (.A(\wfg_drive_spi_top.cfg_lsbfirst_q ),
    .B(_02678_),
    .X(_02683_));
 sky130_fd_sc_hd__o211a_1 _20115_ (.A1(_01663_),
    .A2(_02677_),
    .B1(_02683_),
    .C1(_02672_),
    .X(_01283_));
 sky130_fd_sc_hd__or2_1 _20116_ (.A(\wfg_drive_spi_top.cfg_sspol_q ),
    .B(_02678_),
    .X(_02684_));
 sky130_fd_sc_hd__o211a_1 _20117_ (.A1(_01672_),
    .A2(_02677_),
    .B1(_02684_),
    .C1(_02672_),
    .X(_01284_));
 sky130_fd_sc_hd__or2_1 _20118_ (.A(_01763_),
    .B(_02675_),
    .X(_02685_));
 sky130_fd_sc_hd__buf_2 _20119_ (.A(_02685_),
    .X(_02686_));
 sky130_fd_sc_hd__nor2_2 _20120_ (.A(_01763_),
    .B(_02673_),
    .Y(_02687_));
 sky130_fd_sc_hd__or2_1 _20121_ (.A(\wfg_drive_spi_top.clkcfg_div_q[0] ),
    .B(_02687_),
    .X(_02688_));
 sky130_fd_sc_hd__o211a_1 _20122_ (.A1(_01660_),
    .A2(_02686_),
    .B1(_02688_),
    .C1(_02672_),
    .X(_01285_));
 sky130_fd_sc_hd__or2_1 _20123_ (.A(\wfg_drive_spi_top.clkcfg_div_q[1] ),
    .B(_02687_),
    .X(_02689_));
 sky130_fd_sc_hd__o211a_1 _20124_ (.A1(_01663_),
    .A2(_02686_),
    .B1(_02689_),
    .C1(_02672_),
    .X(_01286_));
 sky130_fd_sc_hd__or2_1 _20125_ (.A(\wfg_drive_spi_top.clkcfg_div_q[2] ),
    .B(_02687_),
    .X(_02690_));
 sky130_fd_sc_hd__o211a_1 _20126_ (.A1(_01666_),
    .A2(_02686_),
    .B1(_02690_),
    .C1(_02672_),
    .X(_01287_));
 sky130_fd_sc_hd__or2_1 _20127_ (.A(\wfg_drive_spi_top.clkcfg_div_q[3] ),
    .B(_02687_),
    .X(_02691_));
 sky130_fd_sc_hd__o211a_1 _20128_ (.A1(_01669_),
    .A2(_02686_),
    .B1(_02691_),
    .C1(_01600_),
    .X(_01288_));
 sky130_fd_sc_hd__or2_1 _20129_ (.A(\wfg_drive_spi_top.clkcfg_div_q[4] ),
    .B(_02687_),
    .X(_02692_));
 sky130_fd_sc_hd__o211a_1 _20130_ (.A1(_01672_),
    .A2(_02686_),
    .B1(_02692_),
    .C1(_01600_),
    .X(_01289_));
 sky130_fd_sc_hd__or2_1 _20131_ (.A(\wfg_drive_spi_top.clkcfg_div_q[5] ),
    .B(_02687_),
    .X(_02693_));
 sky130_fd_sc_hd__o211a_1 _20132_ (.A1(_01675_),
    .A2(_02686_),
    .B1(_02693_),
    .C1(_01600_),
    .X(_01290_));
 sky130_fd_sc_hd__or2_1 _20133_ (.A(\wfg_drive_spi_top.clkcfg_div_q[6] ),
    .B(_02687_),
    .X(_02694_));
 sky130_fd_sc_hd__o211a_1 _20134_ (.A1(_01679_),
    .A2(_02686_),
    .B1(_02694_),
    .C1(_01600_),
    .X(_01291_));
 sky130_fd_sc_hd__or2_1 _20135_ (.A(\wfg_drive_spi_top.clkcfg_div_q[7] ),
    .B(_02687_),
    .X(_02695_));
 sky130_fd_sc_hd__o211a_1 _20136_ (.A1(_01682_),
    .A2(_02686_),
    .B1(_02695_),
    .C1(_01600_),
    .X(_01292_));
 sky130_fd_sc_hd__dfrtp_1 _20137_ (.CLK(clknet_leaf_99_io_wbs_clk),
    .D(_00004_),
    .RESET_B(_00040_),
    .Q(\wfg_core_top.wfg_core.subcycle_count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _20138_ (.CLK(clknet_leaf_99_io_wbs_clk),
    .D(_00011_),
    .RESET_B(_00041_),
    .Q(\wfg_core_top.wfg_core.subcycle_count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _20139_ (.CLK(clknet_leaf_99_io_wbs_clk),
    .D(_00012_),
    .RESET_B(_00042_),
    .Q(\wfg_core_top.wfg_core.subcycle_count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _20140_ (.CLK(clknet_leaf_99_io_wbs_clk),
    .D(_00013_),
    .RESET_B(_00043_),
    .Q(\wfg_core_top.wfg_core.subcycle_count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _20141_ (.CLK(clknet_leaf_99_io_wbs_clk),
    .D(_00014_),
    .RESET_B(_00044_),
    .Q(\wfg_core_top.wfg_core.subcycle_count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _20142_ (.CLK(clknet_leaf_104_io_wbs_clk),
    .D(_00015_),
    .RESET_B(_00045_),
    .Q(\wfg_core_top.wfg_core.subcycle_count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _20143_ (.CLK(clknet_leaf_99_io_wbs_clk),
    .D(_00016_),
    .RESET_B(_00046_),
    .Q(\wfg_core_top.wfg_core.subcycle_count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _20144_ (.CLK(clknet_leaf_99_io_wbs_clk),
    .D(_00017_),
    .RESET_B(_00047_),
    .Q(\wfg_core_top.wfg_core.subcycle_count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _20145_ (.CLK(clknet_leaf_98_io_wbs_clk),
    .D(_00018_),
    .RESET_B(_00048_),
    .Q(\wfg_core_top.wfg_core.subcycle_count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _20146_ (.CLK(clknet_leaf_98_io_wbs_clk),
    .D(_00019_),
    .RESET_B(_00049_),
    .Q(\wfg_core_top.wfg_core.subcycle_count[9] ));
 sky130_fd_sc_hd__dfrtp_1 _20147_ (.CLK(clknet_leaf_79_io_wbs_clk),
    .D(_00005_),
    .RESET_B(_00050_),
    .Q(\wfg_core_top.wfg_core.subcycle_count[10] ));
 sky130_fd_sc_hd__dfrtp_1 _20148_ (.CLK(clknet_leaf_79_io_wbs_clk),
    .D(_00006_),
    .RESET_B(_00051_),
    .Q(\wfg_core_top.wfg_core.subcycle_count[11] ));
 sky130_fd_sc_hd__dfrtp_1 _20149_ (.CLK(clknet_leaf_78_io_wbs_clk),
    .D(_00007_),
    .RESET_B(_00052_),
    .Q(\wfg_core_top.wfg_core.subcycle_count[12] ));
 sky130_fd_sc_hd__dfrtp_1 _20150_ (.CLK(clknet_leaf_78_io_wbs_clk),
    .D(_00008_),
    .RESET_B(_00053_),
    .Q(\wfg_core_top.wfg_core.subcycle_count[13] ));
 sky130_fd_sc_hd__dfrtp_1 _20151_ (.CLK(clknet_leaf_78_io_wbs_clk),
    .D(_00009_),
    .RESET_B(_00054_),
    .Q(\wfg_core_top.wfg_core.subcycle_count[14] ));
 sky130_fd_sc_hd__dfrtp_1 _20152_ (.CLK(clknet_leaf_78_io_wbs_clk),
    .D(_00010_),
    .RESET_B(_00055_),
    .Q(\wfg_core_top.wfg_core.subcycle_count[15] ));
 sky130_fd_sc_hd__dfrtp_1 _20153_ (.CLK(clknet_leaf_96_io_wbs_clk),
    .D(_00472_),
    .RESET_B(_00056_),
    .Q(\wfg_core_top.wfg_core.sync_count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _20154_ (.CLK(clknet_leaf_96_io_wbs_clk),
    .D(_00473_),
    .RESET_B(_00057_),
    .Q(\wfg_core_top.wfg_core.sync_count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _20155_ (.CLK(clknet_leaf_97_io_wbs_clk),
    .D(_00474_),
    .RESET_B(_00058_),
    .Q(\wfg_core_top.wfg_core.sync_count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _20156_ (.CLK(clknet_leaf_97_io_wbs_clk),
    .D(_00475_),
    .RESET_B(_00059_),
    .Q(\wfg_core_top.wfg_core.sync_count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _20157_ (.CLK(clknet_leaf_97_io_wbs_clk),
    .D(_00476_),
    .RESET_B(_00060_),
    .Q(\wfg_core_top.wfg_core.sync_count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _20158_ (.CLK(clknet_leaf_97_io_wbs_clk),
    .D(_00477_),
    .RESET_B(_00061_),
    .Q(\wfg_core_top.wfg_core.sync_count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _20159_ (.CLK(clknet_leaf_97_io_wbs_clk),
    .D(_00478_),
    .RESET_B(_00062_),
    .Q(\wfg_core_top.wfg_core.sync_count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _20160_ (.CLK(clknet_leaf_97_io_wbs_clk),
    .D(_00479_),
    .RESET_B(_00063_),
    .Q(\wfg_core_top.wfg_core.sync_count[7] ));
 sky130_fd_sc_hd__dfrtp_2 _20161_ (.CLK(clknet_leaf_98_io_wbs_clk),
    .D(_00480_),
    .RESET_B(_00064_),
    .Q(\wfg_core_top.wfg_core.temp_subcycle ));
 sky130_fd_sc_hd__dfrtp_2 _20162_ (.CLK(clknet_leaf_97_io_wbs_clk),
    .D(_00481_),
    .RESET_B(_00065_),
    .Q(\wfg_core_top.wfg_core.temp_sync ));
 sky130_fd_sc_hd__dfxtp_1 _20163_ (.CLK(clknet_leaf_15_io_wbs_clk),
    .D(_00482_),
    .Q(\wfg_core_top.wfg_core.subcycle_dly ));
 sky130_fd_sc_hd__dfxtp_1 _20164_ (.CLK(clknet_leaf_16_io_wbs_clk),
    .D(_00483_),
    .Q(\wfg_core_top.wfg_core.sync_dly ));
 sky130_fd_sc_hd__dfrtp_2 _20165_ (.CLK(clknet_leaf_16_io_wbs_clk),
    .D(_00484_),
    .RESET_B(_00066_),
    .Q(\wfg_core_top.wfg_core.subcycle_pls_cnt[0] ));
 sky130_fd_sc_hd__dfrtp_2 _20166_ (.CLK(clknet_leaf_16_io_wbs_clk),
    .D(_00485_),
    .RESET_B(_00067_),
    .Q(\wfg_core_top.wfg_core.subcycle_pls_cnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _20167_ (.CLK(clknet_leaf_16_io_wbs_clk),
    .D(_00486_),
    .RESET_B(_00068_),
    .Q(\wfg_core_top.wfg_core.subcycle_pls_cnt[2] ));
 sky130_fd_sc_hd__dfrtp_1 _20168_ (.CLK(clknet_leaf_16_io_wbs_clk),
    .D(_00487_),
    .RESET_B(_00069_),
    .Q(\wfg_core_top.wfg_core.subcycle_pls_cnt[3] ));
 sky130_fd_sc_hd__dfrtp_1 _20169_ (.CLK(clknet_leaf_16_io_wbs_clk),
    .D(_00488_),
    .RESET_B(_00070_),
    .Q(\wfg_core_top.wfg_core.subcycle_pls_cnt[4] ));
 sky130_fd_sc_hd__dfrtp_1 _20170_ (.CLK(clknet_leaf_17_io_wbs_clk),
    .D(_00489_),
    .RESET_B(_00071_),
    .Q(\wfg_core_top.wfg_core.subcycle_pls_cnt[5] ));
 sky130_fd_sc_hd__dfrtp_1 _20171_ (.CLK(clknet_leaf_40_io_wbs_clk),
    .D(_00490_),
    .RESET_B(_00072_),
    .Q(\wfg_core_top.wfg_core.subcycle_pls_cnt[6] ));
 sky130_fd_sc_hd__dfrtp_1 _20172_ (.CLK(clknet_leaf_40_io_wbs_clk),
    .D(_00491_),
    .RESET_B(_00073_),
    .Q(\wfg_core_top.wfg_core.subcycle_pls_cnt[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20173_ (.CLK(clknet_leaf_99_io_wbs_clk),
    .D(_00492_),
    .Q(\wfg_core_top.cfg_subcycle_q[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20174_ (.CLK(clknet_leaf_100_io_wbs_clk),
    .D(_00493_),
    .Q(\wfg_core_top.cfg_subcycle_q[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20175_ (.CLK(clknet_leaf_99_io_wbs_clk),
    .D(_00494_),
    .Q(\wfg_core_top.cfg_subcycle_q[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20176_ (.CLK(clknet_leaf_98_io_wbs_clk),
    .D(_00495_),
    .Q(\wfg_core_top.cfg_subcycle_q[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20177_ (.CLK(clknet_leaf_100_io_wbs_clk),
    .D(_00496_),
    .Q(\wfg_core_top.cfg_subcycle_q[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20178_ (.CLK(clknet_leaf_99_io_wbs_clk),
    .D(_00497_),
    .Q(\wfg_core_top.cfg_subcycle_q[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20179_ (.CLK(clknet_leaf_99_io_wbs_clk),
    .D(_00498_),
    .Q(\wfg_core_top.cfg_subcycle_q[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20180_ (.CLK(clknet_leaf_98_io_wbs_clk),
    .D(_00499_),
    .Q(\wfg_core_top.cfg_subcycle_q[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20181_ (.CLK(clknet_leaf_98_io_wbs_clk),
    .D(_00500_),
    .Q(\wfg_core_top.cfg_subcycle_q[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20182_ (.CLK(clknet_leaf_98_io_wbs_clk),
    .D(_00501_),
    .Q(\wfg_core_top.cfg_subcycle_q[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20183_ (.CLK(clknet_leaf_79_io_wbs_clk),
    .D(_00502_),
    .Q(\wfg_core_top.cfg_subcycle_q[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20184_ (.CLK(clknet_leaf_79_io_wbs_clk),
    .D(_00503_),
    .Q(\wfg_core_top.cfg_subcycle_q[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20185_ (.CLK(clknet_leaf_78_io_wbs_clk),
    .D(_00504_),
    .Q(\wfg_core_top.cfg_subcycle_q[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20186_ (.CLK(clknet_leaf_79_io_wbs_clk),
    .D(_00505_),
    .Q(\wfg_core_top.cfg_subcycle_q[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20187_ (.CLK(clknet_leaf_80_io_wbs_clk),
    .D(_00506_),
    .Q(\wfg_core_top.cfg_subcycle_q[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20188_ (.CLK(clknet_leaf_79_io_wbs_clk),
    .D(_00507_),
    .Q(\wfg_core_top.cfg_subcycle_q[23] ));
 sky130_fd_sc_hd__dfxtp_1 _20189_ (.CLK(clknet_leaf_95_io_wbs_clk),
    .D(_00508_),
    .Q(\wfg_core_top.cfg_sync_q[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20190_ (.CLK(clknet_leaf_79_io_wbs_clk),
    .D(_00509_),
    .Q(\wfg_core_top.cfg_sync_q[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20191_ (.CLK(clknet_leaf_96_io_wbs_clk),
    .D(_00510_),
    .Q(\wfg_core_top.cfg_sync_q[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20192_ (.CLK(clknet_leaf_96_io_wbs_clk),
    .D(_00511_),
    .Q(\wfg_core_top.cfg_sync_q[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20193_ (.CLK(clknet_leaf_98_io_wbs_clk),
    .D(_00512_),
    .Q(\wfg_core_top.cfg_sync_q[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20194_ (.CLK(clknet_leaf_95_io_wbs_clk),
    .D(_00513_),
    .Q(\wfg_core_top.cfg_sync_q[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20195_ (.CLK(clknet_leaf_95_io_wbs_clk),
    .D(_00514_),
    .Q(\wfg_core_top.cfg_sync_q[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20196_ (.CLK(clknet_leaf_95_io_wbs_clk),
    .D(_00515_),
    .Q(\wfg_core_top.cfg_sync_q[7] ));
 sky130_fd_sc_hd__dfxtp_4 _20197_ (.CLK(clknet_leaf_101_io_wbs_clk),
    .D(_00516_),
    .Q(\wfg_core_top.active_o ));
 sky130_fd_sc_hd__dfxtp_1 _20198_ (.CLK(clknet_leaf_91_io_wbs_clk),
    .D(_00517_),
    .Q(\wfg_subcore_top.wbs_ack_o ));
 sky130_fd_sc_hd__dfstp_1 _20199_ (.CLK(clknet_leaf_23_io_wbs_clk),
    .D(_00001_),
    .SET_B(_00074_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.cur_state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _20200_ (.CLK(clknet_leaf_22_io_wbs_clk),
    .D(\wfg_stim_mem_top.wfg_stim_mem.cur_state[2] ),
    .RESET_B(_00075_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.cur_state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _20201_ (.CLK(clknet_leaf_22_io_wbs_clk),
    .D(_00000_),
    .RESET_B(_00076_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.cur_state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _20202_ (.CLK(clknet_leaf_22_io_wbs_clk),
    .D(_00002_),
    .RESET_B(_00077_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.cur_state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20203_ (.CLK(clknet_leaf_101_io_wbs_clk),
    .D(_00518_),
    .Q(\wfg_core_top.wbs_ack_o ));
 sky130_fd_sc_hd__dfrtp_1 _20204_ (.CLK(clknet_leaf_17_io_wbs_clk),
    .D(\wfg_drive_pat_top.wfg_drive_pat.wfg_sync_i ),
    .RESET_B(_00078_),
    .Q(\wfg_drive_pat_top.wfg_axis_tready_o ));
 sky130_fd_sc_hd__dfrtp_1 _20205_ (.CLK(clknet_leaf_31_io_wbs_clk),
    .D(_00519_),
    .RESET_B(_00079_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[0].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_1 _20206_ (.CLK(clknet_leaf_48_io_wbs_clk),
    .D(_00520_),
    .RESET_B(_00080_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[1].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_1 _20207_ (.CLK(clknet_leaf_46_io_wbs_clk),
    .D(_00521_),
    .RESET_B(_00081_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[2].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_4 _20208_ (.CLK(clknet_leaf_47_io_wbs_clk),
    .D(_00522_),
    .RESET_B(_00082_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[3].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_2 _20209_ (.CLK(clknet_leaf_47_io_wbs_clk),
    .D(_00523_),
    .RESET_B(_00083_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[4].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_4 _20210_ (.CLK(clknet_leaf_45_io_wbs_clk),
    .D(_00524_),
    .RESET_B(_00084_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[5].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_4 _20211_ (.CLK(clknet_leaf_47_io_wbs_clk),
    .D(_00525_),
    .RESET_B(_00085_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[6].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_4 _20212_ (.CLK(clknet_leaf_45_io_wbs_clk),
    .D(_00526_),
    .RESET_B(_00086_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[7].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_4 _20213_ (.CLK(clknet_leaf_45_io_wbs_clk),
    .D(_00527_),
    .RESET_B(_00087_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[8].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_1 _20214_ (.CLK(clknet_leaf_45_io_wbs_clk),
    .D(_00528_),
    .RESET_B(_00088_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[9].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_2 _20215_ (.CLK(clknet_leaf_52_io_wbs_clk),
    .D(_00529_),
    .RESET_B(_00089_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[10].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_4 _20216_ (.CLK(clknet_leaf_52_io_wbs_clk),
    .D(_00530_),
    .RESET_B(_00090_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[11].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_4 _20217_ (.CLK(clknet_leaf_62_io_wbs_clk),
    .D(_00531_),
    .RESET_B(_00091_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[12].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_2 _20218_ (.CLK(clknet_leaf_52_io_wbs_clk),
    .D(_00532_),
    .RESET_B(_00092_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[13].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_2 _20219_ (.CLK(clknet_leaf_52_io_wbs_clk),
    .D(_00533_),
    .RESET_B(_00093_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[14].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_2 _20220_ (.CLK(clknet_leaf_62_io_wbs_clk),
    .D(_00534_),
    .RESET_B(_00094_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[15].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_2 _20221_ (.CLK(clknet_leaf_62_io_wbs_clk),
    .D(_00535_),
    .RESET_B(_00095_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[16].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_2 _20222_ (.CLK(clknet_leaf_61_io_wbs_clk),
    .D(_00536_),
    .RESET_B(_00096_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[17].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_1 _20223_ (.CLK(clknet_leaf_62_io_wbs_clk),
    .D(_00537_),
    .RESET_B(_00097_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[18].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_2 _20224_ (.CLK(clknet_leaf_61_io_wbs_clk),
    .D(_00538_),
    .RESET_B(_00098_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[19].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_1 _20225_ (.CLK(clknet_leaf_61_io_wbs_clk),
    .D(_00539_),
    .RESET_B(_00099_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[20].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_1 _20226_ (.CLK(clknet_leaf_62_io_wbs_clk),
    .D(_00540_),
    .RESET_B(_00100_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[21].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_2 _20227_ (.CLK(clknet_leaf_61_io_wbs_clk),
    .D(_00541_),
    .RESET_B(_00101_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[22].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_1 _20228_ (.CLK(clknet_leaf_59_io_wbs_clk),
    .D(_00542_),
    .RESET_B(_00102_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[23].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_1 _20229_ (.CLK(clknet_leaf_60_io_wbs_clk),
    .D(_00543_),
    .RESET_B(_00103_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[24].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_1 _20230_ (.CLK(clknet_leaf_60_io_wbs_clk),
    .D(_00544_),
    .RESET_B(_00104_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[25].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_1 _20231_ (.CLK(clknet_leaf_59_io_wbs_clk),
    .D(_00545_),
    .RESET_B(_00105_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[26].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_1 _20232_ (.CLK(clknet_leaf_59_io_wbs_clk),
    .D(_00546_),
    .RESET_B(_00106_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[27].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_1 _20233_ (.CLK(clknet_leaf_59_io_wbs_clk),
    .D(_00547_),
    .RESET_B(_00107_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[28].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_2 _20234_ (.CLK(clknet_leaf_61_io_wbs_clk),
    .D(_00548_),
    .RESET_B(_00108_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[29].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_1 _20235_ (.CLK(clknet_leaf_61_io_wbs_clk),
    .D(_00549_),
    .RESET_B(_00109_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[30].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_1 _20236_ (.CLK(clknet_leaf_61_io_wbs_clk),
    .D(_00550_),
    .RESET_B(_00110_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[31].drv.axis_data_ff ));
 sky130_fd_sc_hd__dfrtp_4 _20237_ (.CLK(clknet_leaf_45_io_wbs_clk),
    .D(_00551_),
    .RESET_B(_00111_),
    .Q(net155));
 sky130_fd_sc_hd__dfrtp_4 _20238_ (.CLK(clknet_leaf_62_io_wbs_clk),
    .D(_00552_),
    .RESET_B(_00112_),
    .Q(net166));
 sky130_fd_sc_hd__dfrtp_2 _20239_ (.CLK(clknet_leaf_62_io_wbs_clk),
    .D(_00553_),
    .RESET_B(_00113_),
    .Q(net169));
 sky130_fd_sc_hd__dfrtp_4 _20240_ (.CLK(clknet_leaf_34_io_wbs_clk),
    .D(_00554_),
    .RESET_B(_00114_),
    .Q(net170));
 sky130_fd_sc_hd__dfrtp_4 _20241_ (.CLK(clknet_leaf_34_io_wbs_clk),
    .D(_00555_),
    .RESET_B(_00115_),
    .Q(net171));
 sky130_fd_sc_hd__dfrtp_4 _20242_ (.CLK(clknet_leaf_33_io_wbs_clk),
    .D(_00556_),
    .RESET_B(_00116_),
    .Q(net172));
 sky130_fd_sc_hd__dfrtp_4 _20243_ (.CLK(clknet_leaf_34_io_wbs_clk),
    .D(_00557_),
    .RESET_B(_00117_),
    .Q(net173));
 sky130_fd_sc_hd__dfrtp_4 _20244_ (.CLK(clknet_leaf_33_io_wbs_clk),
    .D(_00558_),
    .RESET_B(_00118_),
    .Q(net174));
 sky130_fd_sc_hd__dfrtp_4 _20245_ (.CLK(clknet_leaf_33_io_wbs_clk),
    .D(_00559_),
    .RESET_B(_00119_),
    .Q(net175));
 sky130_fd_sc_hd__dfrtp_4 _20246_ (.CLK(clknet_leaf_32_io_wbs_clk),
    .D(_00560_),
    .RESET_B(_00120_),
    .Q(net145));
 sky130_fd_sc_hd__dfrtp_4 _20247_ (.CLK(clknet_leaf_31_io_wbs_clk),
    .D(_00561_),
    .RESET_B(_00121_),
    .Q(net146));
 sky130_fd_sc_hd__dfrtp_4 _20248_ (.CLK(clknet_leaf_32_io_wbs_clk),
    .D(_00562_),
    .RESET_B(_00122_),
    .Q(net147));
 sky130_fd_sc_hd__dfrtp_4 _20249_ (.CLK(clknet_leaf_31_io_wbs_clk),
    .D(_00563_),
    .RESET_B(_00123_),
    .Q(net148));
 sky130_fd_sc_hd__dfrtp_4 _20250_ (.CLK(clknet_leaf_47_io_wbs_clk),
    .D(_00564_),
    .RESET_B(_00124_),
    .Q(net149));
 sky130_fd_sc_hd__dfxtp_1 _20251_ (.CLK(clknet_leaf_90_io_wbs_clk),
    .D(_00565_),
    .Q(\wfg_subcore_top.wbs_dat_o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20252_ (.CLK(clknet_leaf_91_io_wbs_clk),
    .D(_00566_),
    .Q(\wfg_subcore_top.wbs_dat_o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20253_ (.CLK(clknet_leaf_91_io_wbs_clk),
    .D(_00567_),
    .Q(\wfg_subcore_top.wbs_dat_o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20254_ (.CLK(clknet_leaf_91_io_wbs_clk),
    .D(_00568_),
    .Q(\wfg_subcore_top.wbs_dat_o[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20255_ (.CLK(clknet_leaf_11_io_wbs_clk),
    .D(_00569_),
    .Q(\wfg_subcore_top.wbs_dat_o[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20256_ (.CLK(clknet_leaf_102_io_wbs_clk),
    .D(_00570_),
    .Q(\wfg_subcore_top.wbs_dat_o[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20257_ (.CLK(clknet_leaf_11_io_wbs_clk),
    .D(_00571_),
    .Q(\wfg_subcore_top.wbs_dat_o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20258_ (.CLK(clknet_leaf_102_io_wbs_clk),
    .D(_00572_),
    .Q(\wfg_subcore_top.wbs_dat_o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20259_ (.CLK(clknet_leaf_11_io_wbs_clk),
    .D(_00573_),
    .Q(\wfg_subcore_top.wbs_dat_o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20260_ (.CLK(clknet_leaf_91_io_wbs_clk),
    .D(_00574_),
    .Q(\wfg_subcore_top.wbs_dat_o[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20261_ (.CLK(clknet_leaf_90_io_wbs_clk),
    .D(_00575_),
    .Q(\wfg_subcore_top.wbs_dat_o[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20262_ (.CLK(clknet_leaf_90_io_wbs_clk),
    .D(_00576_),
    .Q(\wfg_subcore_top.wbs_dat_o[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20263_ (.CLK(clknet_leaf_90_io_wbs_clk),
    .D(_00577_),
    .Q(\wfg_subcore_top.wbs_dat_o[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20264_ (.CLK(clknet_leaf_89_io_wbs_clk),
    .D(_00578_),
    .Q(\wfg_subcore_top.wbs_dat_o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20265_ (.CLK(clknet_leaf_88_io_wbs_clk),
    .D(_00579_),
    .Q(\wfg_subcore_top.wbs_dat_o[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20266_ (.CLK(clknet_leaf_90_io_wbs_clk),
    .D(_00580_),
    .Q(\wfg_subcore_top.wbs_dat_o[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20267_ (.CLK(clknet_leaf_89_io_wbs_clk),
    .D(_00581_),
    .Q(\wfg_subcore_top.wbs_dat_o[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20268_ (.CLK(clknet_leaf_90_io_wbs_clk),
    .D(_00582_),
    .Q(\wfg_subcore_top.wbs_dat_o[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20269_ (.CLK(clknet_leaf_89_io_wbs_clk),
    .D(_00583_),
    .Q(\wfg_subcore_top.wbs_dat_o[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20270_ (.CLK(clknet_leaf_89_io_wbs_clk),
    .D(_00584_),
    .Q(\wfg_subcore_top.wbs_dat_o[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20271_ (.CLK(clknet_leaf_88_io_wbs_clk),
    .D(_00585_),
    .Q(\wfg_subcore_top.wbs_dat_o[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20272_ (.CLK(clknet_leaf_84_io_wbs_clk),
    .D(_00586_),
    .Q(\wfg_subcore_top.wbs_dat_o[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20273_ (.CLK(clknet_leaf_84_io_wbs_clk),
    .D(_00587_),
    .Q(\wfg_subcore_top.wbs_dat_o[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20274_ (.CLK(clknet_leaf_84_io_wbs_clk),
    .D(_00588_),
    .Q(\wfg_subcore_top.wbs_dat_o[23] ));
 sky130_fd_sc_hd__dfrtp_4 _20275_ (.CLK(clknet_leaf_47_io_wbs_clk),
    .D(_00589_),
    .RESET_B(_00125_),
    .Q(net150));
 sky130_fd_sc_hd__dfrtp_4 _20276_ (.CLK(clknet_leaf_47_io_wbs_clk),
    .D(_00590_),
    .RESET_B(_00126_),
    .Q(net151));
 sky130_fd_sc_hd__dfrtp_4 _20277_ (.CLK(clknet_leaf_47_io_wbs_clk),
    .D(_00591_),
    .RESET_B(_00127_),
    .Q(net152));
 sky130_fd_sc_hd__dfrtp_4 _20278_ (.CLK(clknet_leaf_46_io_wbs_clk),
    .D(_00592_),
    .RESET_B(_00128_),
    .Q(net153));
 sky130_fd_sc_hd__dfrtp_4 _20279_ (.CLK(clknet_leaf_46_io_wbs_clk),
    .D(_00593_),
    .RESET_B(_00129_),
    .Q(net154));
 sky130_fd_sc_hd__dfrtp_4 _20280_ (.CLK(clknet_leaf_48_io_wbs_clk),
    .D(_00594_),
    .RESET_B(_00130_),
    .Q(net156));
 sky130_fd_sc_hd__dfrtp_4 _20281_ (.CLK(clknet_leaf_45_io_wbs_clk),
    .D(_00595_),
    .RESET_B(_00131_),
    .Q(net157));
 sky130_fd_sc_hd__dfrtp_4 _20282_ (.CLK(clknet_leaf_45_io_wbs_clk),
    .D(_00596_),
    .RESET_B(_00132_),
    .Q(net158));
 sky130_fd_sc_hd__dfrtp_4 _20283_ (.CLK(clknet_leaf_62_io_wbs_clk),
    .D(_00597_),
    .RESET_B(_00133_),
    .Q(net159));
 sky130_fd_sc_hd__dfrtp_4 _20284_ (.CLK(clknet_leaf_61_io_wbs_clk),
    .D(_00598_),
    .RESET_B(_00134_),
    .Q(net160));
 sky130_fd_sc_hd__dfrtp_4 _20285_ (.CLK(clknet_leaf_60_io_wbs_clk),
    .D(_00599_),
    .RESET_B(_00135_),
    .Q(net161));
 sky130_fd_sc_hd__dfrtp_4 _20286_ (.CLK(clknet_leaf_60_io_wbs_clk),
    .D(_00600_),
    .RESET_B(_00136_),
    .Q(net162));
 sky130_fd_sc_hd__dfrtp_4 _20287_ (.CLK(clknet_leaf_62_io_wbs_clk),
    .D(_00601_),
    .RESET_B(_00137_),
    .Q(net163));
 sky130_fd_sc_hd__dfrtp_4 _20288_ (.CLK(clknet_leaf_60_io_wbs_clk),
    .D(_00602_),
    .RESET_B(_00138_),
    .Q(net164));
 sky130_fd_sc_hd__dfrtp_4 _20289_ (.CLK(clknet_leaf_60_io_wbs_clk),
    .D(_00603_),
    .RESET_B(_00139_),
    .Q(net165));
 sky130_fd_sc_hd__dfrtp_4 _20290_ (.CLK(clknet_leaf_45_io_wbs_clk),
    .D(_00604_),
    .RESET_B(_00140_),
    .Q(net167));
 sky130_fd_sc_hd__dfrtp_2 _20291_ (.CLK(clknet_leaf_62_io_wbs_clk),
    .D(_00605_),
    .RESET_B(_00141_),
    .Q(net168));
 sky130_fd_sc_hd__dfrtp_4 _20292_ (.CLK(clknet_leaf_45_io_wbs_clk),
    .D(_00606_),
    .RESET_B(_00142_),
    .Q(net176));
 sky130_fd_sc_hd__dfxtp_1 _20293_ (.CLK(clknet_leaf_39_io_wbs_clk),
    .D(_00607_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20294_ (.CLK(clknet_leaf_17_io_wbs_clk),
    .D(_00608_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20295_ (.CLK(clknet_leaf_89_io_wbs_clk),
    .D(_00609_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20296_ (.CLK(clknet_leaf_18_io_wbs_clk),
    .D(_00610_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20297_ (.CLK(clknet_leaf_18_io_wbs_clk),
    .D(_00611_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20298_ (.CLK(clknet_leaf_90_io_wbs_clk),
    .D(_00612_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20299_ (.CLK(clknet_leaf_18_io_wbs_clk),
    .D(_00613_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20300_ (.CLK(clknet_leaf_18_io_wbs_clk),
    .D(_00614_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20301_ (.CLK(clknet_leaf_17_io_wbs_clk),
    .D(_00615_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20302_ (.CLK(clknet_leaf_17_io_wbs_clk),
    .D(_00616_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20303_ (.CLK(clknet_leaf_17_io_wbs_clk),
    .D(_00617_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20304_ (.CLK(clknet_leaf_16_io_wbs_clk),
    .D(_00618_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20305_ (.CLK(clknet_leaf_16_io_wbs_clk),
    .D(_00619_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20306_ (.CLK(clknet_leaf_41_io_wbs_clk),
    .D(_00620_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20307_ (.CLK(clknet_leaf_40_io_wbs_clk),
    .D(_00621_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20308_ (.CLK(clknet_leaf_89_io_wbs_clk),
    .D(_00622_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20309_ (.CLK(clknet_leaf_74_io_wbs_clk),
    .D(_00623_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20310_ (.CLK(clknet_leaf_41_io_wbs_clk),
    .D(_00624_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[17] ));
 sky130_fd_sc_hd__dfxtp_2 _20311_ (.CLK(clknet_leaf_71_io_wbs_clk),
    .D(_00625_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[18] ));
 sky130_fd_sc_hd__dfxtp_2 _20312_ (.CLK(clknet_leaf_71_io_wbs_clk),
    .D(_00626_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[19] ));
 sky130_fd_sc_hd__dfxtp_2 _20313_ (.CLK(clknet_leaf_70_io_wbs_clk),
    .D(_00627_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20314_ (.CLK(clknet_leaf_74_io_wbs_clk),
    .D(_00628_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[21] ));
 sky130_fd_sc_hd__dfxtp_2 _20315_ (.CLK(clknet_leaf_67_io_wbs_clk),
    .D(_00629_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20316_ (.CLK(clknet_leaf_40_io_wbs_clk),
    .D(_00630_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[23] ));
 sky130_fd_sc_hd__dfxtp_2 _20317_ (.CLK(clknet_leaf_66_io_wbs_clk),
    .D(_00631_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[24] ));
 sky130_fd_sc_hd__dfxtp_2 _20318_ (.CLK(clknet_leaf_64_io_wbs_clk),
    .D(_00632_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[25] ));
 sky130_fd_sc_hd__dfxtp_2 _20319_ (.CLK(clknet_leaf_68_io_wbs_clk),
    .D(_00633_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[26] ));
 sky130_fd_sc_hd__dfxtp_2 _20320_ (.CLK(clknet_leaf_66_io_wbs_clk),
    .D(_00634_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[27] ));
 sky130_fd_sc_hd__dfxtp_2 _20321_ (.CLK(clknet_leaf_66_io_wbs_clk),
    .D(_00635_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[28] ));
 sky130_fd_sc_hd__dfxtp_2 _20322_ (.CLK(clknet_leaf_68_io_wbs_clk),
    .D(_00636_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[29] ));
 sky130_fd_sc_hd__dfxtp_2 _20323_ (.CLK(clknet_leaf_67_io_wbs_clk),
    .D(_00637_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[30] ));
 sky130_fd_sc_hd__dfxtp_2 _20324_ (.CLK(clknet_leaf_67_io_wbs_clk),
    .D(_00638_),
    .Q(\wfg_drive_pat_top.wbs_dat_o[31] ));
 sky130_fd_sc_hd__dfxtp_1 _20325_ (.CLK(clknet_leaf_36_io_wbs_clk),
    .D(_00639_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[0].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20326_ (.CLK(clknet_leaf_42_io_wbs_clk),
    .D(_00640_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[1].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20327_ (.CLK(clknet_leaf_41_io_wbs_clk),
    .D(_00641_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[2].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20328_ (.CLK(clknet_leaf_21_io_wbs_clk),
    .D(_00642_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[3].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20329_ (.CLK(clknet_leaf_20_io_wbs_clk),
    .D(_00643_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[4].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20330_ (.CLK(clknet_leaf_21_io_wbs_clk),
    .D(_00644_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[5].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20331_ (.CLK(clknet_leaf_21_io_wbs_clk),
    .D(_00645_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[6].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20332_ (.CLK(clknet_leaf_21_io_wbs_clk),
    .D(_00646_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[7].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20333_ (.CLK(clknet_leaf_36_io_wbs_clk),
    .D(_00647_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[8].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20334_ (.CLK(clknet_leaf_43_io_wbs_clk),
    .D(_00648_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[9].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20335_ (.CLK(clknet_leaf_37_io_wbs_clk),
    .D(_00649_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[10].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20336_ (.CLK(clknet_leaf_36_io_wbs_clk),
    .D(_00650_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[11].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20337_ (.CLK(clknet_leaf_32_io_wbs_clk),
    .D(_00651_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[12].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20338_ (.CLK(clknet_leaf_43_io_wbs_clk),
    .D(_00652_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[13].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20339_ (.CLK(clknet_leaf_42_io_wbs_clk),
    .D(_00653_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[14].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20340_ (.CLK(clknet_leaf_43_io_wbs_clk),
    .D(_00654_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[15].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20341_ (.CLK(clknet_leaf_47_io_wbs_clk),
    .D(_00655_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[16].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20342_ (.CLK(clknet_leaf_44_io_wbs_clk),
    .D(_00656_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[17].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20343_ (.CLK(clknet_leaf_44_io_wbs_clk),
    .D(_00657_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[18].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20344_ (.CLK(clknet_leaf_70_io_wbs_clk),
    .D(_00658_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[19].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20345_ (.CLK(clknet_leaf_69_io_wbs_clk),
    .D(_00659_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[20].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20346_ (.CLK(clknet_leaf_69_io_wbs_clk),
    .D(_00660_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[21].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20347_ (.CLK(clknet_leaf_69_io_wbs_clk),
    .D(_00661_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[22].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20348_ (.CLK(clknet_leaf_64_io_wbs_clk),
    .D(_00662_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[23].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20349_ (.CLK(clknet_leaf_64_io_wbs_clk),
    .D(_00663_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[24].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20350_ (.CLK(clknet_leaf_65_io_wbs_clk),
    .D(_00664_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[25].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20351_ (.CLK(clknet_leaf_63_io_wbs_clk),
    .D(_00665_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[26].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20352_ (.CLK(clknet_leaf_65_io_wbs_clk),
    .D(_00666_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[27].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20353_ (.CLK(clknet_leaf_66_io_wbs_clk),
    .D(_00667_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[28].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20354_ (.CLK(clknet_leaf_64_io_wbs_clk),
    .D(_00668_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[29].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20355_ (.CLK(clknet_leaf_67_io_wbs_clk),
    .D(_00669_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[30].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20356_ (.CLK(clknet_leaf_67_io_wbs_clk),
    .D(_00670_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[31].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__dfxtp_1 _20357_ (.CLK(clknet_leaf_40_io_wbs_clk),
    .D(_00671_),
    .Q(\wfg_drive_pat_top.cfg_core_sel_q ));
 sky130_fd_sc_hd__dfxtp_1 _20358_ (.CLK(clknet_leaf_39_io_wbs_clk),
    .D(_00672_),
    .Q(\wfg_drive_pat_top.cfg_begin_q[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20359_ (.CLK(clknet_leaf_40_io_wbs_clk),
    .D(_00673_),
    .Q(\wfg_drive_pat_top.cfg_begin_q[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20360_ (.CLK(clknet_leaf_41_io_wbs_clk),
    .D(_00674_),
    .Q(\wfg_drive_pat_top.cfg_begin_q[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20361_ (.CLK(clknet_leaf_20_io_wbs_clk),
    .D(_00675_),
    .Q(\wfg_drive_pat_top.cfg_begin_q[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20362_ (.CLK(clknet_leaf_20_io_wbs_clk),
    .D(_00676_),
    .Q(\wfg_drive_pat_top.cfg_begin_q[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20363_ (.CLK(clknet_leaf_39_io_wbs_clk),
    .D(_00677_),
    .Q(\wfg_drive_pat_top.cfg_begin_q[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20364_ (.CLK(clknet_leaf_39_io_wbs_clk),
    .D(_00678_),
    .Q(\wfg_drive_pat_top.cfg_begin_q[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20365_ (.CLK(clknet_leaf_39_io_wbs_clk),
    .D(_00679_),
    .Q(\wfg_drive_pat_top.cfg_begin_q[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20366_ (.CLK(clknet_leaf_38_io_wbs_clk),
    .D(_00680_),
    .Q(\wfg_drive_pat_top.cfg_end_q[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20367_ (.CLK(clknet_leaf_41_io_wbs_clk),
    .D(_00681_),
    .Q(\wfg_drive_pat_top.cfg_end_q[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20368_ (.CLK(clknet_leaf_39_io_wbs_clk),
    .D(_00682_),
    .Q(\wfg_drive_pat_top.cfg_end_q[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20369_ (.CLK(clknet_leaf_35_io_wbs_clk),
    .D(_00683_),
    .Q(\wfg_drive_pat_top.cfg_end_q[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20370_ (.CLK(clknet_leaf_38_io_wbs_clk),
    .D(_00684_),
    .Q(\wfg_drive_pat_top.cfg_end_q[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20371_ (.CLK(clknet_leaf_39_io_wbs_clk),
    .D(_00685_),
    .Q(\wfg_drive_pat_top.cfg_end_q[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20372_ (.CLK(clknet_leaf_38_io_wbs_clk),
    .D(_00686_),
    .Q(\wfg_drive_pat_top.cfg_end_q[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20373_ (.CLK(clknet_leaf_38_io_wbs_clk),
    .D(_00687_),
    .Q(\wfg_drive_pat_top.cfg_end_q[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20374_ (.CLK(clknet_leaf_38_io_wbs_clk),
    .D(_00688_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20375_ (.CLK(clknet_leaf_41_io_wbs_clk),
    .D(_00689_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20376_ (.CLK(clknet_leaf_41_io_wbs_clk),
    .D(_00690_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20377_ (.CLK(clknet_leaf_20_io_wbs_clk),
    .D(_00691_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20378_ (.CLK(clknet_leaf_20_io_wbs_clk),
    .D(_00692_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20379_ (.CLK(clknet_leaf_35_io_wbs_clk),
    .D(_00693_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20380_ (.CLK(clknet_leaf_35_io_wbs_clk),
    .D(_00694_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20381_ (.CLK(clknet_leaf_35_io_wbs_clk),
    .D(_00695_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20382_ (.CLK(clknet_leaf_36_io_wbs_clk),
    .D(_00696_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20383_ (.CLK(clknet_leaf_41_io_wbs_clk),
    .D(_00697_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20384_ (.CLK(clknet_leaf_37_io_wbs_clk),
    .D(_00698_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20385_ (.CLK(clknet_leaf_36_io_wbs_clk),
    .D(_00699_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20386_ (.CLK(clknet_leaf_37_io_wbs_clk),
    .D(_00700_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20387_ (.CLK(clknet_leaf_42_io_wbs_clk),
    .D(_00701_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20388_ (.CLK(clknet_leaf_42_io_wbs_clk),
    .D(_00702_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20389_ (.CLK(clknet_leaf_44_io_wbs_clk),
    .D(_00703_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20390_ (.CLK(clknet_leaf_44_io_wbs_clk),
    .D(_00704_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20391_ (.CLK(clknet_leaf_44_io_wbs_clk),
    .D(_00705_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20392_ (.CLK(clknet_leaf_70_io_wbs_clk),
    .D(_00706_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20393_ (.CLK(clknet_leaf_70_io_wbs_clk),
    .D(_00707_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20394_ (.CLK(clknet_leaf_70_io_wbs_clk),
    .D(_00708_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20395_ (.CLK(clknet_leaf_70_io_wbs_clk),
    .D(_00709_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20396_ (.CLK(clknet_leaf_69_io_wbs_clk),
    .D(_00710_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20397_ (.CLK(clknet_leaf_64_io_wbs_clk),
    .D(_00711_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[23] ));
 sky130_fd_sc_hd__dfxtp_1 _20398_ (.CLK(clknet_leaf_64_io_wbs_clk),
    .D(_00712_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[24] ));
 sky130_fd_sc_hd__dfxtp_1 _20399_ (.CLK(clknet_leaf_65_io_wbs_clk),
    .D(_00713_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[25] ));
 sky130_fd_sc_hd__dfxtp_1 _20400_ (.CLK(clknet_leaf_63_io_wbs_clk),
    .D(_00714_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[26] ));
 sky130_fd_sc_hd__dfxtp_1 _20401_ (.CLK(clknet_leaf_65_io_wbs_clk),
    .D(_00715_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[27] ));
 sky130_fd_sc_hd__dfxtp_1 _20402_ (.CLK(clknet_leaf_65_io_wbs_clk),
    .D(_00716_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[28] ));
 sky130_fd_sc_hd__dfxtp_1 _20403_ (.CLK(clknet_leaf_64_io_wbs_clk),
    .D(_00717_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[29] ));
 sky130_fd_sc_hd__dfxtp_1 _20404_ (.CLK(clknet_leaf_68_io_wbs_clk),
    .D(_00718_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[30] ));
 sky130_fd_sc_hd__dfxtp_1 _20405_ (.CLK(clknet_leaf_68_io_wbs_clk),
    .D(_00719_),
    .Q(\wfg_drive_pat_top.patsel0_low_q[31] ));
 sky130_fd_sc_hd__dfxtp_1 _20406_ (.CLK(clknet_leaf_37_io_wbs_clk),
    .D(_00720_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20407_ (.CLK(clknet_leaf_41_io_wbs_clk),
    .D(_00721_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20408_ (.CLK(clknet_leaf_41_io_wbs_clk),
    .D(_00722_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20409_ (.CLK(clknet_leaf_20_io_wbs_clk),
    .D(_00723_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20410_ (.CLK(clknet_leaf_20_io_wbs_clk),
    .D(_00724_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20411_ (.CLK(clknet_leaf_35_io_wbs_clk),
    .D(_00725_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20412_ (.CLK(clknet_leaf_34_io_wbs_clk),
    .D(_00726_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20413_ (.CLK(clknet_leaf_35_io_wbs_clk),
    .D(_00727_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20414_ (.CLK(clknet_leaf_36_io_wbs_clk),
    .D(_00728_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20415_ (.CLK(clknet_leaf_37_io_wbs_clk),
    .D(_00729_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20416_ (.CLK(clknet_leaf_37_io_wbs_clk),
    .D(_00730_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20417_ (.CLK(clknet_leaf_36_io_wbs_clk),
    .D(_00731_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20418_ (.CLK(clknet_leaf_37_io_wbs_clk),
    .D(_00732_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20419_ (.CLK(clknet_leaf_42_io_wbs_clk),
    .D(_00733_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20420_ (.CLK(clknet_leaf_42_io_wbs_clk),
    .D(_00734_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20421_ (.CLK(clknet_leaf_43_io_wbs_clk),
    .D(_00735_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20422_ (.CLK(clknet_leaf_43_io_wbs_clk),
    .D(_00736_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20423_ (.CLK(clknet_leaf_44_io_wbs_clk),
    .D(_00737_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20424_ (.CLK(clknet_leaf_44_io_wbs_clk),
    .D(_00738_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20425_ (.CLK(clknet_leaf_70_io_wbs_clk),
    .D(_00739_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20426_ (.CLK(clknet_leaf_69_io_wbs_clk),
    .D(_00740_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20427_ (.CLK(clknet_leaf_69_io_wbs_clk),
    .D(_00741_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20428_ (.CLK(clknet_leaf_69_io_wbs_clk),
    .D(_00742_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20429_ (.CLK(clknet_leaf_64_io_wbs_clk),
    .D(_00743_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[23] ));
 sky130_fd_sc_hd__dfxtp_1 _20430_ (.CLK(clknet_leaf_64_io_wbs_clk),
    .D(_00744_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[24] ));
 sky130_fd_sc_hd__dfxtp_1 _20431_ (.CLK(clknet_leaf_65_io_wbs_clk),
    .D(_00745_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[25] ));
 sky130_fd_sc_hd__dfxtp_1 _20432_ (.CLK(clknet_leaf_63_io_wbs_clk),
    .D(_00746_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[26] ));
 sky130_fd_sc_hd__dfxtp_1 _20433_ (.CLK(clknet_leaf_65_io_wbs_clk),
    .D(_00747_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[27] ));
 sky130_fd_sc_hd__dfxtp_1 _20434_ (.CLK(clknet_leaf_65_io_wbs_clk),
    .D(_00748_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[28] ));
 sky130_fd_sc_hd__dfxtp_1 _20435_ (.CLK(clknet_leaf_63_io_wbs_clk),
    .D(_00749_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[29] ));
 sky130_fd_sc_hd__dfxtp_1 _20436_ (.CLK(clknet_leaf_63_io_wbs_clk),
    .D(_00750_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[30] ));
 sky130_fd_sc_hd__dfxtp_1 _20437_ (.CLK(clknet_leaf_68_io_wbs_clk),
    .D(_00751_),
    .Q(\wfg_drive_pat_top.patsel1_high_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _20438_ (.CLK(clknet_leaf_11_io_wbs_clk),
    .D(_00024_),
    .RESET_B(_00143_),
    .Q(\wfg_subcore_top.wfg_subcore.subcycle_count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _20439_ (.CLK(clknet_leaf_11_io_wbs_clk),
    .D(_00031_),
    .RESET_B(_00144_),
    .Q(\wfg_subcore_top.wfg_subcore.subcycle_count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _20440_ (.CLK(clknet_leaf_10_io_wbs_clk),
    .D(_00032_),
    .RESET_B(_00145_),
    .Q(\wfg_subcore_top.wfg_subcore.subcycle_count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _20441_ (.CLK(clknet_leaf_10_io_wbs_clk),
    .D(_00033_),
    .RESET_B(_00146_),
    .Q(\wfg_subcore_top.wfg_subcore.subcycle_count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _20442_ (.CLK(clknet_leaf_12_io_wbs_clk),
    .D(_00034_),
    .RESET_B(_00147_),
    .Q(\wfg_subcore_top.wfg_subcore.subcycle_count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _20443_ (.CLK(clknet_leaf_12_io_wbs_clk),
    .D(_00035_),
    .RESET_B(_00148_),
    .Q(\wfg_subcore_top.wfg_subcore.subcycle_count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _20444_ (.CLK(clknet_leaf_12_io_wbs_clk),
    .D(_00036_),
    .RESET_B(_00149_),
    .Q(\wfg_subcore_top.wfg_subcore.subcycle_count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _20445_ (.CLK(clknet_leaf_90_io_wbs_clk),
    .D(_00037_),
    .RESET_B(_00150_),
    .Q(\wfg_subcore_top.wfg_subcore.subcycle_count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _20446_ (.CLK(clknet_leaf_88_io_wbs_clk),
    .D(_00038_),
    .RESET_B(_00151_),
    .Q(\wfg_subcore_top.wfg_subcore.subcycle_count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _20447_ (.CLK(clknet_leaf_15_io_wbs_clk),
    .D(_00039_),
    .RESET_B(_00152_),
    .Q(\wfg_subcore_top.wfg_subcore.subcycle_count[9] ));
 sky130_fd_sc_hd__dfrtp_1 _20448_ (.CLK(clknet_leaf_88_io_wbs_clk),
    .D(_00025_),
    .RESET_B(_00153_),
    .Q(\wfg_subcore_top.wfg_subcore.subcycle_count[10] ));
 sky130_fd_sc_hd__dfrtp_1 _20449_ (.CLK(clknet_leaf_15_io_wbs_clk),
    .D(_00026_),
    .RESET_B(_00154_),
    .Q(\wfg_subcore_top.wfg_subcore.subcycle_count[11] ));
 sky130_fd_sc_hd__dfrtp_1 _20450_ (.CLK(clknet_leaf_87_io_wbs_clk),
    .D(_00027_),
    .RESET_B(_00155_),
    .Q(\wfg_subcore_top.wfg_subcore.subcycle_count[12] ));
 sky130_fd_sc_hd__dfrtp_1 _20451_ (.CLK(clknet_leaf_86_io_wbs_clk),
    .D(_00028_),
    .RESET_B(_00156_),
    .Q(\wfg_subcore_top.wfg_subcore.subcycle_count[13] ));
 sky130_fd_sc_hd__dfrtp_1 _20452_ (.CLK(clknet_leaf_86_io_wbs_clk),
    .D(_00029_),
    .RESET_B(_00157_),
    .Q(\wfg_subcore_top.wfg_subcore.subcycle_count[14] ));
 sky130_fd_sc_hd__dfrtp_1 _20453_ (.CLK(clknet_leaf_87_io_wbs_clk),
    .D(_00030_),
    .RESET_B(_00158_),
    .Q(\wfg_subcore_top.wfg_subcore.subcycle_count[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20454_ (.CLK(clknet_leaf_101_io_wbs_clk),
    .D(_00752_),
    .Q(\wfg_stim_sine_top.wbs_ack_o ));
 sky130_fd_sc_hd__dfrtp_1 _20455_ (.CLK(clknet_leaf_15_io_wbs_clk),
    .D(_00753_),
    .RESET_B(_00159_),
    .Q(\wfg_subcore_top.wfg_subcore.sync_count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _20456_ (.CLK(clknet_leaf_14_io_wbs_clk),
    .D(_00754_),
    .RESET_B(_00160_),
    .Q(\wfg_subcore_top.wfg_subcore.sync_count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _20457_ (.CLK(clknet_leaf_12_io_wbs_clk),
    .D(_00755_),
    .RESET_B(_00161_),
    .Q(\wfg_subcore_top.wfg_subcore.sync_count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _20458_ (.CLK(clknet_leaf_12_io_wbs_clk),
    .D(_00756_),
    .RESET_B(_00162_),
    .Q(\wfg_subcore_top.wfg_subcore.sync_count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _20459_ (.CLK(clknet_leaf_13_io_wbs_clk),
    .D(_00757_),
    .RESET_B(_00163_),
    .Q(\wfg_subcore_top.wfg_subcore.sync_count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _20460_ (.CLK(clknet_leaf_13_io_wbs_clk),
    .D(_00758_),
    .RESET_B(_00164_),
    .Q(\wfg_subcore_top.wfg_subcore.sync_count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _20461_ (.CLK(clknet_leaf_10_io_wbs_clk),
    .D(_00759_),
    .RESET_B(_00165_),
    .Q(\wfg_subcore_top.wfg_subcore.sync_count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _20462_ (.CLK(clknet_leaf_12_io_wbs_clk),
    .D(_00760_),
    .RESET_B(_00166_),
    .Q(\wfg_subcore_top.wfg_subcore.sync_count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _20463_ (.CLK(clknet_leaf_14_io_wbs_clk),
    .D(_00761_),
    .RESET_B(_00167_),
    .Q(\wfg_subcore_top.wfg_subcore.temp_subcycle ));
 sky130_fd_sc_hd__dfrtp_1 _20464_ (.CLK(clknet_leaf_15_io_wbs_clk),
    .D(_00762_),
    .RESET_B(_00168_),
    .Q(\wfg_subcore_top.wfg_subcore.temp_sync ));
 sky130_fd_sc_hd__dfxtp_1 _20465_ (.CLK(clknet_leaf_86_io_wbs_clk),
    .D(_00763_),
    .Q(\wfg_subcore_top.wfg_subcore.subcycle_dly ));
 sky130_fd_sc_hd__dfxtp_1 _20466_ (.CLK(clknet_leaf_15_io_wbs_clk),
    .D(_00764_),
    .Q(\wfg_subcore_top.wfg_subcore.sync_dly ));
 sky130_fd_sc_hd__dfrtp_2 _20467_ (.CLK(clknet_leaf_16_io_wbs_clk),
    .D(_00765_),
    .RESET_B(_00169_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[0] ));
 sky130_fd_sc_hd__dfrtp_1 _20468_ (.CLK(clknet_leaf_86_io_wbs_clk),
    .D(_00766_),
    .RESET_B(_00170_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[1] ));
 sky130_fd_sc_hd__dfrtp_1 _20469_ (.CLK(clknet_leaf_74_io_wbs_clk),
    .D(_00767_),
    .RESET_B(_00171_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[2] ));
 sky130_fd_sc_hd__dfrtp_1 _20470_ (.CLK(clknet_leaf_74_io_wbs_clk),
    .D(_00768_),
    .RESET_B(_00172_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[3] ));
 sky130_fd_sc_hd__dfrtp_1 _20471_ (.CLK(clknet_leaf_74_io_wbs_clk),
    .D(_00769_),
    .RESET_B(_00173_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[4] ));
 sky130_fd_sc_hd__dfrtp_1 _20472_ (.CLK(clknet_leaf_40_io_wbs_clk),
    .D(_00770_),
    .RESET_B(_00174_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[5] ));
 sky130_fd_sc_hd__dfrtp_1 _20473_ (.CLK(clknet_leaf_40_io_wbs_clk),
    .D(_00771_),
    .RESET_B(_00175_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[6] ));
 sky130_fd_sc_hd__dfrtp_1 _20474_ (.CLK(clknet_leaf_40_io_wbs_clk),
    .D(_00772_),
    .RESET_B(_00176_),
    .Q(\wfg_drive_pat_top.wfg_drive_pat.wfg_subcore_subcycle_cnt_i[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20475_ (.CLK(clknet_leaf_92_io_wbs_clk),
    .D(_00773_),
    .Q(\wfg_stim_sine_top.wbs_dat_o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20476_ (.CLK(clknet_leaf_93_io_wbs_clk),
    .D(_00774_),
    .Q(\wfg_stim_sine_top.wbs_dat_o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20477_ (.CLK(clknet_leaf_93_io_wbs_clk),
    .D(_00775_),
    .Q(\wfg_stim_sine_top.wbs_dat_o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20478_ (.CLK(clknet_leaf_93_io_wbs_clk),
    .D(_00776_),
    .Q(\wfg_stim_sine_top.wbs_dat_o[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20479_ (.CLK(clknet_leaf_93_io_wbs_clk),
    .D(_00777_),
    .Q(\wfg_stim_sine_top.wbs_dat_o[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20480_ (.CLK(clknet_leaf_93_io_wbs_clk),
    .D(_00778_),
    .Q(\wfg_stim_sine_top.wbs_dat_o[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20481_ (.CLK(clknet_leaf_93_io_wbs_clk),
    .D(_00779_),
    .Q(\wfg_stim_sine_top.wbs_dat_o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20482_ (.CLK(clknet_leaf_92_io_wbs_clk),
    .D(_00780_),
    .Q(\wfg_stim_sine_top.wbs_dat_o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20483_ (.CLK(clknet_leaf_93_io_wbs_clk),
    .D(_00781_),
    .Q(\wfg_stim_sine_top.wbs_dat_o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20484_ (.CLK(clknet_leaf_93_io_wbs_clk),
    .D(_00782_),
    .Q(\wfg_stim_sine_top.wbs_dat_o[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20485_ (.CLK(clknet_leaf_81_io_wbs_clk),
    .D(_00783_),
    .Q(\wfg_stim_sine_top.wbs_dat_o[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20486_ (.CLK(clknet_leaf_94_io_wbs_clk),
    .D(_00784_),
    .Q(\wfg_stim_sine_top.wbs_dat_o[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20487_ (.CLK(clknet_leaf_81_io_wbs_clk),
    .D(_00785_),
    .Q(\wfg_stim_sine_top.wbs_dat_o[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20488_ (.CLK(clknet_leaf_81_io_wbs_clk),
    .D(_00786_),
    .Q(\wfg_stim_sine_top.wbs_dat_o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20489_ (.CLK(clknet_leaf_81_io_wbs_clk),
    .D(_00787_),
    .Q(\wfg_stim_sine_top.wbs_dat_o[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20490_ (.CLK(clknet_leaf_94_io_wbs_clk),
    .D(_00788_),
    .Q(\wfg_stim_sine_top.wbs_dat_o[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20491_ (.CLK(clknet_leaf_81_io_wbs_clk),
    .D(_00789_),
    .Q(\wfg_stim_sine_top.wbs_dat_o[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20492_ (.CLK(clknet_leaf_81_io_wbs_clk),
    .D(_00790_),
    .Q(\wfg_stim_sine_top.wbs_dat_o[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20493_ (.CLK(clknet_leaf_11_io_wbs_clk),
    .D(_00791_),
    .Q(\wfg_subcore_top.cfg_subcycle_q[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20494_ (.CLK(clknet_leaf_11_io_wbs_clk),
    .D(_00792_),
    .Q(\wfg_subcore_top.cfg_subcycle_q[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20495_ (.CLK(clknet_leaf_90_io_wbs_clk),
    .D(_00793_),
    .Q(\wfg_subcore_top.cfg_subcycle_q[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20496_ (.CLK(clknet_leaf_90_io_wbs_clk),
    .D(_00794_),
    .Q(\wfg_subcore_top.cfg_subcycle_q[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20497_ (.CLK(clknet_leaf_12_io_wbs_clk),
    .D(_00795_),
    .Q(\wfg_subcore_top.cfg_subcycle_q[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20498_ (.CLK(clknet_leaf_12_io_wbs_clk),
    .D(_00796_),
    .Q(\wfg_subcore_top.cfg_subcycle_q[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20499_ (.CLK(clknet_leaf_90_io_wbs_clk),
    .D(_00797_),
    .Q(\wfg_subcore_top.cfg_subcycle_q[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20500_ (.CLK(clknet_leaf_90_io_wbs_clk),
    .D(_00798_),
    .Q(\wfg_subcore_top.cfg_subcycle_q[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20501_ (.CLK(clknet_leaf_88_io_wbs_clk),
    .D(_00799_),
    .Q(\wfg_subcore_top.cfg_subcycle_q[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20502_ (.CLK(clknet_leaf_88_io_wbs_clk),
    .D(_00800_),
    .Q(\wfg_subcore_top.cfg_subcycle_q[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20503_ (.CLK(clknet_leaf_88_io_wbs_clk),
    .D(_00801_),
    .Q(\wfg_subcore_top.cfg_subcycle_q[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20504_ (.CLK(clknet_leaf_88_io_wbs_clk),
    .D(_00802_),
    .Q(\wfg_subcore_top.cfg_subcycle_q[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20505_ (.CLK(clknet_leaf_88_io_wbs_clk),
    .D(_00803_),
    .Q(\wfg_subcore_top.cfg_subcycle_q[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20506_ (.CLK(clknet_leaf_87_io_wbs_clk),
    .D(_00804_),
    .Q(\wfg_subcore_top.cfg_subcycle_q[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20507_ (.CLK(clknet_leaf_87_io_wbs_clk),
    .D(_00805_),
    .Q(\wfg_subcore_top.cfg_subcycle_q[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20508_ (.CLK(clknet_leaf_88_io_wbs_clk),
    .D(_00806_),
    .Q(\wfg_subcore_top.cfg_subcycle_q[23] ));
 sky130_fd_sc_hd__dfxtp_1 _20509_ (.CLK(clknet_leaf_12_io_wbs_clk),
    .D(_00807_),
    .Q(\wfg_subcore_top.cfg_sync_q[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20510_ (.CLK(clknet_leaf_12_io_wbs_clk),
    .D(_00808_),
    .Q(\wfg_subcore_top.cfg_sync_q[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20511_ (.CLK(clknet_leaf_12_io_wbs_clk),
    .D(_00809_),
    .Q(\wfg_subcore_top.cfg_sync_q[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20512_ (.CLK(clknet_leaf_12_io_wbs_clk),
    .D(_00810_),
    .Q(\wfg_subcore_top.cfg_sync_q[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20513_ (.CLK(clknet_leaf_11_io_wbs_clk),
    .D(_00811_),
    .Q(\wfg_subcore_top.cfg_sync_q[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20514_ (.CLK(clknet_leaf_11_io_wbs_clk),
    .D(_00812_),
    .Q(\wfg_subcore_top.cfg_sync_q[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20515_ (.CLK(clknet_leaf_11_io_wbs_clk),
    .D(_00813_),
    .Q(\wfg_subcore_top.cfg_sync_q[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20516_ (.CLK(clknet_leaf_11_io_wbs_clk),
    .D(_00814_),
    .Q(\wfg_subcore_top.cfg_sync_q[7] ));
 sky130_fd_sc_hd__dfxtp_2 _20517_ (.CLK(clknet_leaf_91_io_wbs_clk),
    .D(_00815_),
    .Q(\wfg_subcore_top.active_o ));
 sky130_fd_sc_hd__dfxtp_1 _20518_ (.CLK(clknet_leaf_101_io_wbs_clk),
    .D(_00816_),
    .Q(\wfg_drive_spi_top.wbs_ack_o ));
 sky130_fd_sc_hd__dfxtp_1 _20519_ (.CLK(clknet_leaf_14_io_wbs_clk),
    .D(_00817_),
    .Q(\wfg_drive_spi_top.wbs_dat_o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20520_ (.CLK(clknet_leaf_14_io_wbs_clk),
    .D(_00818_),
    .Q(\wfg_drive_spi_top.wbs_dat_o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20521_ (.CLK(clknet_leaf_14_io_wbs_clk),
    .D(_00819_),
    .Q(\wfg_drive_spi_top.wbs_dat_o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20522_ (.CLK(clknet_leaf_14_io_wbs_clk),
    .D(_00820_),
    .Q(\wfg_drive_spi_top.wbs_dat_o[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20523_ (.CLK(clknet_leaf_13_io_wbs_clk),
    .D(_00821_),
    .Q(\wfg_drive_spi_top.wbs_dat_o[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20524_ (.CLK(clknet_leaf_13_io_wbs_clk),
    .D(_00822_),
    .Q(\wfg_drive_spi_top.wbs_dat_o[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20525_ (.CLK(clknet_leaf_19_io_wbs_clk),
    .D(_00823_),
    .Q(\wfg_drive_spi_top.wbs_dat_o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20526_ (.CLK(clknet_leaf_18_io_wbs_clk),
    .D(_00824_),
    .Q(\wfg_drive_spi_top.wbs_dat_o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20527_ (.CLK(clknet_leaf_14_io_wbs_clk),
    .D(_00825_),
    .Q(\wfg_interconnect_top.ctrl_en_q ));
 sky130_fd_sc_hd__dfxtp_4 _20528_ (.CLK(clknet_leaf_17_io_wbs_clk),
    .D(_00826_),
    .Q(\wfg_interconnect_top.driver0_select_q[0] ));
 sky130_fd_sc_hd__dfxtp_4 _20529_ (.CLK(clknet_leaf_17_io_wbs_clk),
    .D(_00827_),
    .Q(\wfg_interconnect_top.driver0_select_q[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20530_ (.CLK(clknet_leaf_14_io_wbs_clk),
    .D(_00828_),
    .Q(\wfg_interconnect_top.driver1_select_q[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20531_ (.CLK(clknet_leaf_14_io_wbs_clk),
    .D(_00829_),
    .Q(\wfg_interconnect_top.driver1_select_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _20532_ (.CLK(clknet_leaf_74_io_wbs_clk),
    .D(_00830_),
    .RESET_B(_00177_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[0] ));
 sky130_fd_sc_hd__dfrtp_1 _20533_ (.CLK(clknet_leaf_74_io_wbs_clk),
    .D(_00831_),
    .RESET_B(_00178_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[1] ));
 sky130_fd_sc_hd__dfrtp_1 _20534_ (.CLK(clknet_leaf_74_io_wbs_clk),
    .D(_00832_),
    .RESET_B(_00179_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[2] ));
 sky130_fd_sc_hd__dfrtp_1 _20535_ (.CLK(clknet_leaf_74_io_wbs_clk),
    .D(_00833_),
    .RESET_B(_00180_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[3] ));
 sky130_fd_sc_hd__dfrtp_1 _20536_ (.CLK(clknet_leaf_73_io_wbs_clk),
    .D(_00834_),
    .RESET_B(_00181_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[4] ));
 sky130_fd_sc_hd__dfrtp_1 _20537_ (.CLK(clknet_leaf_73_io_wbs_clk),
    .D(_00835_),
    .RESET_B(_00182_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[5] ));
 sky130_fd_sc_hd__dfrtp_1 _20538_ (.CLK(clknet_leaf_73_io_wbs_clk),
    .D(_00836_),
    .RESET_B(_00183_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[6] ));
 sky130_fd_sc_hd__dfrtp_1 _20539_ (.CLK(clknet_leaf_73_io_wbs_clk),
    .D(_00837_),
    .RESET_B(_00184_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[7] ));
 sky130_fd_sc_hd__dfrtp_1 _20540_ (.CLK(clknet_leaf_73_io_wbs_clk),
    .D(_00838_),
    .RESET_B(_00185_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[8] ));
 sky130_fd_sc_hd__dfrtp_1 _20541_ (.CLK(clknet_leaf_71_io_wbs_clk),
    .D(_00839_),
    .RESET_B(_00186_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[9] ));
 sky130_fd_sc_hd__dfrtp_1 _20542_ (.CLK(clknet_leaf_71_io_wbs_clk),
    .D(_00840_),
    .RESET_B(_00187_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[10] ));
 sky130_fd_sc_hd__dfrtp_1 _20543_ (.CLK(clknet_leaf_72_io_wbs_clk),
    .D(_00841_),
    .RESET_B(_00188_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[11] ));
 sky130_fd_sc_hd__dfrtp_1 _20544_ (.CLK(clknet_leaf_72_io_wbs_clk),
    .D(_00842_),
    .RESET_B(_00189_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[12] ));
 sky130_fd_sc_hd__dfrtp_1 _20545_ (.CLK(clknet_leaf_72_io_wbs_clk),
    .D(_00843_),
    .RESET_B(_00190_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[13] ));
 sky130_fd_sc_hd__dfrtp_1 _20546_ (.CLK(clknet_leaf_72_io_wbs_clk),
    .D(_00844_),
    .RESET_B(_00191_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[14] ));
 sky130_fd_sc_hd__dfrtp_1 _20547_ (.CLK(clknet_leaf_73_io_wbs_clk),
    .D(_00845_),
    .RESET_B(_00192_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[15] ));
 sky130_fd_sc_hd__dfrtp_1 _20548_ (.CLK(clknet_leaf_73_io_wbs_clk),
    .D(_00846_),
    .RESET_B(_00193_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[16] ));
 sky130_fd_sc_hd__dfrtp_1 _20549_ (.CLK(clknet_leaf_74_io_wbs_clk),
    .D(_00847_),
    .RESET_B(_00194_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.overflow_chk[17] ));
 sky130_fd_sc_hd__dfrtp_4 _20550_ (.CLK(clknet_leaf_9_io_wbs_clk),
    .D(_00848_),
    .RESET_B(_00195_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.cur_state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _20551_ (.CLK(clknet_leaf_9_io_wbs_clk),
    .D(_00849_),
    .RESET_B(_00196_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.cur_state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _20552_ (.CLK(clknet_leaf_88_io_wbs_clk),
    .D(_00850_),
    .RESET_B(_00197_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.cur_state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20553_ (.CLK(clknet_leaf_101_io_wbs_clk),
    .D(_00851_),
    .Q(\wfg_stim_mem_top.wbs_ack_o ));
 sky130_fd_sc_hd__dfrtp_4 _20554_ (.CLK(clknet_leaf_75_io_wbs_clk),
    .D(_00852_),
    .RESET_B(_00198_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.sin_17[0] ));
 sky130_fd_sc_hd__dfrtp_4 _20555_ (.CLK(clknet_leaf_14_io_wbs_clk),
    .D(_00853_),
    .RESET_B(_00199_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.sin_17[1] ));
 sky130_fd_sc_hd__dfrtp_1 _20556_ (.CLK(clknet_leaf_86_io_wbs_clk),
    .D(_00854_),
    .RESET_B(_00200_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.sin_17[2] ));
 sky130_fd_sc_hd__dfrtp_4 _20557_ (.CLK(clknet_leaf_86_io_wbs_clk),
    .D(_00855_),
    .RESET_B(_00201_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.sin_17[3] ));
 sky130_fd_sc_hd__dfrtp_1 _20558_ (.CLK(clknet_leaf_85_io_wbs_clk),
    .D(_00856_),
    .RESET_B(_00202_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.sin_17[4] ));
 sky130_fd_sc_hd__dfrtp_4 _20559_ (.CLK(clknet_leaf_86_io_wbs_clk),
    .D(_00857_),
    .RESET_B(_00203_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.sin_17[5] ));
 sky130_fd_sc_hd__dfrtp_4 _20560_ (.CLK(clknet_leaf_85_io_wbs_clk),
    .D(_00858_),
    .RESET_B(_00204_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.sin_17[6] ));
 sky130_fd_sc_hd__dfrtp_1 _20561_ (.CLK(clknet_leaf_86_io_wbs_clk),
    .D(_00859_),
    .RESET_B(_00205_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.sin_17[7] ));
 sky130_fd_sc_hd__dfrtp_1 _20562_ (.CLK(clknet_leaf_86_io_wbs_clk),
    .D(_00860_),
    .RESET_B(_00206_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.sin_17[8] ));
 sky130_fd_sc_hd__dfrtp_4 _20563_ (.CLK(clknet_leaf_86_io_wbs_clk),
    .D(_00861_),
    .RESET_B(_00207_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.sin_17[9] ));
 sky130_fd_sc_hd__dfrtp_4 _20564_ (.CLK(clknet_leaf_74_io_wbs_clk),
    .D(_00862_),
    .RESET_B(_00208_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.sin_17[10] ));
 sky130_fd_sc_hd__dfrtp_4 _20565_ (.CLK(clknet_leaf_75_io_wbs_clk),
    .D(_00863_),
    .RESET_B(_00209_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.sin_17[11] ));
 sky130_fd_sc_hd__dfrtp_4 _20566_ (.CLK(clknet_leaf_74_io_wbs_clk),
    .D(_00864_),
    .RESET_B(_00210_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.sin_17[12] ));
 sky130_fd_sc_hd__dfrtp_4 _20567_ (.CLK(clknet_leaf_75_io_wbs_clk),
    .D(_00865_),
    .RESET_B(_00211_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.sin_17[13] ));
 sky130_fd_sc_hd__dfrtp_4 _20568_ (.CLK(clknet_leaf_75_io_wbs_clk),
    .D(_00866_),
    .RESET_B(_00212_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.sin_17[14] ));
 sky130_fd_sc_hd__dfrtp_4 _20569_ (.CLK(clknet_leaf_75_io_wbs_clk),
    .D(_00867_),
    .RESET_B(_00213_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.sin_17[15] ));
 sky130_fd_sc_hd__dfrtp_1 _20570_ (.CLK(clknet_leaf_76_io_wbs_clk),
    .D(_00868_),
    .RESET_B(_00214_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.sin_17[16] ));
 sky130_fd_sc_hd__dfrtp_1 _20571_ (.CLK(clknet_leaf_41_io_wbs_clk),
    .D(_00869_),
    .RESET_B(_00215_),
    .Q(\wfg_interconnect_top.stimulus_0[0] ));
 sky130_fd_sc_hd__dfrtp_1 _20572_ (.CLK(clknet_leaf_73_io_wbs_clk),
    .D(_00870_),
    .RESET_B(_00216_),
    .Q(\wfg_interconnect_top.stimulus_0[1] ));
 sky130_fd_sc_hd__dfrtp_1 _20573_ (.CLK(clknet_leaf_73_io_wbs_clk),
    .D(_00871_),
    .RESET_B(_00217_),
    .Q(\wfg_interconnect_top.stimulus_0[2] ));
 sky130_fd_sc_hd__dfrtp_1 _20574_ (.CLK(clknet_leaf_73_io_wbs_clk),
    .D(_00872_),
    .RESET_B(_00218_),
    .Q(\wfg_interconnect_top.stimulus_0[3] ));
 sky130_fd_sc_hd__dfrtp_1 _20575_ (.CLK(clknet_leaf_73_io_wbs_clk),
    .D(_00873_),
    .RESET_B(_00219_),
    .Q(\wfg_interconnect_top.stimulus_0[4] ));
 sky130_fd_sc_hd__dfrtp_1 _20576_ (.CLK(clknet_leaf_73_io_wbs_clk),
    .D(_00874_),
    .RESET_B(_00220_),
    .Q(\wfg_interconnect_top.stimulus_0[5] ));
 sky130_fd_sc_hd__dfrtp_1 _20577_ (.CLK(clknet_leaf_71_io_wbs_clk),
    .D(_00875_),
    .RESET_B(_00221_),
    .Q(\wfg_interconnect_top.stimulus_0[6] ));
 sky130_fd_sc_hd__dfrtp_1 _20578_ (.CLK(clknet_leaf_71_io_wbs_clk),
    .D(_00876_),
    .RESET_B(_00222_),
    .Q(\wfg_interconnect_top.stimulus_0[7] ));
 sky130_fd_sc_hd__dfrtp_1 _20579_ (.CLK(clknet_leaf_71_io_wbs_clk),
    .D(_00877_),
    .RESET_B(_00223_),
    .Q(\wfg_interconnect_top.stimulus_0[8] ));
 sky130_fd_sc_hd__dfrtp_1 _20580_ (.CLK(clknet_leaf_71_io_wbs_clk),
    .D(_00878_),
    .RESET_B(_00224_),
    .Q(\wfg_interconnect_top.stimulus_0[9] ));
 sky130_fd_sc_hd__dfrtp_1 _20581_ (.CLK(clknet_leaf_71_io_wbs_clk),
    .D(_00879_),
    .RESET_B(_00225_),
    .Q(\wfg_interconnect_top.stimulus_0[10] ));
 sky130_fd_sc_hd__dfrtp_1 _20582_ (.CLK(clknet_leaf_70_io_wbs_clk),
    .D(_00880_),
    .RESET_B(_00226_),
    .Q(\wfg_interconnect_top.stimulus_0[11] ));
 sky130_fd_sc_hd__dfrtp_2 _20583_ (.CLK(clknet_leaf_71_io_wbs_clk),
    .D(_00881_),
    .RESET_B(_00227_),
    .Q(\wfg_interconnect_top.stimulus_0[12] ));
 sky130_fd_sc_hd__dfrtp_1 _20584_ (.CLK(clknet_leaf_69_io_wbs_clk),
    .D(_00882_),
    .RESET_B(_00228_),
    .Q(\wfg_interconnect_top.stimulus_0[13] ));
 sky130_fd_sc_hd__dfrtp_1 _20585_ (.CLK(clknet_leaf_67_io_wbs_clk),
    .D(_00883_),
    .RESET_B(_00229_),
    .Q(\wfg_interconnect_top.stimulus_0[14] ));
 sky130_fd_sc_hd__dfrtp_1 _20586_ (.CLK(clknet_leaf_67_io_wbs_clk),
    .D(_00884_),
    .RESET_B(_00230_),
    .Q(\wfg_interconnect_top.stimulus_0[15] ));
 sky130_fd_sc_hd__dfrtp_2 _20587_ (.CLK(clknet_leaf_71_io_wbs_clk),
    .D(_00885_),
    .RESET_B(_00231_),
    .Q(\wfg_interconnect_top.stimulus_0[16] ));
 sky130_fd_sc_hd__dfrtp_1 _20588_ (.CLK(clknet_leaf_41_io_wbs_clk),
    .D(_00886_),
    .RESET_B(_00232_),
    .Q(\wfg_interconnect_top.stimulus_0[17] ));
 sky130_fd_sc_hd__dfrtp_2 _20589_ (.CLK(clknet_leaf_22_io_wbs_clk),
    .D(_00887_),
    .RESET_B(_00233_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.x[0] ));
 sky130_fd_sc_hd__dfrtp_4 _20590_ (.CLK(clknet_leaf_22_io_wbs_clk),
    .D(_00888_),
    .RESET_B(_00234_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.x[1] ));
 sky130_fd_sc_hd__dfstp_2 _20591_ (.CLK(clknet_leaf_22_io_wbs_clk),
    .D(_00889_),
    .SET_B(_00235_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.x[2] ));
 sky130_fd_sc_hd__dfrtp_4 _20592_ (.CLK(clknet_leaf_22_io_wbs_clk),
    .D(_00890_),
    .RESET_B(_00236_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.x[3] ));
 sky130_fd_sc_hd__dfstp_2 _20593_ (.CLK(clknet_leaf_27_io_wbs_clk),
    .D(_00891_),
    .SET_B(_00237_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.x[4] ));
 sky130_fd_sc_hd__dfstp_2 _20594_ (.CLK(clknet_leaf_27_io_wbs_clk),
    .D(_00892_),
    .SET_B(_00238_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.x[5] ));
 sky130_fd_sc_hd__dfstp_2 _20595_ (.CLK(clknet_leaf_27_io_wbs_clk),
    .D(_00893_),
    .SET_B(_00239_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.x[6] ));
 sky130_fd_sc_hd__dfrtp_4 _20596_ (.CLK(clknet_leaf_27_io_wbs_clk),
    .D(_00894_),
    .RESET_B(_00240_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.x[7] ));
 sky130_fd_sc_hd__dfstp_2 _20597_ (.CLK(clknet_leaf_26_io_wbs_clk),
    .D(_00895_),
    .SET_B(_00241_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.x[8] ));
 sky130_fd_sc_hd__dfstp_2 _20598_ (.CLK(clknet_leaf_29_io_wbs_clk),
    .D(_00896_),
    .SET_B(_00242_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.x[9] ));
 sky130_fd_sc_hd__dfrtp_4 _20599_ (.CLK(clknet_leaf_26_io_wbs_clk),
    .D(_00897_),
    .RESET_B(_00243_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.x[10] ));
 sky130_fd_sc_hd__dfstp_2 _20600_ (.CLK(clknet_leaf_26_io_wbs_clk),
    .D(_00898_),
    .SET_B(_00244_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.x[11] ));
 sky130_fd_sc_hd__dfstp_2 _20601_ (.CLK(clknet_leaf_25_io_wbs_clk),
    .D(_00899_),
    .SET_B(_00245_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.x[12] ));
 sky130_fd_sc_hd__dfrtp_4 _20602_ (.CLK(clknet_leaf_25_io_wbs_clk),
    .D(_00900_),
    .RESET_B(_00246_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.x[13] ));
 sky130_fd_sc_hd__dfrtp_4 _20603_ (.CLK(clknet_leaf_25_io_wbs_clk),
    .D(_00901_),
    .RESET_B(_00247_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.x[14] ));
 sky130_fd_sc_hd__dfstp_2 _20604_ (.CLK(clknet_leaf_25_io_wbs_clk),
    .D(_00902_),
    .SET_B(_00248_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.x[15] ));
 sky130_fd_sc_hd__dfrtp_4 _20605_ (.CLK(clknet_leaf_25_io_wbs_clk),
    .D(_00903_),
    .RESET_B(_00249_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.x[16] ));
 sky130_fd_sc_hd__dfrtp_2 _20606_ (.CLK(clknet_leaf_22_io_wbs_clk),
    .D(_00904_),
    .RESET_B(_00250_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.y[0] ));
 sky130_fd_sc_hd__dfrtp_4 _20607_ (.CLK(clknet_leaf_23_io_wbs_clk),
    .D(_00905_),
    .RESET_B(_00251_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.y[1] ));
 sky130_fd_sc_hd__dfrtp_2 _20608_ (.CLK(clknet_leaf_23_io_wbs_clk),
    .D(_00906_),
    .RESET_B(_00252_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.y[2] ));
 sky130_fd_sc_hd__dfrtp_2 _20609_ (.CLK(clknet_leaf_9_io_wbs_clk),
    .D(_00907_),
    .RESET_B(_00253_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.y[3] ));
 sky130_fd_sc_hd__dfrtp_4 _20610_ (.CLK(clknet_leaf_8_io_wbs_clk),
    .D(_00908_),
    .RESET_B(_00254_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.y[4] ));
 sky130_fd_sc_hd__dfrtp_2 _20611_ (.CLK(clknet_leaf_8_io_wbs_clk),
    .D(_00909_),
    .RESET_B(_00255_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.y[5] ));
 sky130_fd_sc_hd__dfrtp_4 _20612_ (.CLK(clknet_leaf_8_io_wbs_clk),
    .D(_00910_),
    .RESET_B(_00256_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.y[6] ));
 sky130_fd_sc_hd__dfrtp_4 _20613_ (.CLK(clknet_leaf_8_io_wbs_clk),
    .D(_00911_),
    .RESET_B(_00257_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.y[7] ));
 sky130_fd_sc_hd__dfrtp_4 _20614_ (.CLK(clknet_leaf_6_io_wbs_clk),
    .D(_00912_),
    .RESET_B(_00258_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.y[8] ));
 sky130_fd_sc_hd__dfrtp_4 _20615_ (.CLK(clknet_leaf_6_io_wbs_clk),
    .D(_00913_),
    .RESET_B(_00259_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.y[9] ));
 sky130_fd_sc_hd__dfrtp_4 _20616_ (.CLK(clknet_leaf_7_io_wbs_clk),
    .D(_00914_),
    .RESET_B(_00260_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.y[10] ));
 sky130_fd_sc_hd__dfrtp_4 _20617_ (.CLK(clknet_leaf_24_io_wbs_clk),
    .D(_00915_),
    .RESET_B(_00261_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.y[11] ));
 sky130_fd_sc_hd__dfrtp_4 _20618_ (.CLK(clknet_leaf_24_io_wbs_clk),
    .D(_00916_),
    .RESET_B(_00262_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.y[12] ));
 sky130_fd_sc_hd__dfrtp_4 _20619_ (.CLK(clknet_leaf_24_io_wbs_clk),
    .D(_00917_),
    .RESET_B(_00263_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.y[13] ));
 sky130_fd_sc_hd__dfrtp_4 _20620_ (.CLK(clknet_leaf_24_io_wbs_clk),
    .D(_00918_),
    .RESET_B(_00264_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.y[14] ));
 sky130_fd_sc_hd__dfrtp_4 _20621_ (.CLK(clknet_leaf_24_io_wbs_clk),
    .D(_00919_),
    .RESET_B(_00265_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.y[15] ));
 sky130_fd_sc_hd__dfrtp_4 _20622_ (.CLK(clknet_leaf_24_io_wbs_clk),
    .D(_00920_),
    .RESET_B(_00266_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.y[16] ));
 sky130_fd_sc_hd__dfrtp_1 _20623_ (.CLK(clknet_leaf_10_io_wbs_clk),
    .D(_00921_),
    .RESET_B(_00267_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.z[0] ));
 sky130_fd_sc_hd__dfrtp_1 _20624_ (.CLK(clknet_leaf_10_io_wbs_clk),
    .D(_00922_),
    .RESET_B(_00268_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.z[1] ));
 sky130_fd_sc_hd__dfrtp_1 _20625_ (.CLK(clknet_leaf_3_io_wbs_clk),
    .D(_00923_),
    .RESET_B(_00269_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.z[2] ));
 sky130_fd_sc_hd__dfrtp_1 _20626_ (.CLK(clknet_leaf_3_io_wbs_clk),
    .D(_00924_),
    .RESET_B(_00270_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.z[3] ));
 sky130_fd_sc_hd__dfrtp_1 _20627_ (.CLK(clknet_leaf_3_io_wbs_clk),
    .D(_00925_),
    .RESET_B(_00271_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.z[4] ));
 sky130_fd_sc_hd__dfrtp_1 _20628_ (.CLK(clknet_leaf_3_io_wbs_clk),
    .D(_00926_),
    .RESET_B(_00272_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.z[5] ));
 sky130_fd_sc_hd__dfrtp_1 _20629_ (.CLK(clknet_leaf_3_io_wbs_clk),
    .D(_00927_),
    .RESET_B(_00273_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.z[6] ));
 sky130_fd_sc_hd__dfrtp_1 _20630_ (.CLK(clknet_leaf_4_io_wbs_clk),
    .D(_00928_),
    .RESET_B(_00274_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.z[7] ));
 sky130_fd_sc_hd__dfrtp_1 _20631_ (.CLK(clknet_leaf_4_io_wbs_clk),
    .D(_00929_),
    .RESET_B(_00275_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.z[8] ));
 sky130_fd_sc_hd__dfrtp_1 _20632_ (.CLK(clknet_leaf_5_io_wbs_clk),
    .D(_00930_),
    .RESET_B(_00276_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.z[9] ));
 sky130_fd_sc_hd__dfrtp_1 _20633_ (.CLK(clknet_leaf_5_io_wbs_clk),
    .D(_00931_),
    .RESET_B(_00277_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.z[10] ));
 sky130_fd_sc_hd__dfrtp_1 _20634_ (.CLK(clknet_leaf_5_io_wbs_clk),
    .D(_00932_),
    .RESET_B(_00278_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.z[11] ));
 sky130_fd_sc_hd__dfrtp_1 _20635_ (.CLK(clknet_leaf_5_io_wbs_clk),
    .D(_00933_),
    .RESET_B(_00279_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.z[12] ));
 sky130_fd_sc_hd__dfrtp_1 _20636_ (.CLK(clknet_leaf_5_io_wbs_clk),
    .D(_00934_),
    .RESET_B(_00280_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.z[13] ));
 sky130_fd_sc_hd__dfrtp_1 _20637_ (.CLK(clknet_leaf_6_io_wbs_clk),
    .D(_00935_),
    .RESET_B(_00281_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.z[14] ));
 sky130_fd_sc_hd__dfrtp_1 _20638_ (.CLK(clknet_leaf_6_io_wbs_clk),
    .D(_00936_),
    .RESET_B(_00282_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.z[15] ));
 sky130_fd_sc_hd__dfrtp_4 _20639_ (.CLK(clknet_leaf_6_io_wbs_clk),
    .D(_00937_),
    .RESET_B(_00283_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.z[16] ));
 sky130_fd_sc_hd__dfrtp_4 _20640_ (.CLK(clknet_leaf_10_io_wbs_clk),
    .D(_00938_),
    .RESET_B(_00284_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.quadrant[0] ));
 sky130_fd_sc_hd__dfrtp_4 _20641_ (.CLK(clknet_leaf_10_io_wbs_clk),
    .D(_00939_),
    .RESET_B(_00285_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.quadrant[1] ));
 sky130_fd_sc_hd__dfrtp_4 _20642_ (.CLK(clknet_leaf_7_io_wbs_clk),
    .D(_00940_),
    .RESET_B(_00286_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.iteration[0] ));
 sky130_fd_sc_hd__dfrtp_1 _20643_ (.CLK(clknet_leaf_7_io_wbs_clk),
    .D(_00941_),
    .RESET_B(_00287_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.iteration[1] ));
 sky130_fd_sc_hd__dfrtp_4 _20644_ (.CLK(clknet_leaf_7_io_wbs_clk),
    .D(_00942_),
    .RESET_B(_00288_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.iteration[2] ));
 sky130_fd_sc_hd__dfrtp_4 _20645_ (.CLK(clknet_leaf_6_io_wbs_clk),
    .D(_00943_),
    .RESET_B(_00289_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.iteration[3] ));
 sky130_fd_sc_hd__dfrtp_1 _20646_ (.CLK(clknet_leaf_23_io_wbs_clk),
    .D(_00023_),
    .RESET_B(_00290_),
    .Q(\wfg_interconnect_top.stimulus_0[32] ));
 sky130_fd_sc_hd__dfrtp_1 _20647_ (.CLK(clknet_leaf_83_io_wbs_clk),
    .D(_00944_),
    .RESET_B(_00291_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.temp[14] ));
 sky130_fd_sc_hd__dfrtp_1 _20648_ (.CLK(clknet_leaf_83_io_wbs_clk),
    .D(_00945_),
    .RESET_B(_00292_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.temp[15] ));
 sky130_fd_sc_hd__dfrtp_1 _20649_ (.CLK(clknet_leaf_85_io_wbs_clk),
    .D(_00946_),
    .RESET_B(_00293_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.temp[16] ));
 sky130_fd_sc_hd__dfrtp_1 _20650_ (.CLK(clknet_leaf_85_io_wbs_clk),
    .D(_00947_),
    .RESET_B(_00294_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.temp[17] ));
 sky130_fd_sc_hd__dfrtp_1 _20651_ (.CLK(clknet_leaf_85_io_wbs_clk),
    .D(_00948_),
    .RESET_B(_00295_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.temp[18] ));
 sky130_fd_sc_hd__dfrtp_1 _20652_ (.CLK(clknet_leaf_77_io_wbs_clk),
    .D(_00949_),
    .RESET_B(_00296_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.temp[19] ));
 sky130_fd_sc_hd__dfrtp_1 _20653_ (.CLK(clknet_leaf_77_io_wbs_clk),
    .D(_00950_),
    .RESET_B(_00297_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.temp[20] ));
 sky130_fd_sc_hd__dfrtp_1 _20654_ (.CLK(clknet_leaf_75_io_wbs_clk),
    .D(_00951_),
    .RESET_B(_00298_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.temp[21] ));
 sky130_fd_sc_hd__dfrtp_1 _20655_ (.CLK(clknet_leaf_75_io_wbs_clk),
    .D(_00952_),
    .RESET_B(_00299_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.temp[22] ));
 sky130_fd_sc_hd__dfrtp_1 _20656_ (.CLK(clknet_leaf_75_io_wbs_clk),
    .D(_00953_),
    .RESET_B(_00300_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.temp[23] ));
 sky130_fd_sc_hd__dfrtp_1 _20657_ (.CLK(clknet_leaf_76_io_wbs_clk),
    .D(_00954_),
    .RESET_B(_00301_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.temp[24] ));
 sky130_fd_sc_hd__dfrtp_1 _20658_ (.CLK(clknet_leaf_72_io_wbs_clk),
    .D(_00955_),
    .RESET_B(_00302_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.temp[25] ));
 sky130_fd_sc_hd__dfrtp_1 _20659_ (.CLK(clknet_leaf_76_io_wbs_clk),
    .D(_00956_),
    .RESET_B(_00303_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.temp[26] ));
 sky130_fd_sc_hd__dfrtp_1 _20660_ (.CLK(clknet_leaf_76_io_wbs_clk),
    .D(_00957_),
    .RESET_B(_00304_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.temp[27] ));
 sky130_fd_sc_hd__dfrtp_1 _20661_ (.CLK(clknet_leaf_75_io_wbs_clk),
    .D(_00958_),
    .RESET_B(_00305_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.temp[28] ));
 sky130_fd_sc_hd__dfrtp_1 _20662_ (.CLK(clknet_leaf_76_io_wbs_clk),
    .D(_00959_),
    .RESET_B(_00306_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.temp[29] ));
 sky130_fd_sc_hd__dfrtp_1 _20663_ (.CLK(clknet_leaf_74_io_wbs_clk),
    .D(_00960_),
    .RESET_B(_00307_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.temp[30] ));
 sky130_fd_sc_hd__dfrtp_1 _20664_ (.CLK(clknet_leaf_76_io_wbs_clk),
    .D(_00961_),
    .RESET_B(_00308_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.temp[31] ));
 sky130_fd_sc_hd__dfrtp_1 _20665_ (.CLK(clknet_leaf_10_io_wbs_clk),
    .D(_00962_),
    .RESET_B(_00309_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.phase_in[0] ));
 sky130_fd_sc_hd__dfrtp_1 _20666_ (.CLK(clknet_leaf_10_io_wbs_clk),
    .D(_00963_),
    .RESET_B(_00310_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.phase_in[1] ));
 sky130_fd_sc_hd__dfrtp_1 _20667_ (.CLK(clknet_leaf_3_io_wbs_clk),
    .D(_00964_),
    .RESET_B(_00311_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.phase_in[2] ));
 sky130_fd_sc_hd__dfrtp_1 _20668_ (.CLK(clknet_leaf_3_io_wbs_clk),
    .D(_00965_),
    .RESET_B(_00312_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.phase_in[3] ));
 sky130_fd_sc_hd__dfrtp_1 _20669_ (.CLK(clknet_leaf_3_io_wbs_clk),
    .D(_00966_),
    .RESET_B(_00313_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.phase_in[4] ));
 sky130_fd_sc_hd__dfrtp_1 _20670_ (.CLK(clknet_leaf_2_io_wbs_clk),
    .D(_00967_),
    .RESET_B(_00314_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.phase_in[5] ));
 sky130_fd_sc_hd__dfrtp_1 _20671_ (.CLK(clknet_leaf_4_io_wbs_clk),
    .D(_00968_),
    .RESET_B(_00315_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.phase_in[6] ));
 sky130_fd_sc_hd__dfrtp_1 _20672_ (.CLK(clknet_leaf_4_io_wbs_clk),
    .D(_00969_),
    .RESET_B(_00316_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.phase_in[7] ));
 sky130_fd_sc_hd__dfrtp_1 _20673_ (.CLK(clknet_leaf_0_io_wbs_clk),
    .D(_00970_),
    .RESET_B(_00317_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.phase_in[8] ));
 sky130_fd_sc_hd__dfrtp_1 _20674_ (.CLK(clknet_leaf_0_io_wbs_clk),
    .D(_00971_),
    .RESET_B(_00318_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.phase_in[9] ));
 sky130_fd_sc_hd__dfrtp_1 _20675_ (.CLK(clknet_leaf_4_io_wbs_clk),
    .D(_00972_),
    .RESET_B(_00319_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.phase_in[10] ));
 sky130_fd_sc_hd__dfrtp_1 _20676_ (.CLK(clknet_leaf_4_io_wbs_clk),
    .D(_00973_),
    .RESET_B(_00320_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.phase_in[11] ));
 sky130_fd_sc_hd__dfrtp_1 _20677_ (.CLK(clknet_leaf_0_io_wbs_clk),
    .D(_00974_),
    .RESET_B(_00321_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.phase_in[12] ));
 sky130_fd_sc_hd__dfrtp_1 _20678_ (.CLK(clknet_leaf_5_io_wbs_clk),
    .D(_00975_),
    .RESET_B(_00322_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.phase_in[13] ));
 sky130_fd_sc_hd__dfrtp_1 _20679_ (.CLK(clknet_leaf_2_io_wbs_clk),
    .D(_00976_),
    .RESET_B(_00323_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.phase_in[14] ));
 sky130_fd_sc_hd__dfrtp_1 _20680_ (.CLK(clknet_leaf_10_io_wbs_clk),
    .D(_00977_),
    .RESET_B(_00324_),
    .Q(\wfg_stim_sine_top.wfg_stim_sine.phase_in[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20681_ (.CLK(clknet_leaf_92_io_wbs_clk),
    .D(_00978_),
    .Q(\wfg_stim_mem_top.wbs_dat_o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20682_ (.CLK(clknet_leaf_1_io_wbs_clk),
    .D(_00979_),
    .Q(\wfg_stim_mem_top.wbs_dat_o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20683_ (.CLK(clknet_leaf_1_io_wbs_clk),
    .D(_00980_),
    .Q(\wfg_stim_mem_top.wbs_dat_o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20684_ (.CLK(clknet_leaf_2_io_wbs_clk),
    .D(_00981_),
    .Q(\wfg_stim_mem_top.wbs_dat_o[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20685_ (.CLK(clknet_leaf_1_io_wbs_clk),
    .D(_00982_),
    .Q(\wfg_stim_mem_top.wbs_dat_o[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20686_ (.CLK(clknet_leaf_2_io_wbs_clk),
    .D(_00983_),
    .Q(\wfg_stim_mem_top.wbs_dat_o[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20687_ (.CLK(clknet_leaf_2_io_wbs_clk),
    .D(_00984_),
    .Q(\wfg_stim_mem_top.wbs_dat_o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20688_ (.CLK(clknet_leaf_1_io_wbs_clk),
    .D(_00985_),
    .Q(\wfg_stim_mem_top.wbs_dat_o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20689_ (.CLK(clknet_leaf_2_io_wbs_clk),
    .D(_00986_),
    .Q(\wfg_stim_mem_top.wbs_dat_o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20690_ (.CLK(clknet_leaf_2_io_wbs_clk),
    .D(_00987_),
    .Q(\wfg_stim_mem_top.wbs_dat_o[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20691_ (.CLK(clknet_leaf_2_io_wbs_clk),
    .D(_00988_),
    .Q(\wfg_stim_mem_top.wbs_dat_o[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20692_ (.CLK(clknet_leaf_102_io_wbs_clk),
    .D(_00989_),
    .Q(\wfg_stim_mem_top.wbs_dat_o[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20693_ (.CLK(clknet_leaf_102_io_wbs_clk),
    .D(_00990_),
    .Q(\wfg_stim_mem_top.wbs_dat_o[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20694_ (.CLK(clknet_leaf_102_io_wbs_clk),
    .D(_00991_),
    .Q(\wfg_stim_mem_top.wbs_dat_o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20695_ (.CLK(clknet_leaf_102_io_wbs_clk),
    .D(_00992_),
    .Q(\wfg_stim_mem_top.wbs_dat_o[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20696_ (.CLK(clknet_leaf_102_io_wbs_clk),
    .D(_00993_),
    .Q(\wfg_stim_mem_top.wbs_dat_o[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20697_ (.CLK(clknet_leaf_94_io_wbs_clk),
    .D(_00994_),
    .Q(\wfg_stim_mem_top.wbs_dat_o[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20698_ (.CLK(clknet_leaf_92_io_wbs_clk),
    .D(_00995_),
    .Q(\wfg_stim_mem_top.wbs_dat_o[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20699_ (.CLK(clknet_leaf_94_io_wbs_clk),
    .D(_00996_),
    .Q(\wfg_stim_mem_top.wbs_dat_o[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20700_ (.CLK(clknet_leaf_94_io_wbs_clk),
    .D(_00997_),
    .Q(\wfg_stim_mem_top.wbs_dat_o[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20701_ (.CLK(clknet_leaf_94_io_wbs_clk),
    .D(_00998_),
    .Q(\wfg_stim_mem_top.wbs_dat_o[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20702_ (.CLK(clknet_leaf_81_io_wbs_clk),
    .D(_00999_),
    .Q(\wfg_stim_mem_top.wbs_dat_o[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20703_ (.CLK(clknet_leaf_80_io_wbs_clk),
    .D(_01000_),
    .Q(\wfg_stim_mem_top.wbs_dat_o[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20704_ (.CLK(clknet_leaf_81_io_wbs_clk),
    .D(_01001_),
    .Q(\wfg_stim_mem_top.wbs_dat_o[23] ));
 sky130_fd_sc_hd__dfxtp_2 _20705_ (.CLK(clknet_leaf_11_io_wbs_clk),
    .D(_01002_),
    .Q(\wfg_stim_sine_top.ctrl_en_q ));
 sky130_fd_sc_hd__dfxtp_2 _20706_ (.CLK(clknet_leaf_83_io_wbs_clk),
    .D(_01003_),
    .Q(\wfg_stim_sine_top.gain_val_q[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20707_ (.CLK(clknet_leaf_82_io_wbs_clk),
    .D(_01004_),
    .Q(\wfg_stim_sine_top.gain_val_q[1] ));
 sky130_fd_sc_hd__dfxtp_4 _20708_ (.CLK(clknet_leaf_80_io_wbs_clk),
    .D(_01005_),
    .Q(\wfg_stim_sine_top.gain_val_q[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20709_ (.CLK(clknet_leaf_78_io_wbs_clk),
    .D(_01006_),
    .Q(\wfg_stim_sine_top.gain_val_q[3] ));
 sky130_fd_sc_hd__dfxtp_4 _20710_ (.CLK(clknet_leaf_80_io_wbs_clk),
    .D(_01007_),
    .Q(\wfg_stim_sine_top.gain_val_q[4] ));
 sky130_fd_sc_hd__dfxtp_4 _20711_ (.CLK(clknet_leaf_80_io_wbs_clk),
    .D(_01008_),
    .Q(\wfg_stim_sine_top.gain_val_q[5] ));
 sky130_fd_sc_hd__dfxtp_2 _20712_ (.CLK(clknet_leaf_80_io_wbs_clk),
    .D(_01009_),
    .Q(\wfg_stim_sine_top.gain_val_q[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20713_ (.CLK(clknet_leaf_82_io_wbs_clk),
    .D(_01010_),
    .Q(\wfg_stim_sine_top.gain_val_q[7] ));
 sky130_fd_sc_hd__dfxtp_2 _20714_ (.CLK(clknet_leaf_82_io_wbs_clk),
    .D(_01011_),
    .Q(\wfg_stim_sine_top.gain_val_q[8] ));
 sky130_fd_sc_hd__dfxtp_2 _20715_ (.CLK(clknet_leaf_82_io_wbs_clk),
    .D(_01012_),
    .Q(\wfg_stim_sine_top.gain_val_q[9] ));
 sky130_fd_sc_hd__dfxtp_2 _20716_ (.CLK(clknet_leaf_82_io_wbs_clk),
    .D(_01013_),
    .Q(\wfg_stim_sine_top.gain_val_q[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20717_ (.CLK(clknet_leaf_82_io_wbs_clk),
    .D(_01014_),
    .Q(\wfg_stim_sine_top.gain_val_q[11] ));
 sky130_fd_sc_hd__dfxtp_2 _20718_ (.CLK(clknet_leaf_82_io_wbs_clk),
    .D(_01015_),
    .Q(\wfg_stim_sine_top.gain_val_q[12] ));
 sky130_fd_sc_hd__dfxtp_2 _20719_ (.CLK(clknet_leaf_83_io_wbs_clk),
    .D(_01016_),
    .Q(\wfg_stim_sine_top.gain_val_q[13] ));
 sky130_fd_sc_hd__dfxtp_2 _20720_ (.CLK(clknet_leaf_83_io_wbs_clk),
    .D(_01017_),
    .Q(\wfg_stim_sine_top.gain_val_q[14] ));
 sky130_fd_sc_hd__dfxtp_2 _20721_ (.CLK(clknet_leaf_83_io_wbs_clk),
    .D(_01018_),
    .Q(\wfg_stim_sine_top.gain_val_q[15] ));
 sky130_fd_sc_hd__dfxtp_2 _20722_ (.CLK(clknet_leaf_89_io_wbs_clk),
    .D(_01019_),
    .Q(\wfg_stim_sine_top.inc_val_q[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20723_ (.CLK(clknet_leaf_84_io_wbs_clk),
    .D(_01020_),
    .Q(\wfg_stim_sine_top.inc_val_q[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20724_ (.CLK(clknet_leaf_84_io_wbs_clk),
    .D(_01021_),
    .Q(\wfg_stim_sine_top.inc_val_q[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20725_ (.CLK(clknet_leaf_84_io_wbs_clk),
    .D(_01022_),
    .Q(\wfg_stim_sine_top.inc_val_q[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20726_ (.CLK(clknet_leaf_83_io_wbs_clk),
    .D(_01023_),
    .Q(\wfg_stim_sine_top.inc_val_q[4] ));
 sky130_fd_sc_hd__dfxtp_2 _20727_ (.CLK(clknet_leaf_82_io_wbs_clk),
    .D(_01024_),
    .Q(\wfg_stim_sine_top.inc_val_q[5] ));
 sky130_fd_sc_hd__dfxtp_2 _20728_ (.CLK(clknet_leaf_81_io_wbs_clk),
    .D(_01025_),
    .Q(\wfg_stim_sine_top.inc_val_q[6] ));
 sky130_fd_sc_hd__dfxtp_2 _20729_ (.CLK(clknet_leaf_82_io_wbs_clk),
    .D(_01026_),
    .Q(\wfg_stim_sine_top.inc_val_q[7] ));
 sky130_fd_sc_hd__dfxtp_2 _20730_ (.CLK(clknet_leaf_93_io_wbs_clk),
    .D(_01027_),
    .Q(\wfg_stim_sine_top.inc_val_q[8] ));
 sky130_fd_sc_hd__dfxtp_2 _20731_ (.CLK(clknet_leaf_82_io_wbs_clk),
    .D(_01028_),
    .Q(\wfg_stim_sine_top.inc_val_q[9] ));
 sky130_fd_sc_hd__dfxtp_2 _20732_ (.CLK(clknet_leaf_89_io_wbs_clk),
    .D(_01029_),
    .Q(\wfg_stim_sine_top.inc_val_q[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20733_ (.CLK(clknet_leaf_93_io_wbs_clk),
    .D(_01030_),
    .Q(\wfg_stim_sine_top.inc_val_q[11] ));
 sky130_fd_sc_hd__dfxtp_2 _20734_ (.CLK(clknet_leaf_2_io_wbs_clk),
    .D(_01031_),
    .Q(\wfg_stim_sine_top.inc_val_q[12] ));
 sky130_fd_sc_hd__dfxtp_4 _20735_ (.CLK(clknet_leaf_89_io_wbs_clk),
    .D(_01032_),
    .Q(\wfg_stim_sine_top.inc_val_q[13] ));
 sky130_fd_sc_hd__dfxtp_2 _20736_ (.CLK(clknet_leaf_89_io_wbs_clk),
    .D(_01033_),
    .Q(\wfg_stim_sine_top.inc_val_q[14] ));
 sky130_fd_sc_hd__dfxtp_2 _20737_ (.CLK(clknet_leaf_89_io_wbs_clk),
    .D(_01034_),
    .Q(\wfg_stim_sine_top.inc_val_q[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20738_ (.CLK(clknet_leaf_84_io_wbs_clk),
    .D(_01035_),
    .Q(\wfg_stim_sine_top.offset_val_q[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20739_ (.CLK(clknet_leaf_84_io_wbs_clk),
    .D(_01036_),
    .Q(\wfg_stim_sine_top.offset_val_q[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20740_ (.CLK(clknet_leaf_80_io_wbs_clk),
    .D(_01037_),
    .Q(\wfg_stim_sine_top.offset_val_q[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20741_ (.CLK(clknet_leaf_80_io_wbs_clk),
    .D(_01038_),
    .Q(\wfg_stim_sine_top.offset_val_q[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20742_ (.CLK(clknet_leaf_80_io_wbs_clk),
    .D(_01039_),
    .Q(\wfg_stim_sine_top.offset_val_q[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20743_ (.CLK(clknet_leaf_80_io_wbs_clk),
    .D(_01040_),
    .Q(\wfg_stim_sine_top.offset_val_q[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20744_ (.CLK(clknet_leaf_83_io_wbs_clk),
    .D(_01041_),
    .Q(\wfg_stim_sine_top.offset_val_q[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20745_ (.CLK(clknet_leaf_83_io_wbs_clk),
    .D(_01042_),
    .Q(\wfg_stim_sine_top.offset_val_q[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20746_ (.CLK(clknet_leaf_83_io_wbs_clk),
    .D(_01043_),
    .Q(\wfg_stim_sine_top.offset_val_q[8] ));
 sky130_fd_sc_hd__dfxtp_2 _20747_ (.CLK(clknet_leaf_83_io_wbs_clk),
    .D(_01044_),
    .Q(\wfg_stim_sine_top.offset_val_q[9] ));
 sky130_fd_sc_hd__dfxtp_2 _20748_ (.CLK(clknet_leaf_84_io_wbs_clk),
    .D(_01045_),
    .Q(\wfg_stim_sine_top.offset_val_q[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20749_ (.CLK(clknet_leaf_86_io_wbs_clk),
    .D(_01046_),
    .Q(\wfg_stim_sine_top.offset_val_q[11] ));
 sky130_fd_sc_hd__dfxtp_2 _20750_ (.CLK(clknet_leaf_85_io_wbs_clk),
    .D(_01047_),
    .Q(\wfg_stim_sine_top.offset_val_q[12] ));
 sky130_fd_sc_hd__dfxtp_2 _20751_ (.CLK(clknet_leaf_85_io_wbs_clk),
    .D(_01048_),
    .Q(\wfg_stim_sine_top.offset_val_q[13] ));
 sky130_fd_sc_hd__dfxtp_2 _20752_ (.CLK(clknet_leaf_86_io_wbs_clk),
    .D(_01049_),
    .Q(\wfg_stim_sine_top.offset_val_q[14] ));
 sky130_fd_sc_hd__dfxtp_2 _20753_ (.CLK(clknet_leaf_86_io_wbs_clk),
    .D(_01050_),
    .Q(\wfg_stim_sine_top.offset_val_q[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20754_ (.CLK(clknet_leaf_84_io_wbs_clk),
    .D(_01051_),
    .Q(\wfg_stim_sine_top.offset_val_q[16] ));
 sky130_fd_sc_hd__dfxtp_2 _20755_ (.CLK(clknet_leaf_84_io_wbs_clk),
    .D(_01052_),
    .Q(\wfg_stim_sine_top.offset_val_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _20756_ (.CLK(clknet_leaf_23_io_wbs_clk),
    .D(\wfg_stim_mem_top.wfg_stim_mem.cur_state[3] ),
    .RESET_B(_00325_),
    .Q(\wfg_interconnect_top.stimulus_1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _20757_ (.CLK(clknet_leaf_101_io_wbs_clk),
    .D(_01053_),
    .Q(\wfg_interconnect_top.wbs_ack_o ));
 sky130_fd_sc_hd__dfrtp_1 _20758_ (.CLK(clknet_leaf_107_io_wbs_clk),
    .D(_01054_),
    .RESET_B(_00326_),
    .Q(net101));
 sky130_fd_sc_hd__dfrtp_1 _20759_ (.CLK(clknet_leaf_108_io_wbs_clk),
    .D(_01055_),
    .RESET_B(_00327_),
    .Q(net102));
 sky130_fd_sc_hd__dfrtp_1 _20760_ (.CLK(clknet_leaf_108_io_wbs_clk),
    .D(_01056_),
    .RESET_B(_00328_),
    .Q(net103));
 sky130_fd_sc_hd__dfrtp_2 _20761_ (.CLK(clknet_leaf_108_io_wbs_clk),
    .D(_01057_),
    .RESET_B(_00329_),
    .Q(net104));
 sky130_fd_sc_hd__dfrtp_1 _20762_ (.CLK(clknet_leaf_109_io_wbs_clk),
    .D(_01058_),
    .RESET_B(_00330_),
    .Q(net105));
 sky130_fd_sc_hd__dfrtp_1 _20763_ (.CLK(clknet_leaf_109_io_wbs_clk),
    .D(_01059_),
    .RESET_B(_00331_),
    .Q(net106));
 sky130_fd_sc_hd__dfrtp_1 _20764_ (.CLK(clknet_leaf_0_io_wbs_clk),
    .D(_01060_),
    .RESET_B(_00332_),
    .Q(net107));
 sky130_fd_sc_hd__dfrtp_1 _20765_ (.CLK(clknet_leaf_0_io_wbs_clk),
    .D(_01061_),
    .RESET_B(_00333_),
    .Q(net108));
 sky130_fd_sc_hd__dfrtp_1 _20766_ (.CLK(clknet_leaf_0_io_wbs_clk),
    .D(_01062_),
    .RESET_B(_00334_),
    .Q(net109));
 sky130_fd_sc_hd__dfrtp_2 _20767_ (.CLK(clknet_leaf_1_io_wbs_clk),
    .D(_01063_),
    .RESET_B(_00335_),
    .Q(net110));
 sky130_fd_sc_hd__dfrtp_1 _20768_ (.CLK(clknet_leaf_103_io_wbs_clk),
    .D(_01064_),
    .RESET_B(_00336_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.cur_address[10] ));
 sky130_fd_sc_hd__dfrtp_1 _20769_ (.CLK(clknet_leaf_106_io_wbs_clk),
    .D(_01065_),
    .RESET_B(_00337_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.cur_address[11] ));
 sky130_fd_sc_hd__dfrtp_1 _20770_ (.CLK(clknet_leaf_105_io_wbs_clk),
    .D(_01066_),
    .RESET_B(_00338_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.cur_address[12] ));
 sky130_fd_sc_hd__dfrtp_1 _20771_ (.CLK(clknet_leaf_104_io_wbs_clk),
    .D(_01067_),
    .RESET_B(_00339_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.cur_address[13] ));
 sky130_fd_sc_hd__dfrtp_1 _20772_ (.CLK(clknet_leaf_103_io_wbs_clk),
    .D(_01068_),
    .RESET_B(_00340_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.cur_address[14] ));
 sky130_fd_sc_hd__dfrtp_1 _20773_ (.CLK(clknet_leaf_103_io_wbs_clk),
    .D(_01069_),
    .RESET_B(_00341_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.cur_address[15] ));
 sky130_fd_sc_hd__dfrtp_1 _20774_ (.CLK(clknet_leaf_49_io_wbs_clk),
    .D(_01070_),
    .RESET_B(_00342_),
    .Q(\wfg_interconnect_top.stimulus_1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _20775_ (.CLK(clknet_leaf_49_io_wbs_clk),
    .D(_01071_),
    .RESET_B(_00343_),
    .Q(\wfg_interconnect_top.stimulus_1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _20776_ (.CLK(clknet_leaf_51_io_wbs_clk),
    .D(_01072_),
    .RESET_B(_00344_),
    .Q(\wfg_interconnect_top.stimulus_1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _20777_ (.CLK(clknet_leaf_49_io_wbs_clk),
    .D(_01073_),
    .RESET_B(_00345_),
    .Q(\wfg_interconnect_top.stimulus_1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _20778_ (.CLK(clknet_leaf_51_io_wbs_clk),
    .D(_01074_),
    .RESET_B(_00346_),
    .Q(\wfg_interconnect_top.stimulus_1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _20779_ (.CLK(clknet_leaf_51_io_wbs_clk),
    .D(_01075_),
    .RESET_B(_00347_),
    .Q(\wfg_interconnect_top.stimulus_1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _20780_ (.CLK(clknet_leaf_51_io_wbs_clk),
    .D(_01076_),
    .RESET_B(_00348_),
    .Q(\wfg_interconnect_top.stimulus_1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _20781_ (.CLK(clknet_leaf_51_io_wbs_clk),
    .D(_01077_),
    .RESET_B(_00349_),
    .Q(\wfg_interconnect_top.stimulus_1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _20782_ (.CLK(clknet_leaf_50_io_wbs_clk),
    .D(_01078_),
    .RESET_B(_00350_),
    .Q(\wfg_interconnect_top.stimulus_1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _20783_ (.CLK(clknet_leaf_50_io_wbs_clk),
    .D(_01079_),
    .RESET_B(_00351_),
    .Q(\wfg_interconnect_top.stimulus_1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _20784_ (.CLK(clknet_leaf_50_io_wbs_clk),
    .D(_01080_),
    .RESET_B(_00352_),
    .Q(\wfg_interconnect_top.stimulus_1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _20785_ (.CLK(clknet_leaf_54_io_wbs_clk),
    .D(_01081_),
    .RESET_B(_00353_),
    .Q(\wfg_interconnect_top.stimulus_1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _20786_ (.CLK(clknet_leaf_55_io_wbs_clk),
    .D(_01082_),
    .RESET_B(_00354_),
    .Q(\wfg_interconnect_top.stimulus_1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _20787_ (.CLK(clknet_leaf_54_io_wbs_clk),
    .D(_01083_),
    .RESET_B(_00355_),
    .Q(\wfg_interconnect_top.stimulus_1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _20788_ (.CLK(clknet_leaf_53_io_wbs_clk),
    .D(_01084_),
    .RESET_B(_00356_),
    .Q(\wfg_interconnect_top.stimulus_1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _20789_ (.CLK(clknet_leaf_53_io_wbs_clk),
    .D(_01085_),
    .RESET_B(_00357_),
    .Q(\wfg_interconnect_top.stimulus_1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _20790_ (.CLK(clknet_leaf_53_io_wbs_clk),
    .D(_01086_),
    .RESET_B(_00358_),
    .Q(\wfg_interconnect_top.stimulus_1[16] ));
 sky130_fd_sc_hd__dfrtp_1 _20791_ (.CLK(clknet_leaf_53_io_wbs_clk),
    .D(_01087_),
    .RESET_B(_00359_),
    .Q(\wfg_interconnect_top.stimulus_1[17] ));
 sky130_fd_sc_hd__dfrtp_1 _20792_ (.CLK(clknet_leaf_53_io_wbs_clk),
    .D(_01088_),
    .RESET_B(_00360_),
    .Q(\wfg_interconnect_top.stimulus_1[18] ));
 sky130_fd_sc_hd__dfrtp_1 _20793_ (.CLK(clknet_leaf_56_io_wbs_clk),
    .D(_01089_),
    .RESET_B(_00361_),
    .Q(\wfg_interconnect_top.stimulus_1[19] ));
 sky130_fd_sc_hd__dfrtp_1 _20794_ (.CLK(clknet_leaf_56_io_wbs_clk),
    .D(_01090_),
    .RESET_B(_00362_),
    .Q(\wfg_interconnect_top.stimulus_1[20] ));
 sky130_fd_sc_hd__dfrtp_1 _20795_ (.CLK(clknet_leaf_56_io_wbs_clk),
    .D(_01091_),
    .RESET_B(_00363_),
    .Q(\wfg_interconnect_top.stimulus_1[21] ));
 sky130_fd_sc_hd__dfrtp_1 _20796_ (.CLK(clknet_leaf_56_io_wbs_clk),
    .D(_01092_),
    .RESET_B(_00364_),
    .Q(\wfg_interconnect_top.stimulus_1[22] ));
 sky130_fd_sc_hd__dfrtp_1 _20797_ (.CLK(clknet_leaf_57_io_wbs_clk),
    .D(_01093_),
    .RESET_B(_00365_),
    .Q(\wfg_interconnect_top.stimulus_1[23] ));
 sky130_fd_sc_hd__dfrtp_1 _20798_ (.CLK(clknet_leaf_57_io_wbs_clk),
    .D(_01094_),
    .RESET_B(_00366_),
    .Q(\wfg_interconnect_top.stimulus_1[24] ));
 sky130_fd_sc_hd__dfrtp_1 _20799_ (.CLK(clknet_leaf_57_io_wbs_clk),
    .D(_01095_),
    .RESET_B(_00367_),
    .Q(\wfg_interconnect_top.stimulus_1[25] ));
 sky130_fd_sc_hd__dfrtp_1 _20800_ (.CLK(clknet_leaf_57_io_wbs_clk),
    .D(_01096_),
    .RESET_B(_00368_),
    .Q(\wfg_interconnect_top.stimulus_1[26] ));
 sky130_fd_sc_hd__dfrtp_1 _20801_ (.CLK(clknet_leaf_57_io_wbs_clk),
    .D(_01097_),
    .RESET_B(_00369_),
    .Q(\wfg_interconnect_top.stimulus_1[27] ));
 sky130_fd_sc_hd__dfrtp_1 _20802_ (.CLK(clknet_leaf_57_io_wbs_clk),
    .D(_01098_),
    .RESET_B(_00370_),
    .Q(\wfg_interconnect_top.stimulus_1[28] ));
 sky130_fd_sc_hd__dfrtp_1 _20803_ (.CLK(clknet_leaf_57_io_wbs_clk),
    .D(_01099_),
    .RESET_B(_00371_),
    .Q(\wfg_interconnect_top.stimulus_1[29] ));
 sky130_fd_sc_hd__dfrtp_1 _20804_ (.CLK(clknet_leaf_57_io_wbs_clk),
    .D(_01100_),
    .RESET_B(_00372_),
    .Q(\wfg_interconnect_top.stimulus_1[30] ));
 sky130_fd_sc_hd__dfrtp_1 _20805_ (.CLK(clknet_leaf_56_io_wbs_clk),
    .D(_01101_),
    .RESET_B(_00373_),
    .Q(\wfg_interconnect_top.stimulus_1[31] ));
 sky130_fd_sc_hd__dfrtp_1 _20806_ (.CLK(clknet_leaf_50_io_wbs_clk),
    .D(_01102_),
    .RESET_B(_00374_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[0] ));
 sky130_fd_sc_hd__dfrtp_1 _20807_ (.CLK(clknet_leaf_50_io_wbs_clk),
    .D(_01103_),
    .RESET_B(_00375_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[1] ));
 sky130_fd_sc_hd__dfrtp_1 _20808_ (.CLK(clknet_leaf_50_io_wbs_clk),
    .D(_01104_),
    .RESET_B(_00376_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[2] ));
 sky130_fd_sc_hd__dfrtp_1 _20809_ (.CLK(clknet_leaf_51_io_wbs_clk),
    .D(_01105_),
    .RESET_B(_00377_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[3] ));
 sky130_fd_sc_hd__dfrtp_1 _20810_ (.CLK(clknet_leaf_51_io_wbs_clk),
    .D(_01106_),
    .RESET_B(_00378_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[4] ));
 sky130_fd_sc_hd__dfrtp_1 _20811_ (.CLK(clknet_leaf_50_io_wbs_clk),
    .D(_01107_),
    .RESET_B(_00379_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[5] ));
 sky130_fd_sc_hd__dfrtp_1 _20812_ (.CLK(clknet_leaf_50_io_wbs_clk),
    .D(_01108_),
    .RESET_B(_00380_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[6] ));
 sky130_fd_sc_hd__dfrtp_1 _20813_ (.CLK(clknet_leaf_50_io_wbs_clk),
    .D(_01109_),
    .RESET_B(_00381_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[7] ));
 sky130_fd_sc_hd__dfrtp_1 _20814_ (.CLK(clknet_leaf_54_io_wbs_clk),
    .D(_01110_),
    .RESET_B(_00382_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[8] ));
 sky130_fd_sc_hd__dfrtp_1 _20815_ (.CLK(clknet_leaf_54_io_wbs_clk),
    .D(_01111_),
    .RESET_B(_00383_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[9] ));
 sky130_fd_sc_hd__dfrtp_1 _20816_ (.CLK(clknet_leaf_54_io_wbs_clk),
    .D(_01112_),
    .RESET_B(_00384_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[10] ));
 sky130_fd_sc_hd__dfrtp_1 _20817_ (.CLK(clknet_leaf_55_io_wbs_clk),
    .D(_01113_),
    .RESET_B(_00385_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[11] ));
 sky130_fd_sc_hd__dfrtp_1 _20818_ (.CLK(clknet_leaf_55_io_wbs_clk),
    .D(_01114_),
    .RESET_B(_00386_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[12] ));
 sky130_fd_sc_hd__dfrtp_1 _20819_ (.CLK(clknet_leaf_54_io_wbs_clk),
    .D(_01115_),
    .RESET_B(_00387_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[13] ));
 sky130_fd_sc_hd__dfrtp_1 _20820_ (.CLK(clknet_leaf_53_io_wbs_clk),
    .D(_01116_),
    .RESET_B(_00388_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[14] ));
 sky130_fd_sc_hd__dfrtp_1 _20821_ (.CLK(clknet_leaf_53_io_wbs_clk),
    .D(_01117_),
    .RESET_B(_00389_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[15] ));
 sky130_fd_sc_hd__dfrtp_1 _20822_ (.CLK(clknet_leaf_53_io_wbs_clk),
    .D(_01118_),
    .RESET_B(_00390_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[16] ));
 sky130_fd_sc_hd__dfrtp_1 _20823_ (.CLK(clknet_leaf_53_io_wbs_clk),
    .D(_01119_),
    .RESET_B(_00391_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[17] ));
 sky130_fd_sc_hd__dfrtp_1 _20824_ (.CLK(clknet_leaf_55_io_wbs_clk),
    .D(_01120_),
    .RESET_B(_00392_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[18] ));
 sky130_fd_sc_hd__dfrtp_1 _20825_ (.CLK(clknet_leaf_56_io_wbs_clk),
    .D(_01121_),
    .RESET_B(_00393_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[19] ));
 sky130_fd_sc_hd__dfrtp_1 _20826_ (.CLK(clknet_leaf_55_io_wbs_clk),
    .D(_01122_),
    .RESET_B(_00394_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[20] ));
 sky130_fd_sc_hd__dfrtp_1 _20827_ (.CLK(clknet_leaf_55_io_wbs_clk),
    .D(_01123_),
    .RESET_B(_00395_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[21] ));
 sky130_fd_sc_hd__dfrtp_1 _20828_ (.CLK(clknet_leaf_56_io_wbs_clk),
    .D(_01124_),
    .RESET_B(_00396_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[22] ));
 sky130_fd_sc_hd__dfrtp_1 _20829_ (.CLK(clknet_leaf_55_io_wbs_clk),
    .D(_01125_),
    .RESET_B(_00397_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[23] ));
 sky130_fd_sc_hd__dfrtp_1 _20830_ (.CLK(clknet_leaf_55_io_wbs_clk),
    .D(_01126_),
    .RESET_B(_00398_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[24] ));
 sky130_fd_sc_hd__dfrtp_1 _20831_ (.CLK(clknet_leaf_55_io_wbs_clk),
    .D(_01127_),
    .RESET_B(_00399_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[25] ));
 sky130_fd_sc_hd__dfrtp_1 _20832_ (.CLK(clknet_leaf_55_io_wbs_clk),
    .D(_01128_),
    .RESET_B(_00400_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[26] ));
 sky130_fd_sc_hd__dfrtp_1 _20833_ (.CLK(clknet_leaf_56_io_wbs_clk),
    .D(_01129_),
    .RESET_B(_00401_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[27] ));
 sky130_fd_sc_hd__dfrtp_1 _20834_ (.CLK(clknet_leaf_55_io_wbs_clk),
    .D(_01130_),
    .RESET_B(_00402_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[28] ));
 sky130_fd_sc_hd__dfrtp_1 _20835_ (.CLK(clknet_leaf_55_io_wbs_clk),
    .D(_01131_),
    .RESET_B(_00403_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[29] ));
 sky130_fd_sc_hd__dfrtp_1 _20836_ (.CLK(clknet_leaf_56_io_wbs_clk),
    .D(_01132_),
    .RESET_B(_00404_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[30] ));
 sky130_fd_sc_hd__dfrtp_1 _20837_ (.CLK(clknet_leaf_55_io_wbs_clk),
    .D(_01133_),
    .RESET_B(_00405_),
    .Q(\wfg_stim_mem_top.wfg_stim_mem.data_calc[31] ));
 sky130_fd_sc_hd__dfxtp_1 _20838_ (.CLK(clknet_leaf_92_io_wbs_clk),
    .D(_01134_),
    .Q(\wfg_interconnect_top.wbs_dat_o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20839_ (.CLK(clknet_leaf_91_io_wbs_clk),
    .D(_01135_),
    .Q(\wfg_interconnect_top.wbs_dat_o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20840_ (.CLK(clknet_leaf_102_io_wbs_clk),
    .D(_01136_),
    .Q(\wfg_stim_mem_top.ctrl_en_q ));
 sky130_fd_sc_hd__dfxtp_2 _20841_ (.CLK(clknet_leaf_22_io_wbs_clk),
    .D(_01137_),
    .Q(\wfg_stim_mem_top.cfg_gain_q[8] ));
 sky130_fd_sc_hd__dfxtp_4 _20842_ (.CLK(clknet_leaf_34_io_wbs_clk),
    .D(_01138_),
    .Q(\wfg_stim_mem_top.cfg_gain_q[9] ));
 sky130_fd_sc_hd__dfxtp_2 _20843_ (.CLK(clknet_leaf_29_io_wbs_clk),
    .D(_01139_),
    .Q(\wfg_stim_mem_top.cfg_gain_q[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20844_ (.CLK(clknet_leaf_32_io_wbs_clk),
    .D(_01140_),
    .Q(\wfg_stim_mem_top.cfg_gain_q[11] ));
 sky130_fd_sc_hd__dfxtp_4 _20845_ (.CLK(clknet_3_2_0_io_wbs_clk),
    .D(_01141_),
    .Q(\wfg_stim_mem_top.cfg_gain_q[12] ));
 sky130_fd_sc_hd__dfxtp_4 _20846_ (.CLK(clknet_leaf_34_io_wbs_clk),
    .D(_01142_),
    .Q(\wfg_stim_mem_top.cfg_gain_q[13] ));
 sky130_fd_sc_hd__dfxtp_4 _20847_ (.CLK(clknet_leaf_28_io_wbs_clk),
    .D(_01143_),
    .Q(\wfg_stim_mem_top.cfg_gain_q[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20848_ (.CLK(clknet_leaf_28_io_wbs_clk),
    .D(_01144_),
    .Q(\wfg_stim_mem_top.cfg_gain_q[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20849_ (.CLK(clknet_leaf_28_io_wbs_clk),
    .D(_01145_),
    .Q(\wfg_stim_mem_top.cfg_gain_q[16] ));
 sky130_fd_sc_hd__dfxtp_2 _20850_ (.CLK(clknet_leaf_29_io_wbs_clk),
    .D(_01146_),
    .Q(\wfg_stim_mem_top.cfg_gain_q[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20851_ (.CLK(clknet_leaf_29_io_wbs_clk),
    .D(_01147_),
    .Q(\wfg_stim_mem_top.cfg_gain_q[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20852_ (.CLK(clknet_leaf_29_io_wbs_clk),
    .D(_01148_),
    .Q(\wfg_stim_mem_top.cfg_gain_q[19] ));
 sky130_fd_sc_hd__dfxtp_4 _20853_ (.CLK(clknet_leaf_29_io_wbs_clk),
    .D(_01149_),
    .Q(\wfg_stim_mem_top.cfg_gain_q[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20854_ (.CLK(clknet_leaf_29_io_wbs_clk),
    .D(_01150_),
    .Q(\wfg_stim_mem_top.cfg_gain_q[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20855_ (.CLK(clknet_leaf_29_io_wbs_clk),
    .D(_01151_),
    .Q(\wfg_stim_mem_top.cfg_gain_q[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20856_ (.CLK(clknet_leaf_25_io_wbs_clk),
    .D(_01152_),
    .Q(\wfg_stim_mem_top.cfg_gain_q[23] ));
 sky130_fd_sc_hd__dfxtp_2 _20857_ (.CLK(clknet_leaf_2_io_wbs_clk),
    .D(_01153_),
    .Q(\wfg_stim_mem_top.cfg_inc_q[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20858_ (.CLK(clknet_leaf_106_io_wbs_clk),
    .D(_01154_),
    .Q(\wfg_stim_mem_top.cfg_inc_q[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20859_ (.CLK(clknet_leaf_106_io_wbs_clk),
    .D(_01155_),
    .Q(\wfg_stim_mem_top.cfg_inc_q[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20860_ (.CLK(clknet_leaf_106_io_wbs_clk),
    .D(_01156_),
    .Q(\wfg_stim_mem_top.cfg_inc_q[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20861_ (.CLK(clknet_leaf_109_io_wbs_clk),
    .D(_01157_),
    .Q(\wfg_stim_mem_top.cfg_inc_q[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20862_ (.CLK(clknet_leaf_109_io_wbs_clk),
    .D(_01158_),
    .Q(\wfg_stim_mem_top.cfg_inc_q[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20863_ (.CLK(clknet_leaf_1_io_wbs_clk),
    .D(_01159_),
    .Q(\wfg_stim_mem_top.cfg_inc_q[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20864_ (.CLK(clknet_leaf_1_io_wbs_clk),
    .D(_01160_),
    .Q(\wfg_stim_mem_top.cfg_inc_q[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20865_ (.CLK(clknet_leaf_106_io_wbs_clk),
    .D(_01161_),
    .Q(\wfg_stim_mem_top.end_val_q[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20866_ (.CLK(clknet_leaf_107_io_wbs_clk),
    .D(_01162_),
    .Q(\wfg_stim_mem_top.end_val_q[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20867_ (.CLK(clknet_leaf_107_io_wbs_clk),
    .D(_01163_),
    .Q(\wfg_stim_mem_top.end_val_q[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20868_ (.CLK(clknet_leaf_105_io_wbs_clk),
    .D(_01164_),
    .Q(\wfg_stim_mem_top.end_val_q[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20869_ (.CLK(clknet_leaf_107_io_wbs_clk),
    .D(_01165_),
    .Q(\wfg_stim_mem_top.end_val_q[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20870_ (.CLK(clknet_leaf_107_io_wbs_clk),
    .D(_01166_),
    .Q(\wfg_stim_mem_top.end_val_q[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20871_ (.CLK(clknet_leaf_109_io_wbs_clk),
    .D(_01167_),
    .Q(\wfg_stim_mem_top.end_val_q[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20872_ (.CLK(clknet_leaf_1_io_wbs_clk),
    .D(_01168_),
    .Q(\wfg_stim_mem_top.end_val_q[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20873_ (.CLK(clknet_leaf_103_io_wbs_clk),
    .D(_01169_),
    .Q(\wfg_stim_mem_top.end_val_q[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20874_ (.CLK(clknet_leaf_105_io_wbs_clk),
    .D(_01170_),
    .Q(\wfg_stim_mem_top.end_val_q[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20875_ (.CLK(clknet_leaf_105_io_wbs_clk),
    .D(_01171_),
    .Q(\wfg_stim_mem_top.end_val_q[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20876_ (.CLK(clknet_leaf_105_io_wbs_clk),
    .D(_01172_),
    .Q(\wfg_stim_mem_top.end_val_q[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20877_ (.CLK(clknet_leaf_104_io_wbs_clk),
    .D(_01173_),
    .Q(\wfg_stim_mem_top.end_val_q[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20878_ (.CLK(clknet_leaf_105_io_wbs_clk),
    .D(_01174_),
    .Q(\wfg_stim_mem_top.end_val_q[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20879_ (.CLK(clknet_leaf_104_io_wbs_clk),
    .D(_01175_),
    .Q(\wfg_stim_mem_top.end_val_q[14] ));
 sky130_fd_sc_hd__dfxtp_2 _20880_ (.CLK(clknet_leaf_104_io_wbs_clk),
    .D(_01176_),
    .Q(\wfg_stim_mem_top.end_val_q[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20881_ (.CLK(clknet_leaf_106_io_wbs_clk),
    .D(_01177_),
    .Q(\wfg_stim_mem_top.start_val_q[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20882_ (.CLK(clknet_leaf_103_io_wbs_clk),
    .D(_01178_),
    .Q(\wfg_stim_mem_top.start_val_q[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20883_ (.CLK(clknet_leaf_107_io_wbs_clk),
    .D(_01179_),
    .Q(\wfg_stim_mem_top.start_val_q[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20884_ (.CLK(clknet_leaf_105_io_wbs_clk),
    .D(_01180_),
    .Q(\wfg_stim_mem_top.start_val_q[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20885_ (.CLK(clknet_leaf_106_io_wbs_clk),
    .D(_01181_),
    .Q(\wfg_stim_mem_top.start_val_q[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20886_ (.CLK(clknet_leaf_1_io_wbs_clk),
    .D(_01182_),
    .Q(\wfg_stim_mem_top.start_val_q[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20887_ (.CLK(clknet_leaf_1_io_wbs_clk),
    .D(_01183_),
    .Q(\wfg_stim_mem_top.start_val_q[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20888_ (.CLK(clknet_leaf_1_io_wbs_clk),
    .D(_01184_),
    .Q(\wfg_stim_mem_top.start_val_q[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20889_ (.CLK(clknet_leaf_1_io_wbs_clk),
    .D(_01185_),
    .Q(\wfg_stim_mem_top.start_val_q[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20890_ (.CLK(clknet_leaf_105_io_wbs_clk),
    .D(_01186_),
    .Q(\wfg_stim_mem_top.start_val_q[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20891_ (.CLK(clknet_leaf_105_io_wbs_clk),
    .D(_01187_),
    .Q(\wfg_stim_mem_top.start_val_q[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20892_ (.CLK(clknet_leaf_105_io_wbs_clk),
    .D(_01188_),
    .Q(\wfg_stim_mem_top.start_val_q[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20893_ (.CLK(clknet_leaf_104_io_wbs_clk),
    .D(_01189_),
    .Q(\wfg_stim_mem_top.start_val_q[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20894_ (.CLK(clknet_leaf_105_io_wbs_clk),
    .D(_01190_),
    .Q(\wfg_stim_mem_top.start_val_q[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20895_ (.CLK(clknet_leaf_104_io_wbs_clk),
    .D(_01191_),
    .Q(\wfg_stim_mem_top.start_val_q[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20896_ (.CLK(clknet_leaf_104_io_wbs_clk),
    .D(_01192_),
    .Q(\wfg_stim_mem_top.start_val_q[15] ));
 sky130_fd_sc_hd__dfrtp_4 _20897_ (.CLK(clknet_leaf_31_io_wbs_clk),
    .D(\wfg_drive_spi_top.wfg_drive_spi.next_state[0] ),
    .RESET_B(_00406_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.cur_state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _20898_ (.CLK(clknet_leaf_31_io_wbs_clk),
    .D(\wfg_drive_spi_top.wfg_drive_spi.next_state[1] ),
    .RESET_B(_00407_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.cur_state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _20899_ (.CLK(clknet_leaf_31_io_wbs_clk),
    .D(_00021_),
    .RESET_B(_00408_),
    .Q(net178));
 sky130_fd_sc_hd__dfrtp_4 _20900_ (.CLK(clknet_leaf_31_io_wbs_clk),
    .D(_00020_),
    .RESET_B(_00409_),
    .Q(net177));
 sky130_fd_sc_hd__dfrtp_4 _20901_ (.CLK(clknet_leaf_55_io_wbs_clk),
    .D(_00022_),
    .RESET_B(_00410_),
    .Q(net179));
 sky130_fd_sc_hd__dfxtp_1 _20902_ (.CLK(clknet_leaf_101_io_wbs_clk),
    .D(_01193_),
    .Q(\wfg_drive_pat_top.wbs_ack_o ));
 sky130_fd_sc_hd__dfrtp_1 _20903_ (.CLK(clknet_leaf_28_io_wbs_clk),
    .D(_01194_),
    .RESET_B(_00411_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _20904_ (.CLK(clknet_leaf_27_io_wbs_clk),
    .D(_01195_),
    .RESET_B(_00412_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _20905_ (.CLK(clknet_leaf_27_io_wbs_clk),
    .D(_01196_),
    .RESET_B(_00413_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _20906_ (.CLK(clknet_leaf_27_io_wbs_clk),
    .D(_01197_),
    .RESET_B(_00414_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _20907_ (.CLK(clknet_leaf_27_io_wbs_clk),
    .D(_01198_),
    .RESET_B(_00415_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.counter[4] ));
 sky130_fd_sc_hd__dfrtp_1 _20908_ (.CLK(clknet_leaf_27_io_wbs_clk),
    .D(_01199_),
    .RESET_B(_00416_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.counter[5] ));
 sky130_fd_sc_hd__dfrtp_1 _20909_ (.CLK(clknet_leaf_21_io_wbs_clk),
    .D(_01200_),
    .RESET_B(_00417_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.counter[6] ));
 sky130_fd_sc_hd__dfrtp_1 _20910_ (.CLK(clknet_leaf_21_io_wbs_clk),
    .D(_01201_),
    .RESET_B(_00418_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.counter[7] ));
 sky130_fd_sc_hd__dfrtp_1 _20911_ (.CLK(clknet_leaf_28_io_wbs_clk),
    .D(_01202_),
    .RESET_B(_00419_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.clk_div[0] ));
 sky130_fd_sc_hd__dfrtp_1 _20912_ (.CLK(clknet_leaf_27_io_wbs_clk),
    .D(_01203_),
    .RESET_B(_00420_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.clk_div[1] ));
 sky130_fd_sc_hd__dfrtp_1 _20913_ (.CLK(clknet_leaf_28_io_wbs_clk),
    .D(_01204_),
    .RESET_B(_00421_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.clk_div[2] ));
 sky130_fd_sc_hd__dfrtp_1 _20914_ (.CLK(clknet_leaf_22_io_wbs_clk),
    .D(_01205_),
    .RESET_B(_00422_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.clk_div[3] ));
 sky130_fd_sc_hd__dfrtp_1 _20915_ (.CLK(clknet_leaf_21_io_wbs_clk),
    .D(_01206_),
    .RESET_B(_00423_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.clk_div[4] ));
 sky130_fd_sc_hd__dfrtp_1 _20916_ (.CLK(clknet_leaf_21_io_wbs_clk),
    .D(_01207_),
    .RESET_B(_00424_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.clk_div[5] ));
 sky130_fd_sc_hd__dfrtp_1 _20917_ (.CLK(clknet_leaf_21_io_wbs_clk),
    .D(_01208_),
    .RESET_B(_00425_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.clk_div[6] ));
 sky130_fd_sc_hd__dfrtp_1 _20918_ (.CLK(clknet_leaf_21_io_wbs_clk),
    .D(_01209_),
    .RESET_B(_00426_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.clk_div[7] ));
 sky130_fd_sc_hd__dfrtp_1 _20919_ (.CLK(clknet_leaf_48_io_wbs_clk),
    .D(_01210_),
    .RESET_B(_00427_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.current_bit[0] ));
 sky130_fd_sc_hd__dfrtp_1 _20920_ (.CLK(clknet_leaf_48_io_wbs_clk),
    .D(_01211_),
    .RESET_B(_00428_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.current_bit[1] ));
 sky130_fd_sc_hd__dfrtp_1 _20921_ (.CLK(clknet_leaf_48_io_wbs_clk),
    .D(_01212_),
    .RESET_B(_00429_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.current_bit[2] ));
 sky130_fd_sc_hd__dfrtp_1 _20922_ (.CLK(clknet_leaf_48_io_wbs_clk),
    .D(_01213_),
    .RESET_B(_00430_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.current_bit[3] ));
 sky130_fd_sc_hd__dfrtp_1 _20923_ (.CLK(clknet_leaf_31_io_wbs_clk),
    .D(_01214_),
    .RESET_B(_00431_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.current_bit[4] ));
 sky130_fd_sc_hd__dfrtp_1 _20924_ (.CLK(clknet_leaf_33_io_wbs_clk),
    .D(_00003_),
    .RESET_B(_00432_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_cs ));
 sky130_fd_sc_hd__dfrtp_2 _20925_ (.CLK(clknet_leaf_48_io_wbs_clk),
    .D(_01215_),
    .RESET_B(_00433_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 _20926_ (.CLK(clknet_leaf_48_io_wbs_clk),
    .D(_01216_),
    .RESET_B(_00434_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 _20927_ (.CLK(clknet_leaf_49_io_wbs_clk),
    .D(_01217_),
    .RESET_B(_00435_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 _20928_ (.CLK(clknet_leaf_46_io_wbs_clk),
    .D(_01218_),
    .RESET_B(_00436_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 _20929_ (.CLK(clknet_leaf_46_io_wbs_clk),
    .D(_01219_),
    .RESET_B(_00437_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 _20930_ (.CLK(clknet_leaf_51_io_wbs_clk),
    .D(_01220_),
    .RESET_B(_00438_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 _20931_ (.CLK(clknet_leaf_46_io_wbs_clk),
    .D(_01221_),
    .RESET_B(_00439_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[6] ));
 sky130_fd_sc_hd__dfrtp_1 _20932_ (.CLK(clknet_leaf_51_io_wbs_clk),
    .D(_01222_),
    .RESET_B(_00440_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 _20933_ (.CLK(clknet_leaf_51_io_wbs_clk),
    .D(_01223_),
    .RESET_B(_00441_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[8] ));
 sky130_fd_sc_hd__dfrtp_1 _20934_ (.CLK(clknet_leaf_51_io_wbs_clk),
    .D(_01224_),
    .RESET_B(_00442_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[9] ));
 sky130_fd_sc_hd__dfrtp_1 _20935_ (.CLK(clknet_leaf_52_io_wbs_clk),
    .D(_01225_),
    .RESET_B(_00443_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[10] ));
 sky130_fd_sc_hd__dfrtp_1 _20936_ (.CLK(clknet_leaf_52_io_wbs_clk),
    .D(_01226_),
    .RESET_B(_00444_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[11] ));
 sky130_fd_sc_hd__dfrtp_1 _20937_ (.CLK(clknet_leaf_52_io_wbs_clk),
    .D(_01227_),
    .RESET_B(_00445_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[12] ));
 sky130_fd_sc_hd__dfrtp_1 _20938_ (.CLK(clknet_leaf_52_io_wbs_clk),
    .D(_01228_),
    .RESET_B(_00446_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[13] ));
 sky130_fd_sc_hd__dfrtp_1 _20939_ (.CLK(clknet_leaf_53_io_wbs_clk),
    .D(_01229_),
    .RESET_B(_00447_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[14] ));
 sky130_fd_sc_hd__dfrtp_1 _20940_ (.CLK(clknet_leaf_53_io_wbs_clk),
    .D(_01230_),
    .RESET_B(_00448_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[15] ));
 sky130_fd_sc_hd__dfrtp_1 _20941_ (.CLK(clknet_leaf_53_io_wbs_clk),
    .D(_01231_),
    .RESET_B(_00449_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[16] ));
 sky130_fd_sc_hd__dfrtp_1 _20942_ (.CLK(clknet_leaf_53_io_wbs_clk),
    .D(_01232_),
    .RESET_B(_00450_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[17] ));
 sky130_fd_sc_hd__dfrtp_1 _20943_ (.CLK(clknet_leaf_61_io_wbs_clk),
    .D(_01233_),
    .RESET_B(_00451_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[18] ));
 sky130_fd_sc_hd__dfrtp_1 _20944_ (.CLK(clknet_leaf_61_io_wbs_clk),
    .D(_01234_),
    .RESET_B(_00452_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[19] ));
 sky130_fd_sc_hd__dfrtp_1 _20945_ (.CLK(clknet_leaf_59_io_wbs_clk),
    .D(_01235_),
    .RESET_B(_00453_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[20] ));
 sky130_fd_sc_hd__dfrtp_1 _20946_ (.CLK(clknet_leaf_58_io_wbs_clk),
    .D(_01236_),
    .RESET_B(_00454_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[21] ));
 sky130_fd_sc_hd__dfrtp_1 _20947_ (.CLK(clknet_leaf_59_io_wbs_clk),
    .D(_01237_),
    .RESET_B(_00455_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[22] ));
 sky130_fd_sc_hd__dfrtp_2 _20948_ (.CLK(clknet_leaf_59_io_wbs_clk),
    .D(_01238_),
    .RESET_B(_00456_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[23] ));
 sky130_fd_sc_hd__dfrtp_1 _20949_ (.CLK(clknet_leaf_59_io_wbs_clk),
    .D(_01239_),
    .RESET_B(_00457_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[24] ));
 sky130_fd_sc_hd__dfrtp_1 _20950_ (.CLK(clknet_leaf_59_io_wbs_clk),
    .D(_01240_),
    .RESET_B(_00458_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[25] ));
 sky130_fd_sc_hd__dfrtp_1 _20951_ (.CLK(clknet_leaf_58_io_wbs_clk),
    .D(_01241_),
    .RESET_B(_00459_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[26] ));
 sky130_fd_sc_hd__dfrtp_1 _20952_ (.CLK(clknet_leaf_57_io_wbs_clk),
    .D(_01242_),
    .RESET_B(_00460_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[27] ));
 sky130_fd_sc_hd__dfrtp_1 _20953_ (.CLK(clknet_leaf_58_io_wbs_clk),
    .D(_01243_),
    .RESET_B(_00461_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[28] ));
 sky130_fd_sc_hd__dfrtp_1 _20954_ (.CLK(clknet_leaf_58_io_wbs_clk),
    .D(_01244_),
    .RESET_B(_00462_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[29] ));
 sky130_fd_sc_hd__dfrtp_1 _20955_ (.CLK(clknet_leaf_58_io_wbs_clk),
    .D(_01245_),
    .RESET_B(_00463_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[30] ));
 sky130_fd_sc_hd__dfrtp_1 _20956_ (.CLK(clknet_leaf_58_io_wbs_clk),
    .D(_01246_),
    .RESET_B(_00464_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_data[31] ));
 sky130_fd_sc_hd__dfrtp_1 _20957_ (.CLK(clknet_leaf_31_io_wbs_clk),
    .D(_01247_),
    .RESET_B(_00465_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.spi_clk ));
 sky130_fd_sc_hd__dfrtp_1 _20958_ (.CLK(clknet_leaf_33_io_wbs_clk),
    .D(_01248_),
    .RESET_B(_00466_),
    .Q(\wfg_drive_spi_top.wfg_axis_tready_o ));
 sky130_fd_sc_hd__dfrtp_4 _20959_ (.CLK(clknet_leaf_49_io_wbs_clk),
    .D(_01249_),
    .RESET_B(_00467_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.lsbfirst ));
 sky130_fd_sc_hd__dfrtp_1 _20960_ (.CLK(clknet_leaf_33_io_wbs_clk),
    .D(_01250_),
    .RESET_B(_00468_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.cpol ));
 sky130_fd_sc_hd__dfrtp_1 _20961_ (.CLK(clknet_leaf_33_io_wbs_clk),
    .D(_01251_),
    .RESET_B(_00469_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.cspol ));
 sky130_fd_sc_hd__dfrtp_4 _20962_ (.CLK(clknet_leaf_31_io_wbs_clk),
    .D(_01252_),
    .RESET_B(_00470_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.byte_cnt[0] ));
 sky130_fd_sc_hd__dfrtp_4 _20963_ (.CLK(clknet_leaf_19_io_wbs_clk),
    .D(_01253_),
    .RESET_B(_00471_),
    .Q(\wfg_drive_spi_top.wfg_drive_spi.byte_cnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20964_ (.CLK(clknet_leaf_98_io_wbs_clk),
    .D(_01254_),
    .Q(\wfg_core_top.wbs_dat_o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20965_ (.CLK(clknet_leaf_101_io_wbs_clk),
    .D(_01255_),
    .Q(\wfg_core_top.wbs_dat_o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20966_ (.CLK(clknet_leaf_100_io_wbs_clk),
    .D(_01256_),
    .Q(\wfg_core_top.wbs_dat_o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20967_ (.CLK(clknet_leaf_100_io_wbs_clk),
    .D(_01257_),
    .Q(\wfg_core_top.wbs_dat_o[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20968_ (.CLK(clknet_leaf_100_io_wbs_clk),
    .D(_01258_),
    .Q(\wfg_core_top.wbs_dat_o[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20969_ (.CLK(clknet_leaf_100_io_wbs_clk),
    .D(_01259_),
    .Q(\wfg_core_top.wbs_dat_o[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20970_ (.CLK(clknet_leaf_100_io_wbs_clk),
    .D(_01260_),
    .Q(\wfg_core_top.wbs_dat_o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20971_ (.CLK(clknet_leaf_100_io_wbs_clk),
    .D(_01261_),
    .Q(\wfg_core_top.wbs_dat_o[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20972_ (.CLK(clknet_leaf_100_io_wbs_clk),
    .D(_01262_),
    .Q(\wfg_core_top.wbs_dat_o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20973_ (.CLK(clknet_leaf_98_io_wbs_clk),
    .D(_01263_),
    .Q(\wfg_core_top.wbs_dat_o[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20974_ (.CLK(clknet_leaf_98_io_wbs_clk),
    .D(_01264_),
    .Q(\wfg_core_top.wbs_dat_o[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20975_ (.CLK(clknet_leaf_98_io_wbs_clk),
    .D(_01265_),
    .Q(\wfg_core_top.wbs_dat_o[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20976_ (.CLK(clknet_leaf_95_io_wbs_clk),
    .D(_01266_),
    .Q(\wfg_core_top.wbs_dat_o[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20977_ (.CLK(clknet_leaf_94_io_wbs_clk),
    .D(_01267_),
    .Q(\wfg_core_top.wbs_dat_o[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20978_ (.CLK(clknet_leaf_95_io_wbs_clk),
    .D(_01268_),
    .Q(\wfg_core_top.wbs_dat_o[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20979_ (.CLK(clknet_leaf_95_io_wbs_clk),
    .D(_01269_),
    .Q(\wfg_core_top.wbs_dat_o[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20980_ (.CLK(clknet_leaf_95_io_wbs_clk),
    .D(_01270_),
    .Q(\wfg_core_top.wbs_dat_o[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20981_ (.CLK(clknet_leaf_95_io_wbs_clk),
    .D(_01271_),
    .Q(\wfg_core_top.wbs_dat_o[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20982_ (.CLK(clknet_leaf_96_io_wbs_clk),
    .D(_01272_),
    .Q(\wfg_core_top.wbs_dat_o[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20983_ (.CLK(clknet_leaf_95_io_wbs_clk),
    .D(_01273_),
    .Q(\wfg_core_top.wbs_dat_o[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20984_ (.CLK(clknet_leaf_96_io_wbs_clk),
    .D(_01274_),
    .Q(\wfg_core_top.wbs_dat_o[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20985_ (.CLK(clknet_leaf_80_io_wbs_clk),
    .D(_01275_),
    .Q(\wfg_core_top.wbs_dat_o[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20986_ (.CLK(clknet_leaf_80_io_wbs_clk),
    .D(_01276_),
    .Q(\wfg_core_top.wbs_dat_o[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20987_ (.CLK(clknet_leaf_79_io_wbs_clk),
    .D(_01277_),
    .Q(\wfg_core_top.wbs_dat_o[23] ));
 sky130_fd_sc_hd__dfxtp_1 _20988_ (.CLK(clknet_leaf_18_io_wbs_clk),
    .D(_01278_),
    .Q(\wfg_drive_spi_top.ctrl_en_q ));
 sky130_fd_sc_hd__dfxtp_1 _20989_ (.CLK(clknet_leaf_18_io_wbs_clk),
    .D(_01279_),
    .Q(\wfg_drive_spi_top.cfg_core_sel_q ));
 sky130_fd_sc_hd__dfxtp_1 _20990_ (.CLK(clknet_leaf_17_io_wbs_clk),
    .D(_01280_),
    .Q(\wfg_drive_spi_top.cfg_cpol_q ));
 sky130_fd_sc_hd__dfxtp_1 _20991_ (.CLK(clknet_leaf_17_io_wbs_clk),
    .D(_01281_),
    .Q(\wfg_drive_spi_top.cfg_dff_q[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20992_ (.CLK(clknet_leaf_19_io_wbs_clk),
    .D(_01282_),
    .Q(\wfg_drive_spi_top.cfg_dff_q[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20993_ (.CLK(clknet_leaf_19_io_wbs_clk),
    .D(_01283_),
    .Q(\wfg_drive_spi_top.cfg_lsbfirst_q ));
 sky130_fd_sc_hd__dfxtp_1 _20994_ (.CLK(clknet_leaf_19_io_wbs_clk),
    .D(_01284_),
    .Q(\wfg_drive_spi_top.cfg_sspol_q ));
 sky130_fd_sc_hd__dfxtp_1 _20995_ (.CLK(clknet_leaf_19_io_wbs_clk),
    .D(_01285_),
    .Q(\wfg_drive_spi_top.clkcfg_div_q[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20996_ (.CLK(clknet_leaf_19_io_wbs_clk),
    .D(_01286_),
    .Q(\wfg_drive_spi_top.clkcfg_div_q[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20997_ (.CLK(clknet_leaf_19_io_wbs_clk),
    .D(_01287_),
    .Q(\wfg_drive_spi_top.clkcfg_div_q[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20998_ (.CLK(clknet_leaf_19_io_wbs_clk),
    .D(_01288_),
    .Q(\wfg_drive_spi_top.clkcfg_div_q[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20999_ (.CLK(clknet_leaf_21_io_wbs_clk),
    .D(_01289_),
    .Q(\wfg_drive_spi_top.clkcfg_div_q[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21000_ (.CLK(clknet_leaf_19_io_wbs_clk),
    .D(_01290_),
    .Q(\wfg_drive_spi_top.clkcfg_div_q[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21001_ (.CLK(clknet_leaf_21_io_wbs_clk),
    .D(_01291_),
    .Q(\wfg_drive_spi_top.clkcfg_div_q[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21002_ (.CLK(clknet_leaf_21_io_wbs_clk),
    .D(_01292_),
    .Q(\wfg_drive_spi_top.clkcfg_div_q[7] ));
 sky130_fd_sc_hd__conb_1 wfg_top_181 (.LO(net181));
 sky130_fd_sc_hd__conb_1 wfg_top_182 (.LO(net182));
 sky130_fd_sc_hd__conb_1 wfg_top_183 (.LO(net183));
 sky130_fd_sc_hd__conb_1 wfg_top_184 (.LO(net184));
 sky130_fd_sc_hd__conb_1 wfg_top_185 (.LO(net185));
 sky130_fd_sc_hd__conb_1 wfg_top_186 (.LO(net186));
 sky130_fd_sc_hd__conb_1 wfg_top_187 (.LO(net187));
 sky130_fd_sc_hd__conb_1 wfg_top_188 (.LO(net188));
 sky130_fd_sc_hd__conb_1 wfg_top_189 (.LO(net189));
 sky130_fd_sc_hd__conb_1 wfg_top_190 (.LO(net190));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_io_wbs_clk (.A(clknet_3_0_0_io_wbs_clk),
    .X(clknet_leaf_0_io_wbs_clk));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5973 ();
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(dout1[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(dout1[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input3 (.A(dout1[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(dout1[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(dout1[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(dout1[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(dout1[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(dout1[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 input9 (.A(dout1[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(dout1[18]),
    .X(net10));
 sky130_fd_sc_hd__dlymetal6s2s_1 input11 (.A(dout1[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(dout1[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(dout1[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(dout1[21]),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(dout1[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(dout1[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(dout1[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(dout1[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(dout1[26]),
    .X(net19));
 sky130_fd_sc_hd__dlymetal6s2s_1 input20 (.A(dout1[27]),
    .X(net20));
 sky130_fd_sc_hd__dlymetal6s2s_1 input21 (.A(dout1[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(dout1[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 input23 (.A(dout1[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(dout1[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_4 input25 (.A(dout1[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_2 input26 (.A(dout1[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(dout1[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(dout1[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_2 input29 (.A(dout1[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(dout1[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(dout1[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(dout1[9]),
    .X(net32));
 sky130_fd_sc_hd__dlymetal6s2s_1 input33 (.A(io_wbs_adr[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(io_wbs_adr[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(io_wbs_adr[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(io_wbs_adr[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(io_wbs_adr[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(io_wbs_adr[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(io_wbs_adr[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(io_wbs_adr[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(io_wbs_adr[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(io_wbs_adr[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(io_wbs_adr[19]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(io_wbs_adr[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(io_wbs_adr[20]),
    .X(net45));
 sky130_fd_sc_hd__buf_2 input46 (.A(io_wbs_adr[21]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(io_wbs_adr[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(io_wbs_adr[23]),
    .X(net48));
 sky130_fd_sc_hd__dlymetal6s2s_1 input49 (.A(io_wbs_adr[24]),
    .X(net49));
 sky130_fd_sc_hd__dlymetal6s2s_1 input50 (.A(io_wbs_adr[25]),
    .X(net50));
 sky130_fd_sc_hd__dlymetal6s2s_1 input51 (.A(io_wbs_adr[26]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(io_wbs_adr[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(io_wbs_adr[28]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(io_wbs_adr[29]),
    .X(net54));
 sky130_fd_sc_hd__buf_2 input55 (.A(io_wbs_adr[2]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(io_wbs_adr[30]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(io_wbs_adr[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_4 input58 (.A(io_wbs_adr[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_2 input59 (.A(io_wbs_adr[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(io_wbs_adr[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 input61 (.A(io_wbs_adr[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(io_wbs_adr[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(io_wbs_adr[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(io_wbs_adr[9]),
    .X(net64));
 sky130_fd_sc_hd__buf_2 input65 (.A(io_wbs_cyc),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_4 input66 (.A(io_wbs_datwr[0]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 input67 (.A(io_wbs_datwr[10]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 input68 (.A(io_wbs_datwr[11]),
    .X(net68));
 sky130_fd_sc_hd__buf_2 input69 (.A(io_wbs_datwr[12]),
    .X(net69));
 sky130_fd_sc_hd__buf_2 input70 (.A(io_wbs_datwr[13]),
    .X(net70));
 sky130_fd_sc_hd__buf_4 input71 (.A(io_wbs_datwr[14]),
    .X(net71));
 sky130_fd_sc_hd__buf_2 input72 (.A(io_wbs_datwr[15]),
    .X(net72));
 sky130_fd_sc_hd__buf_8 input73 (.A(io_wbs_datwr[16]),
    .X(net73));
 sky130_fd_sc_hd__buf_8 input74 (.A(io_wbs_datwr[17]),
    .X(net74));
 sky130_fd_sc_hd__buf_6 input75 (.A(io_wbs_datwr[18]),
    .X(net75));
 sky130_fd_sc_hd__buf_6 input76 (.A(io_wbs_datwr[19]),
    .X(net76));
 sky130_fd_sc_hd__buf_8 input77 (.A(io_wbs_datwr[1]),
    .X(net77));
 sky130_fd_sc_hd__buf_6 input78 (.A(io_wbs_datwr[20]),
    .X(net78));
 sky130_fd_sc_hd__buf_6 input79 (.A(io_wbs_datwr[21]),
    .X(net79));
 sky130_fd_sc_hd__buf_6 input80 (.A(io_wbs_datwr[22]),
    .X(net80));
 sky130_fd_sc_hd__buf_6 input81 (.A(io_wbs_datwr[23]),
    .X(net81));
 sky130_fd_sc_hd__buf_2 input82 (.A(io_wbs_datwr[24]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_4 input83 (.A(io_wbs_datwr[25]),
    .X(net83));
 sky130_fd_sc_hd__buf_2 input84 (.A(io_wbs_datwr[26]),
    .X(net84));
 sky130_fd_sc_hd__buf_2 input85 (.A(io_wbs_datwr[27]),
    .X(net85));
 sky130_fd_sc_hd__buf_2 input86 (.A(io_wbs_datwr[28]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_4 input87 (.A(io_wbs_datwr[29]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_4 input88 (.A(io_wbs_datwr[2]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_4 input89 (.A(io_wbs_datwr[30]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_4 input90 (.A(io_wbs_datwr[31]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_4 input91 (.A(io_wbs_datwr[3]),
    .X(net91));
 sky130_fd_sc_hd__buf_4 input92 (.A(io_wbs_datwr[4]),
    .X(net92));
 sky130_fd_sc_hd__buf_4 input93 (.A(io_wbs_datwr[5]),
    .X(net93));
 sky130_fd_sc_hd__buf_2 input94 (.A(io_wbs_datwr[6]),
    .X(net94));
 sky130_fd_sc_hd__buf_2 input95 (.A(io_wbs_datwr[7]),
    .X(net95));
 sky130_fd_sc_hd__buf_2 input96 (.A(io_wbs_datwr[8]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 input97 (.A(io_wbs_datwr[9]),
    .X(net97));
 sky130_fd_sc_hd__buf_8 input98 (.A(io_wbs_rst),
    .X(net98));
 sky130_fd_sc_hd__buf_4 input99 (.A(io_wbs_stb),
    .X(net99));
 sky130_fd_sc_hd__buf_2 input100 (.A(io_wbs_we),
    .X(net100));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(addr1[0]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(addr1[1]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(addr1[2]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(addr1[3]));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .X(addr1[4]));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .X(addr1[5]));
 sky130_fd_sc_hd__buf_2 output107 (.A(net107),
    .X(addr1[6]));
 sky130_fd_sc_hd__buf_2 output108 (.A(net108),
    .X(addr1[7]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net109),
    .X(addr1[8]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net110),
    .X(addr1[9]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net111),
    .X(csb1));
 sky130_fd_sc_hd__buf_2 output112 (.A(net112),
    .X(io_wbs_ack));
 sky130_fd_sc_hd__buf_2 output113 (.A(net113),
    .X(io_wbs_datrd[0]));
 sky130_fd_sc_hd__buf_2 output114 (.A(net114),
    .X(io_wbs_datrd[10]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net115),
    .X(io_wbs_datrd[11]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net116),
    .X(io_wbs_datrd[12]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net117),
    .X(io_wbs_datrd[13]));
 sky130_fd_sc_hd__buf_2 output118 (.A(net118),
    .X(io_wbs_datrd[14]));
 sky130_fd_sc_hd__buf_2 output119 (.A(net119),
    .X(io_wbs_datrd[15]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net120),
    .X(io_wbs_datrd[16]));
 sky130_fd_sc_hd__buf_2 output121 (.A(net121),
    .X(io_wbs_datrd[17]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net122),
    .X(io_wbs_datrd[18]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net123),
    .X(io_wbs_datrd[19]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net124),
    .X(io_wbs_datrd[1]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net125),
    .X(io_wbs_datrd[20]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net126),
    .X(io_wbs_datrd[21]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net127),
    .X(io_wbs_datrd[22]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net128),
    .X(io_wbs_datrd[23]));
 sky130_fd_sc_hd__buf_2 output129 (.A(net129),
    .X(io_wbs_datrd[24]));
 sky130_fd_sc_hd__buf_2 output130 (.A(net130),
    .X(io_wbs_datrd[25]));
 sky130_fd_sc_hd__buf_2 output131 (.A(net131),
    .X(io_wbs_datrd[26]));
 sky130_fd_sc_hd__buf_2 output132 (.A(net132),
    .X(io_wbs_datrd[27]));
 sky130_fd_sc_hd__buf_2 output133 (.A(net133),
    .X(io_wbs_datrd[28]));
 sky130_fd_sc_hd__buf_2 output134 (.A(net134),
    .X(io_wbs_datrd[29]));
 sky130_fd_sc_hd__buf_2 output135 (.A(net135),
    .X(io_wbs_datrd[2]));
 sky130_fd_sc_hd__buf_2 output136 (.A(net136),
    .X(io_wbs_datrd[30]));
 sky130_fd_sc_hd__buf_2 output137 (.A(net137),
    .X(io_wbs_datrd[31]));
 sky130_fd_sc_hd__buf_2 output138 (.A(net138),
    .X(io_wbs_datrd[3]));
 sky130_fd_sc_hd__buf_2 output139 (.A(net139),
    .X(io_wbs_datrd[4]));
 sky130_fd_sc_hd__buf_2 output140 (.A(net140),
    .X(io_wbs_datrd[5]));
 sky130_fd_sc_hd__buf_2 output141 (.A(net141),
    .X(io_wbs_datrd[6]));
 sky130_fd_sc_hd__buf_2 output142 (.A(net142),
    .X(io_wbs_datrd[7]));
 sky130_fd_sc_hd__buf_2 output143 (.A(net143),
    .X(io_wbs_datrd[8]));
 sky130_fd_sc_hd__buf_2 output144 (.A(net144),
    .X(io_wbs_datrd[9]));
 sky130_fd_sc_hd__buf_2 output145 (.A(net145),
    .X(wfg_drive_pat_dout_o[0]));
 sky130_fd_sc_hd__buf_2 output146 (.A(net146),
    .X(wfg_drive_pat_dout_o[10]));
 sky130_fd_sc_hd__buf_2 output147 (.A(net147),
    .X(wfg_drive_pat_dout_o[11]));
 sky130_fd_sc_hd__buf_2 output148 (.A(net148),
    .X(wfg_drive_pat_dout_o[12]));
 sky130_fd_sc_hd__buf_2 output149 (.A(net149),
    .X(wfg_drive_pat_dout_o[13]));
 sky130_fd_sc_hd__buf_2 output150 (.A(net150),
    .X(wfg_drive_pat_dout_o[14]));
 sky130_fd_sc_hd__buf_2 output151 (.A(net151),
    .X(wfg_drive_pat_dout_o[15]));
 sky130_fd_sc_hd__buf_2 output152 (.A(net152),
    .X(wfg_drive_pat_dout_o[16]));
 sky130_fd_sc_hd__buf_2 output153 (.A(net153),
    .X(wfg_drive_pat_dout_o[17]));
 sky130_fd_sc_hd__buf_2 output154 (.A(net154),
    .X(wfg_drive_pat_dout_o[18]));
 sky130_fd_sc_hd__buf_2 output155 (.A(net155),
    .X(wfg_drive_pat_dout_o[19]));
 sky130_fd_sc_hd__buf_2 output156 (.A(net156),
    .X(wfg_drive_pat_dout_o[1]));
 sky130_fd_sc_hd__buf_2 output157 (.A(net157),
    .X(wfg_drive_pat_dout_o[20]));
 sky130_fd_sc_hd__buf_2 output158 (.A(net158),
    .X(wfg_drive_pat_dout_o[21]));
 sky130_fd_sc_hd__buf_2 output159 (.A(net159),
    .X(wfg_drive_pat_dout_o[22]));
 sky130_fd_sc_hd__buf_2 output160 (.A(net160),
    .X(wfg_drive_pat_dout_o[23]));
 sky130_fd_sc_hd__buf_2 output161 (.A(net161),
    .X(wfg_drive_pat_dout_o[24]));
 sky130_fd_sc_hd__buf_2 output162 (.A(net162),
    .X(wfg_drive_pat_dout_o[25]));
 sky130_fd_sc_hd__buf_2 output163 (.A(net163),
    .X(wfg_drive_pat_dout_o[26]));
 sky130_fd_sc_hd__buf_2 output164 (.A(net164),
    .X(wfg_drive_pat_dout_o[27]));
 sky130_fd_sc_hd__buf_2 output165 (.A(net165),
    .X(wfg_drive_pat_dout_o[28]));
 sky130_fd_sc_hd__buf_2 output166 (.A(net166),
    .X(wfg_drive_pat_dout_o[29]));
 sky130_fd_sc_hd__buf_2 output167 (.A(net167),
    .X(wfg_drive_pat_dout_o[2]));
 sky130_fd_sc_hd__buf_2 output168 (.A(net168),
    .X(wfg_drive_pat_dout_o[30]));
 sky130_fd_sc_hd__buf_2 output169 (.A(net169),
    .X(wfg_drive_pat_dout_o[31]));
 sky130_fd_sc_hd__buf_2 output170 (.A(net170),
    .X(wfg_drive_pat_dout_o[3]));
 sky130_fd_sc_hd__buf_2 output171 (.A(net171),
    .X(wfg_drive_pat_dout_o[4]));
 sky130_fd_sc_hd__buf_2 output172 (.A(net172),
    .X(wfg_drive_pat_dout_o[5]));
 sky130_fd_sc_hd__buf_2 output173 (.A(net173),
    .X(wfg_drive_pat_dout_o[6]));
 sky130_fd_sc_hd__buf_2 output174 (.A(net174),
    .X(wfg_drive_pat_dout_o[7]));
 sky130_fd_sc_hd__buf_2 output175 (.A(net175),
    .X(wfg_drive_pat_dout_o[8]));
 sky130_fd_sc_hd__buf_2 output176 (.A(net176),
    .X(wfg_drive_pat_dout_o[9]));
 sky130_fd_sc_hd__buf_2 output177 (.A(net177),
    .X(wfg_drive_spi_cs_no));
 sky130_fd_sc_hd__buf_2 output178 (.A(net178),
    .X(wfg_drive_spi_sclk_o));
 sky130_fd_sc_hd__buf_2 output179 (.A(net179),
    .X(wfg_drive_spi_sdo_o));
 sky130_fd_sc_hd__conb_1 wfg_top_180 (.LO(net180));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_io_wbs_clk (.A(clknet_3_0_0_io_wbs_clk),
    .X(clknet_leaf_1_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_io_wbs_clk (.A(clknet_3_0_0_io_wbs_clk),
    .X(clknet_leaf_2_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_io_wbs_clk (.A(clknet_3_0_0_io_wbs_clk),
    .X(clknet_leaf_3_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_io_wbs_clk (.A(clknet_3_0_0_io_wbs_clk),
    .X(clknet_leaf_4_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_io_wbs_clk (.A(clknet_opt_1_0_io_wbs_clk),
    .X(clknet_leaf_5_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_io_wbs_clk (.A(clknet_opt_2_0_io_wbs_clk),
    .X(clknet_leaf_6_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_io_wbs_clk (.A(clknet_3_2_0_io_wbs_clk),
    .X(clknet_leaf_7_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_io_wbs_clk (.A(clknet_3_2_0_io_wbs_clk),
    .X(clknet_leaf_8_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_io_wbs_clk (.A(clknet_3_2_0_io_wbs_clk),
    .X(clknet_leaf_9_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_io_wbs_clk (.A(clknet_3_2_0_io_wbs_clk),
    .X(clknet_leaf_10_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_io_wbs_clk (.A(clknet_3_0_0_io_wbs_clk),
    .X(clknet_leaf_11_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_io_wbs_clk (.A(clknet_3_1_0_io_wbs_clk),
    .X(clknet_leaf_12_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_io_wbs_clk (.A(clknet_3_3_0_io_wbs_clk),
    .X(clknet_leaf_13_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_io_wbs_clk (.A(clknet_3_3_0_io_wbs_clk),
    .X(clknet_leaf_14_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_io_wbs_clk (.A(clknet_3_3_0_io_wbs_clk),
    .X(clknet_leaf_15_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_io_wbs_clk (.A(clknet_3_3_0_io_wbs_clk),
    .X(clknet_leaf_16_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_io_wbs_clk (.A(clknet_3_3_0_io_wbs_clk),
    .X(clknet_leaf_17_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_io_wbs_clk (.A(clknet_3_3_0_io_wbs_clk),
    .X(clknet_leaf_18_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_io_wbs_clk (.A(clknet_3_3_0_io_wbs_clk),
    .X(clknet_leaf_19_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_io_wbs_clk (.A(clknet_3_3_0_io_wbs_clk),
    .X(clknet_leaf_20_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_io_wbs_clk (.A(clknet_3_2_0_io_wbs_clk),
    .X(clknet_leaf_21_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_io_wbs_clk (.A(clknet_3_2_0_io_wbs_clk),
    .X(clknet_leaf_22_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_io_wbs_clk (.A(clknet_3_2_0_io_wbs_clk),
    .X(clknet_leaf_23_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_io_wbs_clk (.A(clknet_3_2_0_io_wbs_clk),
    .X(clknet_leaf_24_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_io_wbs_clk (.A(clknet_3_2_0_io_wbs_clk),
    .X(clknet_leaf_25_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_io_wbs_clk (.A(clknet_3_2_0_io_wbs_clk),
    .X(clknet_leaf_26_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_io_wbs_clk (.A(clknet_3_2_0_io_wbs_clk),
    .X(clknet_leaf_27_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_io_wbs_clk (.A(clknet_3_2_0_io_wbs_clk),
    .X(clknet_leaf_28_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_io_wbs_clk (.A(clknet_3_2_0_io_wbs_clk),
    .X(clknet_leaf_29_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_io_wbs_clk (.A(clknet_3_4_0_io_wbs_clk),
    .X(clknet_leaf_31_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_io_wbs_clk (.A(clknet_3_4_0_io_wbs_clk),
    .X(clknet_leaf_32_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_io_wbs_clk (.A(clknet_3_3_0_io_wbs_clk),
    .X(clknet_leaf_33_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_io_wbs_clk (.A(clknet_3_3_0_io_wbs_clk),
    .X(clknet_leaf_34_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_io_wbs_clk (.A(clknet_3_3_0_io_wbs_clk),
    .X(clknet_leaf_35_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_io_wbs_clk (.A(clknet_3_4_0_io_wbs_clk),
    .X(clknet_leaf_36_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_io_wbs_clk (.A(clknet_3_4_0_io_wbs_clk),
    .X(clknet_leaf_37_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_io_wbs_clk (.A(clknet_3_4_0_io_wbs_clk),
    .X(clknet_leaf_38_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_io_wbs_clk (.A(clknet_3_4_0_io_wbs_clk),
    .X(clknet_leaf_39_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_io_wbs_clk (.A(clknet_3_4_0_io_wbs_clk),
    .X(clknet_leaf_40_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_io_wbs_clk (.A(clknet_3_4_0_io_wbs_clk),
    .X(clknet_leaf_41_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_io_wbs_clk (.A(clknet_3_4_0_io_wbs_clk),
    .X(clknet_leaf_42_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_io_wbs_clk (.A(clknet_3_6_0_io_wbs_clk),
    .X(clknet_leaf_43_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_io_wbs_clk (.A(clknet_3_6_0_io_wbs_clk),
    .X(clknet_leaf_44_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_io_wbs_clk (.A(clknet_3_6_0_io_wbs_clk),
    .X(clknet_leaf_45_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_io_wbs_clk (.A(clknet_3_6_0_io_wbs_clk),
    .X(clknet_leaf_46_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_io_wbs_clk (.A(clknet_3_6_0_io_wbs_clk),
    .X(clknet_leaf_47_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_io_wbs_clk (.A(clknet_3_4_0_io_wbs_clk),
    .X(clknet_leaf_48_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_io_wbs_clk (.A(clknet_3_6_0_io_wbs_clk),
    .X(clknet_leaf_49_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_io_wbs_clk (.A(clknet_3_6_0_io_wbs_clk),
    .X(clknet_leaf_50_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_io_wbs_clk (.A(clknet_3_6_0_io_wbs_clk),
    .X(clknet_leaf_51_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_io_wbs_clk (.A(clknet_3_6_0_io_wbs_clk),
    .X(clknet_leaf_52_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_io_wbs_clk (.A(clknet_3_7_0_io_wbs_clk),
    .X(clknet_leaf_53_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_io_wbs_clk (.A(clknet_3_7_0_io_wbs_clk),
    .X(clknet_leaf_54_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_io_wbs_clk (.A(clknet_3_7_0_io_wbs_clk),
    .X(clknet_leaf_55_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_io_wbs_clk (.A(clknet_3_7_0_io_wbs_clk),
    .X(clknet_leaf_56_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_io_wbs_clk (.A(clknet_opt_4_0_io_wbs_clk),
    .X(clknet_leaf_57_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_io_wbs_clk (.A(clknet_3_7_0_io_wbs_clk),
    .X(clknet_leaf_58_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_io_wbs_clk (.A(clknet_3_7_0_io_wbs_clk),
    .X(clknet_leaf_59_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_io_wbs_clk (.A(clknet_3_7_0_io_wbs_clk),
    .X(clknet_leaf_60_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_io_wbs_clk (.A(clknet_3_7_0_io_wbs_clk),
    .X(clknet_leaf_61_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_io_wbs_clk (.A(clknet_3_7_0_io_wbs_clk),
    .X(clknet_leaf_62_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_io_wbs_clk (.A(clknet_3_7_0_io_wbs_clk),
    .X(clknet_leaf_63_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_io_wbs_clk (.A(clknet_3_7_0_io_wbs_clk),
    .X(clknet_leaf_64_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_io_wbs_clk (.A(clknet_3_7_0_io_wbs_clk),
    .X(clknet_leaf_65_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_io_wbs_clk (.A(clknet_3_7_0_io_wbs_clk),
    .X(clknet_leaf_66_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_io_wbs_clk (.A(clknet_3_7_0_io_wbs_clk),
    .X(clknet_leaf_67_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_io_wbs_clk (.A(clknet_3_7_0_io_wbs_clk),
    .X(clknet_leaf_68_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_io_wbs_clk (.A(clknet_3_6_0_io_wbs_clk),
    .X(clknet_leaf_69_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_io_wbs_clk (.A(clknet_3_6_0_io_wbs_clk),
    .X(clknet_leaf_70_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_io_wbs_clk (.A(clknet_3_6_0_io_wbs_clk),
    .X(clknet_leaf_71_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_io_wbs_clk (.A(clknet_3_5_0_io_wbs_clk),
    .X(clknet_leaf_72_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_io_wbs_clk (.A(clknet_3_5_0_io_wbs_clk),
    .X(clknet_leaf_73_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_io_wbs_clk (.A(clknet_3_5_0_io_wbs_clk),
    .X(clknet_leaf_74_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_io_wbs_clk (.A(clknet_3_5_0_io_wbs_clk),
    .X(clknet_leaf_75_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_io_wbs_clk (.A(clknet_3_5_0_io_wbs_clk),
    .X(clknet_leaf_76_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_io_wbs_clk (.A(clknet_3_5_0_io_wbs_clk),
    .X(clknet_leaf_77_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_io_wbs_clk (.A(clknet_opt_3_0_io_wbs_clk),
    .X(clknet_leaf_78_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_io_wbs_clk (.A(clknet_3_1_0_io_wbs_clk),
    .X(clknet_leaf_79_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_io_wbs_clk (.A(clknet_3_5_0_io_wbs_clk),
    .X(clknet_leaf_80_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_io_wbs_clk (.A(clknet_3_1_0_io_wbs_clk),
    .X(clknet_leaf_81_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_io_wbs_clk (.A(clknet_3_5_0_io_wbs_clk),
    .X(clknet_leaf_82_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_io_wbs_clk (.A(clknet_3_5_0_io_wbs_clk),
    .X(clknet_leaf_83_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_io_wbs_clk (.A(clknet_3_1_0_io_wbs_clk),
    .X(clknet_leaf_84_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_io_wbs_clk (.A(clknet_3_5_0_io_wbs_clk),
    .X(clknet_leaf_85_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_io_wbs_clk (.A(clknet_3_3_0_io_wbs_clk),
    .X(clknet_leaf_86_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_io_wbs_clk (.A(clknet_3_3_0_io_wbs_clk),
    .X(clknet_leaf_87_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_io_wbs_clk (.A(clknet_3_1_0_io_wbs_clk),
    .X(clknet_leaf_88_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_io_wbs_clk (.A(clknet_3_1_0_io_wbs_clk),
    .X(clknet_leaf_89_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_io_wbs_clk (.A(clknet_3_1_0_io_wbs_clk),
    .X(clknet_leaf_90_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_io_wbs_clk (.A(clknet_3_1_0_io_wbs_clk),
    .X(clknet_leaf_91_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_io_wbs_clk (.A(clknet_3_1_0_io_wbs_clk),
    .X(clknet_leaf_92_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_io_wbs_clk (.A(clknet_3_1_0_io_wbs_clk),
    .X(clknet_leaf_93_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_io_wbs_clk (.A(clknet_3_1_0_io_wbs_clk),
    .X(clknet_leaf_94_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_io_wbs_clk (.A(clknet_3_1_0_io_wbs_clk),
    .X(clknet_leaf_95_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_io_wbs_clk (.A(clknet_3_1_0_io_wbs_clk),
    .X(clknet_leaf_96_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_io_wbs_clk (.A(clknet_3_1_0_io_wbs_clk),
    .X(clknet_leaf_97_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_io_wbs_clk (.A(clknet_3_1_0_io_wbs_clk),
    .X(clknet_leaf_98_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_io_wbs_clk (.A(clknet_3_1_0_io_wbs_clk),
    .X(clknet_leaf_99_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_io_wbs_clk (.A(clknet_3_1_0_io_wbs_clk),
    .X(clknet_leaf_100_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_io_wbs_clk (.A(clknet_3_1_0_io_wbs_clk),
    .X(clknet_leaf_101_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_io_wbs_clk (.A(clknet_3_0_0_io_wbs_clk),
    .X(clknet_leaf_102_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_io_wbs_clk (.A(clknet_3_0_0_io_wbs_clk),
    .X(clknet_leaf_103_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_io_wbs_clk (.A(clknet_3_0_0_io_wbs_clk),
    .X(clknet_leaf_104_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_io_wbs_clk (.A(clknet_3_0_0_io_wbs_clk),
    .X(clknet_leaf_105_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_io_wbs_clk (.A(clknet_3_0_0_io_wbs_clk),
    .X(clknet_leaf_106_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_io_wbs_clk (.A(clknet_3_0_0_io_wbs_clk),
    .X(clknet_leaf_107_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_io_wbs_clk (.A(clknet_3_0_0_io_wbs_clk),
    .X(clknet_leaf_108_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_io_wbs_clk (.A(clknet_3_0_0_io_wbs_clk),
    .X(clknet_leaf_109_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_io_wbs_clk (.A(io_wbs_clk),
    .X(clknet_0_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0_io_wbs_clk (.A(clknet_0_io_wbs_clk),
    .X(clknet_1_0_0_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_1_io_wbs_clk (.A(clknet_1_0_0_io_wbs_clk),
    .X(clknet_1_0_1_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_0_io_wbs_clk (.A(clknet_0_io_wbs_clk),
    .X(clknet_1_1_0_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_1_io_wbs_clk (.A(clknet_1_1_0_io_wbs_clk),
    .X(clknet_1_1_1_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_io_wbs_clk (.A(clknet_1_0_1_io_wbs_clk),
    .X(clknet_2_0_0_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_io_wbs_clk (.A(clknet_1_0_1_io_wbs_clk),
    .X(clknet_2_1_0_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_io_wbs_clk (.A(clknet_1_1_1_io_wbs_clk),
    .X(clknet_2_2_0_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_io_wbs_clk (.A(clknet_1_1_1_io_wbs_clk),
    .X(clknet_2_3_0_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_io_wbs_clk (.A(clknet_2_0_0_io_wbs_clk),
    .X(clknet_3_0_0_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_io_wbs_clk (.A(clknet_2_0_0_io_wbs_clk),
    .X(clknet_3_1_0_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_io_wbs_clk (.A(clknet_2_1_0_io_wbs_clk),
    .X(clknet_3_2_0_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_io_wbs_clk (.A(clknet_2_1_0_io_wbs_clk),
    .X(clknet_3_3_0_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_io_wbs_clk (.A(clknet_2_2_0_io_wbs_clk),
    .X(clknet_3_4_0_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_io_wbs_clk (.A(clknet_2_2_0_io_wbs_clk),
    .X(clknet_3_5_0_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_io_wbs_clk (.A(clknet_2_3_0_io_wbs_clk),
    .X(clknet_3_6_0_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_io_wbs_clk (.A(clknet_2_3_0_io_wbs_clk),
    .X(clknet_3_7_0_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_0_io_wbs_clk (.A(clknet_3_0_0_io_wbs_clk),
    .X(clknet_opt_1_0_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_0_io_wbs_clk (.A(clknet_3_2_0_io_wbs_clk),
    .X(clknet_opt_2_0_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_3_0_io_wbs_clk (.A(clknet_3_5_0_io_wbs_clk),
    .X(clknet_opt_3_0_io_wbs_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_4_0_io_wbs_clk (.A(clknet_3_7_0_io_wbs_clk),
    .X(clknet_opt_4_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20201__D (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13741__B1_N (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13399__A (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20924__D (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10302__C1 (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10299__B1 (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10297__C1 (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10294__C1 (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10291__C1 (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10286__C1 (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10283__C1 (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10280__B1 (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10075__S (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20646__D (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17078__B1 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17072__A2 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17071__A (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13916__B (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13902__A2 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13861__A (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20137__RESET_B (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18426__C1 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18424__C1 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18422__C1 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18420__C1 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18418__C1 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18416__C1 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18414__C1 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18412__C1 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18410__C1 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20756__RESET_B (.DIODE(_00325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20773__RESET_B (.DIODE(_00341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20557__D (.DIODE(_00855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20567__D (.DIODE(_00865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17823__S (.DIODE(_01320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17820__S (.DIODE(_01320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17817__S (.DIODE(_01320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17814__S (.DIODE(_01320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17811__S (.DIODE(_01320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17808__S (.DIODE(_01320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17805__S (.DIODE(_01320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17802__S (.DIODE(_01320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17799__S (.DIODE(_01320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17796__S (.DIODE(_01320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18328__B1 (.DIODE(_01351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18107__A (.DIODE(_01351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18104__A (.DIODE(_01351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18101__A (.DIODE(_01351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17883__A (.DIODE(_01351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17839__A (.DIODE(_01351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18096__A2 (.DIODE(_01378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18094__B (.DIODE(_01378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18093__B (.DIODE(_01378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18091__A (.DIODE(_01378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17874__C (.DIODE(_01378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18103__A2_N (.DIODE(_01384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18100__A2_N (.DIODE(_01384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18098__A2 (.DIODE(_01384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18095__A2 (.DIODE(_01384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18089__A2 (.DIODE(_01384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17892__A (.DIODE(_01384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17884__B (.DIODE(_01384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17883__B (.DIODE(_01384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17880__B (.DIODE(_01384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18109__A2 (.DIODE(_01387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17914__B1 (.DIODE(_01387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17912__B1 (.DIODE(_01387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17908__B1 (.DIODE(_01387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17905__B1 (.DIODE(_01387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17902__A1 (.DIODE(_01387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17899__B1 (.DIODE(_01387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17895__C1 (.DIODE(_01387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17891__B1 (.DIODE(_01387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17886__A0 (.DIODE(_01387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18092__A2 (.DIODE(_01394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18086__A2 (.DIODE(_01394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18083__A2 (.DIODE(_01394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18080__A2 (.DIODE(_01394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18077__A2 (.DIODE(_01394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18074__A2 (.DIODE(_01394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18071__A2 (.DIODE(_01394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18068__A2 (.DIODE(_01394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18065__A2 (.DIODE(_01394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17896__A3 (.DIODE(_01394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17919__A (.DIODE(_01411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17922__D (.DIODE(_01413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17924__C (.DIODE(_01414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17924__D (.DIODE(_01415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17954__A_N (.DIODE(_01416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17936__C (.DIODE(_01416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17933__C (.DIODE(_01416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17931__B_N (.DIODE(_01416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17952__A1 (.DIODE(_01420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17932__B (.DIODE(_01420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17929__A (.DIODE(_01420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19065__A2 (.DIODE(_01427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18020__A2 (.DIODE(_01427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18017__A2 (.DIODE(_01427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18014__A2 (.DIODE(_01427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17982__A2 (.DIODE(_01427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17974__A2 (.DIODE(_01427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17967__A (.DIODE(_01427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17965__A2 (.DIODE(_01427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17960__A2 (.DIODE(_01427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17944__A2 (.DIODE(_01427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19414__A (.DIODE(_01429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19412__A (.DIODE(_01429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19407__A (.DIODE(_01429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17984__B1 (.DIODE(_01429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17981__B1 (.DIODE(_01429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17976__B1 (.DIODE(_01429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17973__B1 (.DIODE(_01429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17968__B1 (.DIODE(_01429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17938__A (.DIODE(_01429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18042__B1 (.DIODE(_01430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18038__B1 (.DIODE(_01430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18034__B1 (.DIODE(_01430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18030__B1 (.DIODE(_01430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18026__B1 (.DIODE(_01430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18022__B1 (.DIODE(_01430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17988__A (.DIODE(_01430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17964__B1 (.DIODE(_01430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17960__B1 (.DIODE(_01430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17944__B1 (.DIODE(_01430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17985__A2 (.DIODE(_01432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17983__A2 (.DIODE(_01432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17977__A2 (.DIODE(_01432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17975__A2 (.DIODE(_01432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17969__A2 (.DIODE(_01432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17966__A2 (.DIODE(_01432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17959__A2 (.DIODE(_01432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17943__A2 (.DIODE(_01432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18497__A (.DIODE(_01433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18482__A (.DIODE(_01433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18018__B (.DIODE(_01433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18015__B (.DIODE(_01433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18012__B (.DIODE(_01433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18009__B (.DIODE(_01433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18006__B (.DIODE(_01433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17963__A (.DIODE(_01433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17942__A (.DIODE(_01433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18003__B (.DIODE(_01434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18000__B (.DIODE(_01434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17997__B (.DIODE(_01434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17992__B (.DIODE(_01434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17989__B (.DIODE(_01434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17984__A2 (.DIODE(_01434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17976__A2 (.DIODE(_01434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17968__A2 (.DIODE(_01434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17959__B1 (.DIODE(_01434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17943__B1 (.DIODE(_01434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17944__C1 (.DIODE(_01435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17948__D (.DIODE(_01439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18042__A2 (.DIODE(_01444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18038__A2 (.DIODE(_01444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18034__A2 (.DIODE(_01444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18030__A2 (.DIODE(_01444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17995__A (.DIODE(_01444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17953__A (.DIODE(_01444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18041__A2 (.DIODE(_01446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18037__A2 (.DIODE(_01446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18033__A2 (.DIODE(_01446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18029__A2 (.DIODE(_01446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17996__A (.DIODE(_01446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17955__A (.DIODE(_01446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17960__C1 (.DIODE(_01450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19968__B (.DIODE(_01453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18041__B1 (.DIODE(_01453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18037__B1 (.DIODE(_01453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18033__B1 (.DIODE(_01453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18029__B1 (.DIODE(_01453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18025__B1 (.DIODE(_01453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18021__B1 (.DIODE(_01453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17981__A2 (.DIODE(_01453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17973__A2 (.DIODE(_01453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17964__A2 (.DIODE(_01453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18011__A2 (.DIODE(_01456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18008__A2 (.DIODE(_01456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18005__A2 (.DIODE(_01456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18002__A2 (.DIODE(_01456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17999__A2 (.DIODE(_01456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17994__A2 (.DIODE(_01456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17991__A2 (.DIODE(_01456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17987__A2 (.DIODE(_01456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17979__A2 (.DIODE(_01456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17971__A2 (.DIODE(_01456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18020__B1 (.DIODE(_01472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18017__B1 (.DIODE(_01472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18014__B1 (.DIODE(_01472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18011__B1 (.DIODE(_01472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18008__B1 (.DIODE(_01472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18005__B1 (.DIODE(_01472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18002__B1 (.DIODE(_01472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17999__B1 (.DIODE(_01472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17994__B1 (.DIODE(_01472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17991__B1 (.DIODE(_01472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18026__A2 (.DIODE(_01477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18022__A2 (.DIODE(_01477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18019__A2 (.DIODE(_01477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18016__A2 (.DIODE(_01477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18013__A2 (.DIODE(_01477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18010__A2 (.DIODE(_01477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18007__A2 (.DIODE(_01477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18004__A2 (.DIODE(_01477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18001__A2 (.DIODE(_01477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17998__A2 (.DIODE(_01477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18032__A (.DIODE(_01503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18035__A (.DIODE(_01504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18039__A (.DIODE(_01507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18043__A (.DIODE(_01510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18061__B (.DIODE(_01514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18059__B (.DIODE(_01514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18057__B (.DIODE(_01514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18055__B (.DIODE(_01514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18053__B (.DIODE(_01514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18051__B (.DIODE(_01514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18049__B (.DIODE(_01514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18047__B (.DIODE(_01514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18058__A (.DIODE(_01520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18060__A (.DIODE(_01521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18062__A (.DIODE(_01522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18140__A2 (.DIODE(_01554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18137__A2 (.DIODE(_01554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18134__A2 (.DIODE(_01554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18131__A2 (.DIODE(_01554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18128__A2 (.DIODE(_01554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18125__A2 (.DIODE(_01554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18122__A2 (.DIODE(_01554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18119__A2 (.DIODE(_01554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18116__A2 (.DIODE(_01554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18113__A2 (.DIODE(_01554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18140__C1 (.DIODE(_01556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18137__C1 (.DIODE(_01556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18134__C1 (.DIODE(_01556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18131__C1 (.DIODE(_01556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18128__C1 (.DIODE(_01556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18125__C1 (.DIODE(_01556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18122__C1 (.DIODE(_01556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18119__C1 (.DIODE(_01556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18116__C1 (.DIODE(_01556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18113__C1 (.DIODE(_01556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19932__A (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19896__A (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19865__A (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19828__A (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18885__A (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18429__A (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18333__B (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18320__A (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18210__A (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18164__A (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20097__A (.DIODE(_01589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20076__A (.DIODE(_01589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20052__A (.DIODE(_01589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19460__A (.DIODE(_01589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19427__A (.DIODE(_01589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19186__A (.DIODE(_01589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19165__A (.DIODE(_01589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19142__A (.DIODE(_01589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19109__A (.DIODE(_01589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18165__A (.DIODE(_01589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19049__A (.DIODE(_01590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19045__S (.DIODE(_01590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19043__S (.DIODE(_01590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18645__B1 (.DIODE(_01590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18640__B1 (.DIODE(_01590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18635__B1 (.DIODE(_01590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18205__A (.DIODE(_01590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18198__S (.DIODE(_01590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18196__S (.DIODE(_01590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18167__A (.DIODE(_01590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20044__A (.DIODE(_01591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20036__A (.DIODE(_01591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19232__B1 (.DIODE(_01591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19230__B1 (.DIODE(_01591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19223__B1 (.DIODE(_01591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19220__B1 (.DIODE(_01591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18406__A (.DIODE(_01591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18190__A (.DIODE(_01591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18179__A (.DIODE(_01591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18168__A (.DIODE(_01591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18178__A (.DIODE(_01592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18177__A (.DIODE(_01592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18176__A (.DIODE(_01592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18175__A (.DIODE(_01592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18174__A (.DIODE(_01592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18173__A (.DIODE(_01592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18172__A (.DIODE(_01592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18171__A (.DIODE(_01592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18170__A (.DIODE(_01592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18169__A (.DIODE(_01592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18189__A (.DIODE(_01593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18188__A (.DIODE(_01593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18187__A (.DIODE(_01593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18186__A (.DIODE(_01593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18185__A (.DIODE(_01593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18184__A (.DIODE(_01593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18183__A (.DIODE(_01593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18182__A (.DIODE(_01593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18181__A (.DIODE(_01593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18180__A (.DIODE(_01593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18204__A (.DIODE(_01594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18203__A (.DIODE(_01594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18202__A (.DIODE(_01594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18201__A (.DIODE(_01594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18200__A (.DIODE(_01594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18195__A (.DIODE(_01594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18194__A (.DIODE(_01594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18193__A (.DIODE(_01594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18192__A (.DIODE(_01594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18191__A (.DIODE(_01594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19034__A (.DIODE(_01597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19019__A (.DIODE(_01597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18478__A (.DIODE(_01597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18467__A (.DIODE(_01597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18389__A (.DIODE(_01597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18378__A (.DIODE(_01597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18367__A (.DIODE(_01597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18356__A (.DIODE(_01597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18345__A (.DIODE(_01597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18206__A (.DIODE(_01597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18344__A (.DIODE(_01598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18343__A (.DIODE(_01598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18342__A (.DIODE(_01598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18339__A (.DIODE(_01598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18338__A (.DIODE(_01598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18337__A (.DIODE(_01598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18336__A (.DIODE(_01598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18209__A (.DIODE(_01598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18208__A (.DIODE(_01598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18207__A (.DIODE(_01598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18853__A (.DIODE(_01599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18821__A (.DIODE(_01599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18784__A (.DIODE(_01599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18741__A (.DIODE(_01599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18709__A (.DIODE(_01599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18677__A (.DIODE(_01599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18311__A (.DIODE(_01599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18274__A (.DIODE(_01599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18236__A (.DIODE(_01599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18211__A (.DIODE(_01599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20136__C1 (.DIODE(_01600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20134__C1 (.DIODE(_01600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20132__C1 (.DIODE(_01600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20130__C1 (.DIODE(_01600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20128__C1 (.DIODE(_01600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20101__C1 (.DIODE(_01600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19780__C1 (.DIODE(_01600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19228__C1 (.DIODE(_01600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18234__A (.DIODE(_01600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18230__A (.DIODE(_01600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19887__A0 (.DIODE(_01601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19644__A0 (.DIODE(_01601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19592__A0 (.DIODE(_01601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19539__A0 (.DIODE(_01601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19138__A1 (.DIODE(_01601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18935__A0 (.DIODE(_01601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18831__A0 (.DIODE(_01601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18783__A1 (.DIODE(_01601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18678__A0 (.DIODE(_01601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18229__A0 (.DIODE(_01601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18492__B (.DIODE(_01602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18324__B (.DIODE(_01602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18215__A (.DIODE(_01602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19912__A (.DIODE(_01604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19564__A (.DIODE(_01604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19062__A (.DIODE(_01604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18754__A (.DIODE(_01604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18226__A (.DIODE(_01604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20102__C (.DIODE(_01605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19506__B (.DIODE(_01605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19191__B (.DIODE(_01605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19130__B (.DIODE(_01605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18650__B (.DIODE(_01605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18328__A1 (.DIODE(_01605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18327__B (.DIODE(_01605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18226__B (.DIODE(_01605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19506__C (.DIODE(_01607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18650__C (.DIODE(_01607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18481__A (.DIODE(_01607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18321__A (.DIODE(_01607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18226__C (.DIODE(_01607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18648__C (.DIODE(_01613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18225__D (.DIODE(_01613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19787__A0 (.DIODE(_01620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19647__A0 (.DIODE(_01620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19595__A0 (.DIODE(_01620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19542__A0 (.DIODE(_01620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19140__A1 (.DIODE(_01620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18938__A0 (.DIODE(_01620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18834__A0 (.DIODE(_01620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18785__A0 (.DIODE(_01620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18681__A0 (.DIODE(_01620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18233__A0 (.DIODE(_01620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18272__A (.DIODE(_01623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18269__A (.DIODE(_01623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18265__A (.DIODE(_01623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18262__A (.DIODE(_01623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18259__A (.DIODE(_01623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18255__A (.DIODE(_01623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18251__A (.DIODE(_01623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18247__A (.DIODE(_01623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18243__A (.DIODE(_01623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18239__A (.DIODE(_01623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19790__A0 (.DIODE(_01624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19650__A0 (.DIODE(_01624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19598__A0 (.DIODE(_01624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19545__A0 (.DIODE(_01624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19143__A1 (.DIODE(_01624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18942__A0 (.DIODE(_01624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18838__A0 (.DIODE(_01624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18788__A0 (.DIODE(_01624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18685__A0 (.DIODE(_01624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18238__A0 (.DIODE(_01624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19793__A0 (.DIODE(_01627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19654__A0 (.DIODE(_01627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19601__A0 (.DIODE(_01627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19549__A0 (.DIODE(_01627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19145__A1 (.DIODE(_01627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18945__A0 (.DIODE(_01627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18841__A0 (.DIODE(_01627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18791__A0 (.DIODE(_01627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18688__A0 (.DIODE(_01627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18242__A0 (.DIODE(_01627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19900__A0 (.DIODE(_01630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19797__A0 (.DIODE(_01630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19657__A0 (.DIODE(_01630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19552__A0 (.DIODE(_01630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19147__A1 (.DIODE(_01630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18948__A0 (.DIODE(_01630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18844__A0 (.DIODE(_01630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18794__A0 (.DIODE(_01630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18691__A0 (.DIODE(_01630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18246__A0 (.DIODE(_01630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19800__A0 (.DIODE(_01633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19660__A0 (.DIODE(_01633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19607__A0 (.DIODE(_01633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19555__A0 (.DIODE(_01633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19149__A1 (.DIODE(_01633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18952__A0 (.DIODE(_01633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18847__A0 (.DIODE(_01633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18798__A1 (.DIODE(_01633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18694__A0 (.DIODE(_01633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18250__A0 (.DIODE(_01633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19906__A0 (.DIODE(_01636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19803__A0 (.DIODE(_01636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19663__A0 (.DIODE(_01636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19610__A0 (.DIODE(_01636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19151__A1 (.DIODE(_01636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18955__A0 (.DIODE(_01636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18850__A0 (.DIODE(_01636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18799__A0 (.DIODE(_01636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18697__A0 (.DIODE(_01636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18254__A0 (.DIODE(_01636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19806__A0 (.DIODE(_01639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19666__A0 (.DIODE(_01639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19613__A0 (.DIODE(_01639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19561__A0 (.DIODE(_01639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19153__A1 (.DIODE(_01639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18958__A0 (.DIODE(_01639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18854__A0 (.DIODE(_01639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18803__A1 (.DIODE(_01639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18700__A0 (.DIODE(_01639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18258__A0 (.DIODE(_01639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18300__S (.DIODE(_01646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18296__S (.DIODE(_01646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18292__S (.DIODE(_01646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18288__S (.DIODE(_01646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18284__S (.DIODE(_01646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18281__S (.DIODE(_01646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18278__S (.DIODE(_01646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18275__S (.DIODE(_01646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18271__S (.DIODE(_01646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18268__S (.DIODE(_01646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18309__A (.DIODE(_01651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18305__A (.DIODE(_01651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18301__A (.DIODE(_01651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18297__A (.DIODE(_01651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18293__A (.DIODE(_01651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18289__A (.DIODE(_01651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18285__A (.DIODE(_01651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18282__A (.DIODE(_01651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18279__A (.DIODE(_01651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18276__A (.DIODE(_01651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20122__A1 (.DIODE(_01660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20109__A1 (.DIODE(_01660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20101__A1 (.DIODE(_01660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19780__A1 (.DIODE(_01660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19237__A1 (.DIODE(_01660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19231__A1 (.DIODE(_01660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19228__A1 (.DIODE(_01660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19174__A1 (.DIODE(_01660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18762__A1 (.DIODE(_01660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18288__A0 (.DIODE(_01660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20124__A1 (.DIODE(_01663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20115__A1 (.DIODE(_01663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19919__A1 (.DIODE(_01663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19239__A1 (.DIODE(_01663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19233__A1 (.DIODE(_01663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19176__A1 (.DIODE(_01663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18809__A0 (.DIODE(_01663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18763__A0 (.DIODE(_01663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18656__A0 (.DIODE(_01663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18292__A0 (.DIODE(_01663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20126__A1 (.DIODE(_01666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20111__A1 (.DIODE(_01666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19573__A0 (.DIODE(_01666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19521__A0 (.DIODE(_01666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19178__A1 (.DIODE(_01666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18916__A0 (.DIODE(_01666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18812__A0 (.DIODE(_01666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18766__A0 (.DIODE(_01666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18659__A0 (.DIODE(_01666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18296__A0 (.DIODE(_01666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20128__A1 (.DIODE(_01669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20113__A1 (.DIODE(_01669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19576__A0 (.DIODE(_01669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19524__A0 (.DIODE(_01669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19180__A1 (.DIODE(_01669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18920__A0 (.DIODE(_01669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18815__A0 (.DIODE(_01669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18769__A0 (.DIODE(_01669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18662__A0 (.DIODE(_01669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18300__A0 (.DIODE(_01669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20130__A1 (.DIODE(_01672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20117__A1 (.DIODE(_01672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19579__A0 (.DIODE(_01672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19527__A0 (.DIODE(_01672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19182__A1 (.DIODE(_01672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18923__A0 (.DIODE(_01672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18818__A0 (.DIODE(_01672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18772__A0 (.DIODE(_01672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18665__A0 (.DIODE(_01672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18304__A0 (.DIODE(_01672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20132__A1 (.DIODE(_01675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20107__A1 (.DIODE(_01675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19582__A0 (.DIODE(_01675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19530__A0 (.DIODE(_01675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19184__A1 (.DIODE(_01675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18926__A0 (.DIODE(_01675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18822__A0 (.DIODE(_01675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18775__A0 (.DIODE(_01675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18668__A0 (.DIODE(_01675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18308__A0 (.DIODE(_01675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18675__A (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18672__A (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18669__A (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18666__A (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18663__A (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18660__A (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18657__A (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18654__A (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18318__A (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18314__A (.DIODE(_01678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20134__A1 (.DIODE(_01679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19638__A0 (.DIODE(_01679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19586__A0 (.DIODE(_01679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19533__A0 (.DIODE(_01679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19187__A1 (.DIODE(_01679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18929__A0 (.DIODE(_01679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18825__A0 (.DIODE(_01679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18779__A1 (.DIODE(_01679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18671__A0 (.DIODE(_01679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18313__A0 (.DIODE(_01679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20136__A1 (.DIODE(_01682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19641__A0 (.DIODE(_01682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19589__A0 (.DIODE(_01682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19536__A0 (.DIODE(_01682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19189__A1 (.DIODE(_01682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18932__A0 (.DIODE(_01682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18828__A0 (.DIODE(_01682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18781__A1 (.DIODE(_01682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18674__A0 (.DIODE(_01682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18317__A0 (.DIODE(_01682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19488__A (.DIODE(_01685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19484__A (.DIODE(_01685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19480__A (.DIODE(_01685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19476__A (.DIODE(_01685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19419__A (.DIODE(_01685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19192__A (.DIODE(_01685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18574__A (.DIODE(_01685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18530__A (.DIODE(_01685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18517__A (.DIODE(_01685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18329__A (.DIODE(_01685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20102__D (.DIODE(_01686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19416__B (.DIODE(_01686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19225__B (.DIODE(_01686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19195__B (.DIODE(_01686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19069__B (.DIODE(_01686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19029__B (.DIODE(_01686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18500__B (.DIODE(_01686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18401__B (.DIODE(_01686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18332__B (.DIODE(_01686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18323__A (.DIODE(_01686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19414__B (.DIODE(_01690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18651__A (.DIODE(_01690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18497__B (.DIODE(_01690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18326__A (.DIODE(_01690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20101__A2 (.DIODE(_01691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19780__A2 (.DIODE(_01691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19779__A1 (.DIODE(_01691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19508__B (.DIODE(_01691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19507__A1 (.DIODE(_01691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19228__A2 (.DIODE(_01691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19218__C (.DIODE(_01691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19191__C (.DIODE(_01691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18328__A3 (.DIODE(_01691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18327__D (.DIODE(_01691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18355__A (.DIODE(_01700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18354__A (.DIODE(_01700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18353__A (.DIODE(_01700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18352__A (.DIODE(_01700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18351__A (.DIODE(_01700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18350__A (.DIODE(_01700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18349__A (.DIODE(_01700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18348__A (.DIODE(_01700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18347__A (.DIODE(_01700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18346__A (.DIODE(_01700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18388__A (.DIODE(_01703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18387__A (.DIODE(_01703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18386__A (.DIODE(_01703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18385__A (.DIODE(_01703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18384__A (.DIODE(_01703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18383__A (.DIODE(_01703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18382__A (.DIODE(_01703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18381__A (.DIODE(_01703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18380__A (.DIODE(_01703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18379__A (.DIODE(_01703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18466__A (.DIODE(_01704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18465__A (.DIODE(_01704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18464__A (.DIODE(_01704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18463__A (.DIODE(_01704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18462__A (.DIODE(_01704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18461__A (.DIODE(_01704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18393__A (.DIODE(_01704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18392__A (.DIODE(_01704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18391__A (.DIODE(_01704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18390__A (.DIODE(_01704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19772__A (.DIODE(_01706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19767__A (.DIODE(_01706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19407__C (.DIODE(_01706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19201__A (.DIODE(_01706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19198__A (.DIODE(_01706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19079__A (.DIODE(_01706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19057__A (.DIODE(_01706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18482__C (.DIODE(_01706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18396__B (.DIODE(_01706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18459__B1 (.DIODE(_01707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18457__B1 (.DIODE(_01707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18455__B1 (.DIODE(_01707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18452__B1 (.DIODE(_01707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18427__A (.DIODE(_01707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18397__A (.DIODE(_01707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20100__A2 (.DIODE(_01709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20040__C (.DIODE(_01709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20039__B (.DIODE(_01709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19227__A2 (.DIODE(_01709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19203__A2 (.DIODE(_01709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19190__A2 (.DIODE(_01709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18400__C (.DIODE(_01709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18399__B (.DIODE(_01709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18459__A2 (.DIODE(_01710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18457__A2 (.DIODE(_01710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18455__A2 (.DIODE(_01710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18433__A (.DIODE(_01710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18408__A (.DIODE(_01710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18404__A2 (.DIODE(_01710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20041__B (.DIODE(_01713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20037__B (.DIODE(_01713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19416__C (.DIODE(_01713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19069__C (.DIODE(_01713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18500__C (.DIODE(_01713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18403__B (.DIODE(_01713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18460__A2 (.DIODE(_01714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18458__A2 (.DIODE(_01714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18456__A2 (.DIODE(_01714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18432__A (.DIODE(_01714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18407__A (.DIODE(_01714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18404__C1 (.DIODE(_01714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18431__A2 (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18426__A2 (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18424__A2 (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18422__A2 (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18420__A2 (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18418__A2 (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18416__A2 (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18414__A2 (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18412__A2 (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18410__A2 (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19509__A (.DIODE(_01730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19504__A (.DIODE(_01730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19500__A (.DIODE(_01730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19496__A (.DIODE(_01730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19492__A (.DIODE(_01730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19070__A (.DIODE(_01730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18616__A (.DIODE(_01730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18544__A (.DIODE(_01730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18453__A (.DIODE(_01730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18430__A (.DIODE(_01730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18540__C1 (.DIODE(_01744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18535__C1 (.DIODE(_01744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18526__C1 (.DIODE(_01744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18522__C1 (.DIODE(_01744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18512__C1 (.DIODE(_01744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18504__C1 (.DIODE(_01744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18460__C1 (.DIODE(_01744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18458__C1 (.DIODE(_01744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18456__C1 (.DIODE(_01744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18454__C1 (.DIODE(_01744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18477__A (.DIODE(_01748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18476__A (.DIODE(_01748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18475__A (.DIODE(_01748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18474__A (.DIODE(_01748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18473__A (.DIODE(_01748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18472__A (.DIODE(_01748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18471__A (.DIODE(_01748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18470__A (.DIODE(_01748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18469__A (.DIODE(_01748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18468__A (.DIODE(_01748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19018__A (.DIODE(_01749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19017__A (.DIODE(_01749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19016__A (.DIODE(_01749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19015__A (.DIODE(_01749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19014__A (.DIODE(_01749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19013__A (.DIODE(_01749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19012__A (.DIODE(_01749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19011__A (.DIODE(_01749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18480__A (.DIODE(_01749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18479__A (.DIODE(_01749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18571__B (.DIODE(_01751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18527__B (.DIODE(_01751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18513__B (.DIODE(_01751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18505__A (.DIODE(_01751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18483__A (.DIODE(_01751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18631__A2 (.DIODE(_01752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18628__A2 (.DIODE(_01752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18620__A2 (.DIODE(_01752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18617__A2 (.DIODE(_01752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18613__A2 (.DIODE(_01752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18605__A2 (.DIODE(_01752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18579__A2 (.DIODE(_01752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18570__A2 (.DIODE(_01752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18566__A2 (.DIODE(_01752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18484__A (.DIODE(_01752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18646__A2 (.DIODE(_01753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18641__A2 (.DIODE(_01753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18636__A2 (.DIODE(_01753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18625__A2 (.DIODE(_01753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18610__A2 (.DIODE(_01753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18602__A2 (.DIODE(_01753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18597__A2 (.DIODE(_01753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18592__A2 (.DIODE(_01753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18587__A2 (.DIODE(_01753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18504__A2 (.DIODE(_01753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18500__A (.DIODE(_01754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18495__A (.DIODE(_01754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18491__B1 (.DIODE(_01754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18488__A (.DIODE(_01754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19061__C1 (.DIODE(_01755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18491__A1 (.DIODE(_01755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18487__C (.DIODE(_01755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19781__A (.DIODE(_01756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19616__B (.DIODE(_01756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19072__B (.DIODE(_01756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19064__B (.DIODE(_01756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18908__B (.DIODE(_01756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18488__B (.DIODE(_01756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18572__B1 (.DIODE(_01757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18558__A (.DIODE(_01757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18528__B1 (.DIODE(_01757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18515__B1 (.DIODE(_01757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18489__A (.DIODE(_01757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18643__B (.DIODE(_01758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18638__B (.DIODE(_01758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18633__B (.DIODE(_01758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18629__B1 (.DIODE(_01758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18626__B1 (.DIODE(_01758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18618__B1 (.DIODE(_01758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18614__B1 (.DIODE(_01758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18611__B1 (.DIODE(_01758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18603__B1 (.DIODE(_01758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18490__A (.DIODE(_01758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18556__A2 (.DIODE(_01759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18552__A2 (.DIODE(_01759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18548__A2 (.DIODE(_01759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18543__A2 (.DIODE(_01759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18539__A2 (.DIODE(_01759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18534__A2 (.DIODE(_01759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18525__A2 (.DIODE(_01759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18521__A2 (.DIODE(_01759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18511__A2 (.DIODE(_01759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18503__A2 (.DIODE(_01759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18577__A2 (.DIODE(_01760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18573__A2 (.DIODE(_01760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18568__A2 (.DIODE(_01760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18564__A2 (.DIODE(_01760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18529__A2 (.DIODE(_01760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18516__A2 (.DIODE(_01760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18508__A (.DIODE(_01760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18496__A2 (.DIODE(_01760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19200__B (.DIODE(_01761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18493__B (.DIODE(_01761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19859__A (.DIODE(_01762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19511__B (.DIODE(_01762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18804__A (.DIODE(_01762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18494__A (.DIODE(_01762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20120__A (.DIODE(_01763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20118__A (.DIODE(_01763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19768__B (.DIODE(_01763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19415__B (.DIODE(_01763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19235__A (.DIODE(_01763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19234__A (.DIODE(_01763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19202__B (.DIODE(_01763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19074__B (.DIODE(_01763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19067__A3 (.DIODE(_01763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18495__B (.DIODE(_01763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18582__A (.DIODE(_01764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18573__B1 (.DIODE(_01764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18514__A (.DIODE(_01764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18509__A (.DIODE(_01764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18496__B1 (.DIODE(_01764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18572__A2 (.DIODE(_01766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18528__A2 (.DIODE(_01766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18515__A2 (.DIODE(_01766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18506__A (.DIODE(_01766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18498__A (.DIODE(_01766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18629__A2 (.DIODE(_01767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18626__A2 (.DIODE(_01767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18618__A2 (.DIODE(_01767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18614__A2 (.DIODE(_01767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18611__A2 (.DIODE(_01767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18603__A2 (.DIODE(_01767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18576__A2 (.DIODE(_01767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18567__A2 (.DIODE(_01767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18563__A2 (.DIODE(_01767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18499__A (.DIODE(_01767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18642__B (.DIODE(_01768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18637__B (.DIODE(_01768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18632__B (.DIODE(_01768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18621__B (.DIODE(_01768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18606__B (.DIODE(_01768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18598__B (.DIODE(_01768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18593__B (.DIODE(_01768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18588__B (.DIODE(_01768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18580__B (.DIODE(_01768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18502__A2 (.DIODE(_01768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18572__C1 (.DIODE(_01769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18536__A (.DIODE(_01769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18528__C1 (.DIODE(_01769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18515__C1 (.DIODE(_01769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18501__A (.DIODE(_01769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18644__B1 (.DIODE(_01770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18639__B1 (.DIODE(_01770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18634__B1 (.DIODE(_01770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18623__B1 (.DIODE(_01770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18608__B1 (.DIODE(_01770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18532__B1 (.DIODE(_01770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18523__B1 (.DIODE(_01770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18519__B1 (.DIODE(_01770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18507__B1 (.DIODE(_01770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18502__B1 (.DIODE(_01770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18559__A2 (.DIODE(_01774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18554__A2 (.DIODE(_01774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18550__A2 (.DIODE(_01774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18546__A2 (.DIODE(_01774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18541__A2 (.DIODE(_01774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18537__A2 (.DIODE(_01774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18532__A2 (.DIODE(_01774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18523__A2 (.DIODE(_01774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18519__A2 (.DIODE(_01774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18507__A2 (.DIODE(_01774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18560__A2 (.DIODE(_01776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18555__A2 (.DIODE(_01776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18551__A2 (.DIODE(_01776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18547__A2 (.DIODE(_01776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18542__A2 (.DIODE(_01776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18538__A2 (.DIODE(_01776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18533__A2 (.DIODE(_01776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18524__A2 (.DIODE(_01776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18520__A2 (.DIODE(_01776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18510__A2 (.DIODE(_01776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18644__A2 (.DIODE(_01777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18639__A2 (.DIODE(_01777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18634__A2 (.DIODE(_01777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18623__A2 (.DIODE(_01777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18608__A2 (.DIODE(_01777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18538__B1 (.DIODE(_01777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18533__B1 (.DIODE(_01777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18524__B1 (.DIODE(_01777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18520__B1 (.DIODE(_01777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18510__B1 (.DIODE(_01777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18512__B1 (.DIODE(_01779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18577__B1 (.DIODE(_01781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18568__B1 (.DIODE(_01781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18564__B1 (.DIODE(_01781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18560__B1 (.DIODE(_01781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18555__B1 (.DIODE(_01781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18551__B1 (.DIODE(_01781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18547__B1 (.DIODE(_01781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18542__B1 (.DIODE(_01781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18529__B1 (.DIODE(_01781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18516__B1 (.DIODE(_01781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18517__C (.DIODE(_01783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18530__C (.DIODE(_01793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18583__A (.DIODE(_01798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18576__B1 (.DIODE(_01798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18567__B1 (.DIODE(_01798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18563__B1 (.DIODE(_01798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18559__B1 (.DIODE(_01798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18554__B1 (.DIODE(_01798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18550__B1 (.DIODE(_01798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18546__B1 (.DIODE(_01798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18541__B1 (.DIODE(_01798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18537__B1 (.DIODE(_01798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18613__C1 (.DIODE(_01805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18605__C1 (.DIODE(_01805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18579__C1 (.DIODE(_01805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18570__C1 (.DIODE(_01805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18566__C1 (.DIODE(_01805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18562__C1 (.DIODE(_01805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18557__C1 (.DIODE(_01805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18553__C1 (.DIODE(_01805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18549__C1 (.DIODE(_01805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18545__C1 (.DIODE(_01805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18549__B1 (.DIODE(_01808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18553__B1 (.DIODE(_01811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18622__B (.DIODE(_01815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18607__B (.DIODE(_01815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18599__B (.DIODE(_01815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18594__B (.DIODE(_01815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18589__B (.DIODE(_01815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18581__B (.DIODE(_01815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18578__A2 (.DIODE(_01815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18569__A2 (.DIODE(_01815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18565__A2 (.DIODE(_01815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18561__A2 (.DIODE(_01815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18562__B1 (.DIODE(_01818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18574__C (.DIODE(_01827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18630__A2 (.DIODE(_01834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18627__A2 (.DIODE(_01834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18619__A2 (.DIODE(_01834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18615__A2 (.DIODE(_01834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18612__A2 (.DIODE(_01834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18604__A2 (.DIODE(_01834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18600__A2 (.DIODE(_01834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18595__A2 (.DIODE(_01834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18590__A2 (.DIODE(_01834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18584__A2 (.DIODE(_01834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18630__C1 (.DIODE(_01835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18627__C1 (.DIODE(_01835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18619__C1 (.DIODE(_01835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18615__C1 (.DIODE(_01835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18612__C1 (.DIODE(_01835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18604__C1 (.DIODE(_01835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18600__B1 (.DIODE(_01835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18595__B1 (.DIODE(_01835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18590__B1 (.DIODE(_01835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18584__B1 (.DIODE(_01835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19836__A (.DIODE(_01837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19784__A (.DIODE(_01837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19605__A (.DIODE(_01837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19559__A (.DIODE(_01837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18624__B1 (.DIODE(_01837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18609__B1 (.DIODE(_01837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18601__B1 (.DIODE(_01837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18596__B1 (.DIODE(_01837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18591__B1 (.DIODE(_01837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18586__B1 (.DIODE(_01837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18605__B1 (.DIODE(_01852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18613__B1 (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18803__C1 (.DIODE(_01861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18798__C1 (.DIODE(_01861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18783__C1 (.DIODE(_01861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18781__C1 (.DIODE(_01861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18779__C1 (.DIODE(_01861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18762__C1 (.DIODE(_01861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18631__C1 (.DIODE(_01861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18628__C1 (.DIODE(_01861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18620__C1 (.DIODE(_01861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18617__C1 (.DIODE(_01861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19915__A0 (.DIODE(_01884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19862__A0 (.DIODE(_01884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19835__A0 (.DIODE(_01884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19619__A0 (.DIODE(_01884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19567__A0 (.DIODE(_01884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19514__A0 (.DIODE(_01884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19508__A (.DIODE(_01884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18910__A0 (.DIODE(_01884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18806__A0 (.DIODE(_01884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18653__A0 (.DIODE(_01884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18908__C (.DIODE(_01887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18804__B (.DIODE(_01887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18755__B (.DIODE(_01887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18651__B (.DIODE(_01887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18751__S (.DIODE(_01888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18748__S (.DIODE(_01888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18716__A (.DIODE(_01888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18684__A (.DIODE(_01888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18652__A (.DIODE(_01888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18681__S (.DIODE(_01889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18678__S (.DIODE(_01889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18674__S (.DIODE(_01889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18671__S (.DIODE(_01889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18668__S (.DIODE(_01889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18665__S (.DIODE(_01889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18662__S (.DIODE(_01889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18659__S (.DIODE(_01889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18656__S (.DIODE(_01889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18653__S (.DIODE(_01889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18707__A (.DIODE(_01906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18704__A (.DIODE(_01906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18701__A (.DIODE(_01906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18698__A (.DIODE(_01906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18695__A (.DIODE(_01906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18692__A (.DIODE(_01906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18689__A (.DIODE(_01906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18686__A (.DIODE(_01906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18682__A (.DIODE(_01906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18679__A (.DIODE(_01906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18713__S (.DIODE(_01911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18710__S (.DIODE(_01911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18706__S (.DIODE(_01911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18703__S (.DIODE(_01911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18700__S (.DIODE(_01911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18697__S (.DIODE(_01911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18694__S (.DIODE(_01911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18691__S (.DIODE(_01911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18688__S (.DIODE(_01911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18685__S (.DIODE(_01911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18739__A (.DIODE(_01928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18736__A (.DIODE(_01928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18733__A (.DIODE(_01928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18730__A (.DIODE(_01928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18727__A (.DIODE(_01928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18724__A (.DIODE(_01928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18721__A (.DIODE(_01928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18718__A (.DIODE(_01928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18714__A (.DIODE(_01928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18711__A (.DIODE(_01928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18745__S (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18742__S (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18738__S (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18735__S (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18732__S (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18729__S (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18726__S (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18723__S (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18720__S (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18717__S (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18776__A (.DIODE(_01950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18773__A (.DIODE(_01950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18770__A (.DIODE(_01950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18767__A (.DIODE(_01950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18764__A (.DIODE(_01950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18758__A (.DIODE(_01950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18752__A (.DIODE(_01950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18749__A (.DIODE(_01950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18746__A (.DIODE(_01950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18743__A (.DIODE(_01950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20105__A (.DIODE(_01959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20103__A (.DIODE(_01959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19770__B (.DIODE(_01959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19412__B (.DIODE(_01959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19411__B (.DIODE(_01959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19229__A (.DIODE(_01959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19218__B (.DIODE(_01959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19130__A (.DIODE(_01959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19076__B (.DIODE(_01959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18755__A (.DIODE(_01959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18799__S (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18794__S (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18791__S (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18788__S (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18756__A (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18802__B (.DIODE(_01961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18797__B (.DIODE(_01961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18785__S (.DIODE(_01961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18775__S (.DIODE(_01961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18772__S (.DIODE(_01961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18769__S (.DIODE(_01961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18766__S (.DIODE(_01961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18763__S (.DIODE(_01961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18760__A (.DIODE(_01961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18757__S (.DIODE(_01961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18819__A (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18816__A (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18813__A (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18810__A (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18807__A (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18800__A (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18795__A (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18792__A (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18789__A (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18786__A (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18905__S (.DIODE(_01992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18902__S (.DIODE(_01992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18869__A (.DIODE(_01992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18837__A (.DIODE(_01992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18805__A (.DIODE(_01992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18834__S (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18831__S (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18828__S (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18825__S (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18822__S (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18818__S (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18815__S (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18812__S (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18809__S (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18806__S (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18851__A (.DIODE(_02004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18848__A (.DIODE(_02004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18845__A (.DIODE(_02004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18842__A (.DIODE(_02004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18839__A (.DIODE(_02004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18835__A (.DIODE(_02004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18832__A (.DIODE(_02004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18829__A (.DIODE(_02004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18826__A (.DIODE(_02004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18823__A (.DIODE(_02004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18866__S (.DIODE(_02015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18863__S (.DIODE(_02015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18860__S (.DIODE(_02015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18857__S (.DIODE(_02015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18854__S (.DIODE(_02015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18850__S (.DIODE(_02015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18847__S (.DIODE(_02015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18844__S (.DIODE(_02015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18841__S (.DIODE(_02015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18838__S (.DIODE(_02015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18883__A (.DIODE(_02026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18880__A (.DIODE(_02026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18877__A (.DIODE(_02026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18874__A (.DIODE(_02026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18871__A (.DIODE(_02026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18867__A (.DIODE(_02026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18864__A (.DIODE(_02026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18861__A (.DIODE(_02026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18858__A (.DIODE(_02026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18855__A (.DIODE(_02026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18899__S (.DIODE(_02037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18896__S (.DIODE(_02037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18893__S (.DIODE(_02037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18890__S (.DIODE(_02037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18887__S (.DIODE(_02037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18882__S (.DIODE(_02037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18879__S (.DIODE(_02037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18876__S (.DIODE(_02037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18873__S (.DIODE(_02037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18870__S (.DIODE(_02037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19796__A (.DIODE(_02048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19653__A (.DIODE(_02048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19622__A (.DIODE(_02048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19585__A (.DIODE(_02048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19548__A (.DIODE(_02048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19517__A (.DIODE(_02048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18983__A (.DIODE(_02048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18951__A (.DIODE(_02048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18919__A (.DIODE(_02048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18886__A (.DIODE(_02048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18917__A (.DIODE(_02049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18914__A (.DIODE(_02049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18911__A (.DIODE(_02049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18906__A (.DIODE(_02049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18903__A (.DIODE(_02049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18900__A (.DIODE(_02049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18897__A (.DIODE(_02049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18894__A (.DIODE(_02049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18891__A (.DIODE(_02049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18888__A (.DIODE(_02049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19008__S (.DIODE(_02064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19005__S (.DIODE(_02064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18973__A (.DIODE(_02064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18941__A (.DIODE(_02064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18909__A (.DIODE(_02064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18938__S (.DIODE(_02065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18935__S (.DIODE(_02065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18932__S (.DIODE(_02065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18929__S (.DIODE(_02065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18926__S (.DIODE(_02065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18923__S (.DIODE(_02065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18920__S (.DIODE(_02065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18916__S (.DIODE(_02065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18913__S (.DIODE(_02065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18910__S (.DIODE(_02065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18949__A (.DIODE(_02072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18946__A (.DIODE(_02072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18943__A (.DIODE(_02072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18939__A (.DIODE(_02072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18936__A (.DIODE(_02072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18933__A (.DIODE(_02072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18930__A (.DIODE(_02072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18927__A (.DIODE(_02072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18924__A (.DIODE(_02072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18921__A (.DIODE(_02072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18970__S (.DIODE(_02087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18967__S (.DIODE(_02087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18964__S (.DIODE(_02087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18961__S (.DIODE(_02087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18958__S (.DIODE(_02087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18955__S (.DIODE(_02087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18952__S (.DIODE(_02087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18948__S (.DIODE(_02087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18945__S (.DIODE(_02087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18942__S (.DIODE(_02087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18981__A (.DIODE(_02094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18978__A (.DIODE(_02094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18975__A (.DIODE(_02094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18971__A (.DIODE(_02094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18968__A (.DIODE(_02094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18965__A (.DIODE(_02094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18962__A (.DIODE(_02094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18959__A (.DIODE(_02094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18956__A (.DIODE(_02094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18953__A (.DIODE(_02094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19002__S (.DIODE(_02109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18999__S (.DIODE(_02109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18996__S (.DIODE(_02109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18993__S (.DIODE(_02109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18990__S (.DIODE(_02109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18987__S (.DIODE(_02109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18984__S (.DIODE(_02109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18980__S (.DIODE(_02109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18977__S (.DIODE(_02109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18974__S (.DIODE(_02109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19515__A (.DIODE(_02116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19009__A (.DIODE(_02116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19006__A (.DIODE(_02116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19003__A (.DIODE(_02116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19000__A (.DIODE(_02116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18997__A (.DIODE(_02116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18994__A (.DIODE(_02116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18991__A (.DIODE(_02116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18988__A (.DIODE(_02116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18985__A (.DIODE(_02116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19033__A (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19032__A (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19027__A (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19026__A (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19025__A (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19024__A (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19023__A (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19022__A (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19021__A (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19020__A (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19048__A (.DIODE(_02139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19047__A (.DIODE(_02139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19042__A (.DIODE(_02139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19041__A (.DIODE(_02139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19040__A (.DIODE(_02139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19039__A (.DIODE(_02139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19038__A (.DIODE(_02139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19037__A (.DIODE(_02139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19036__A (.DIODE(_02139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19035__A (.DIODE(_02139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19335__A (.DIODE(_02142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19324__A (.DIODE(_02142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19313__A (.DIODE(_02142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19302__A (.DIODE(_02142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19291__A (.DIODE(_02142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19280__A (.DIODE(_02142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19269__A (.DIODE(_02142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19255__A (.DIODE(_02142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19244__A (.DIODE(_02142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19050__A (.DIODE(_02142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19067__A1 (.DIODE(_02153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19120__A2 (.DIODE(_02158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19117__A2 (.DIODE(_02158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19104__A2 (.DIODE(_02158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19098__A2 (.DIODE(_02158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19092__A2 (.DIODE(_02158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19089__A2 (.DIODE(_02158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19083__A2 (.DIODE(_02158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19073__A (.DIODE(_02158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19123__A2 (.DIODE(_02160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19114__A2 (.DIODE(_02160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19111__A2 (.DIODE(_02160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19107__A2 (.DIODE(_02160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19101__A2 (.DIODE(_02160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19075__A (.DIODE(_02160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19123__B1 (.DIODE(_02162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19114__B1 (.DIODE(_02162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19111__B1 (.DIODE(_02162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19107__B1 (.DIODE(_02162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19101__B1 (.DIODE(_02162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19077__A (.DIODE(_02162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19121__B1 (.DIODE(_02165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19118__B1 (.DIODE(_02165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19105__B1 (.DIODE(_02165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19099__B1 (.DIODE(_02165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19093__B1 (.DIODE(_02165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19090__B1 (.DIODE(_02165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19084__B1 (.DIODE(_02165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19080__A (.DIODE(_02165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19094__B1 (.DIODE(_02175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19097__B1 (.DIODE(_02177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19100__B1 (.DIODE(_02179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19106__B1 (.DIODE(_02183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19140__C1 (.DIODE(_02186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19138__C1 (.DIODE(_02186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19129__C1 (.DIODE(_02186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19127__C1 (.DIODE(_02186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19125__C1 (.DIODE(_02186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19122__C1 (.DIODE(_02186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19119__C1 (.DIODE(_02186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19116__C1 (.DIODE(_02186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19113__C1 (.DIODE(_02186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19110__C1 (.DIODE(_02186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20100__A1 (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20099__A (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19778__C (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19227__A1 (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19226__A (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19190__A1 (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19135__B (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19185__B (.DIODE(_02204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19183__B (.DIODE(_02204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19181__B (.DIODE(_02204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19159__A (.DIODE(_02204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19136__A (.DIODE(_02204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19163__C1 (.DIODE(_02209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19161__C1 (.DIODE(_02209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19157__C1 (.DIODE(_02209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19155__C1 (.DIODE(_02209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19153__C1 (.DIODE(_02209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19151__C1 (.DIODE(_02209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19149__C1 (.DIODE(_02209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19147__C1 (.DIODE(_02209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19145__C1 (.DIODE(_02209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19143__C1 (.DIODE(_02209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19180__A2 (.DIODE(_02217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19178__A2 (.DIODE(_02217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19176__A2 (.DIODE(_02217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19174__A2 (.DIODE(_02217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19172__A2 (.DIODE(_02217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19170__A2 (.DIODE(_02217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19168__A2 (.DIODE(_02217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19166__A2 (.DIODE(_02217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19163__A2 (.DIODE(_02217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19161__A2 (.DIODE(_02217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19179__B (.DIODE(_02218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19177__B (.DIODE(_02218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19175__B (.DIODE(_02218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19173__B (.DIODE(_02218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19171__B (.DIODE(_02218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19169__B (.DIODE(_02218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19167__B (.DIODE(_02218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19164__B (.DIODE(_02218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19162__B (.DIODE(_02218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19160__B (.DIODE(_02218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19184__C1 (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19182__C1 (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19180__C1 (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19178__C1 (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19176__C1 (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19174__C1 (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19172__C1 (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19170__C1 (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19168__C1 (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19166__C1 (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19239__C1 (.DIODE(_02233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19237__C1 (.DIODE(_02233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19216__C1 (.DIODE(_02233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19214__C1 (.DIODE(_02233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19212__C1 (.DIODE(_02233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19210__C1 (.DIODE(_02233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19208__C1 (.DIODE(_02233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19206__C1 (.DIODE(_02233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19189__C1 (.DIODE(_02233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19187__C1 (.DIODE(_02233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19218__A_N (.DIODE(_02238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19203__A1 (.DIODE(_02238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19202__A (.DIODE(_02238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19200__A (.DIODE(_02238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19195__A (.DIODE(_02238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20100__A3 (.DIODE(_02239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20099__B (.DIODE(_02239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19201__B (.DIODE(_02239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19198__B (.DIODE(_02239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19196__C (.DIODE(_02239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19770__A (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19768__A (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19225__A (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19772__B (.DIODE(_02260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19767__B (.DIODE(_02260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19676__C (.DIODE(_02260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19227__A3 (.DIODE(_02260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19226__B (.DIODE(_02260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19268__A (.DIODE(_02271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19267__A (.DIODE(_02271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19266__A (.DIODE(_02271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19262__A (.DIODE(_02271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19261__A (.DIODE(_02271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19260__A (.DIODE(_02271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19259__A (.DIODE(_02271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19258__A (.DIODE(_02271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19257__A (.DIODE(_02271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19256__A (.DIODE(_02271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19290__A (.DIODE(_02275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19289__A (.DIODE(_02275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19288__A (.DIODE(_02275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19287__A (.DIODE(_02275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19286__A (.DIODE(_02275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19285__A (.DIODE(_02275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19284__A (.DIODE(_02275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19283__A (.DIODE(_02275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19282__A (.DIODE(_02275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19281__A (.DIODE(_02275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19312__A (.DIODE(_02277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19311__A (.DIODE(_02277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19310__A (.DIODE(_02277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19309__A (.DIODE(_02277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19308__A (.DIODE(_02277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19307__A (.DIODE(_02277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19306__A (.DIODE(_02277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19305__A (.DIODE(_02277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19304__A (.DIODE(_02277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19303__A (.DIODE(_02277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19323__A (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19322__A (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19321__A (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19320__A (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19319__A (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19318__A (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19317__A (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19316__A (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19315__A (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19314__A (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19334__A (.DIODE(_02279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19333__A (.DIODE(_02279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19332__A (.DIODE(_02279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19331__A (.DIODE(_02279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19330__A (.DIODE(_02279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19329__A (.DIODE(_02279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19328__A (.DIODE(_02279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19327__A (.DIODE(_02279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19326__A (.DIODE(_02279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19325__A (.DIODE(_02279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19345__A (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19344__A (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19343__A (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19342__A (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19341__A (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19340__A (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19339__A (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19338__A (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19337__A (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19336__A (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19716__A (.DIODE(_02281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19705__A (.DIODE(_02281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19694__A (.DIODE(_02281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19683__A (.DIODE(_02281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19402__A (.DIODE(_02281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19391__A (.DIODE(_02281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19380__A (.DIODE(_02281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19369__A (.DIODE(_02281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19358__A (.DIODE(_02281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19347__A (.DIODE(_02281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19357__A (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19356__A (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19355__A (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19354__A (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19353__A (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19352__A (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19351__A (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19350__A (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19349__A (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19348__A (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19368__A (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19367__A (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19366__A (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19365__A (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19364__A (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19363__A (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19362__A (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19361__A (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19360__A (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19359__A (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19390__A (.DIODE(_02285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19389__A (.DIODE(_02285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19388__A (.DIODE(_02285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19387__A (.DIODE(_02285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19386__A (.DIODE(_02285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19385__A (.DIODE(_02285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19384__A (.DIODE(_02285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19383__A (.DIODE(_02285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19382__A (.DIODE(_02285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19381__A (.DIODE(_02285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19401__A (.DIODE(_02286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19400__A (.DIODE(_02286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19399__A (.DIODE(_02286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19398__A (.DIODE(_02286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19397__A (.DIODE(_02286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19396__A (.DIODE(_02286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19395__A (.DIODE(_02286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19394__A (.DIODE(_02286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19393__A (.DIODE(_02286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19392__A (.DIODE(_02286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19682__A (.DIODE(_02287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19681__A (.DIODE(_02287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19680__A (.DIODE(_02287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19679__A (.DIODE(_02287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19678__A (.DIODE(_02287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19675__A (.DIODE(_02287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19406__A (.DIODE(_02287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19405__A (.DIODE(_02287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19404__A (.DIODE(_02287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19403__A (.DIODE(_02287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19482__B (.DIODE(_02289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19478__B (.DIODE(_02289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19474__B (.DIODE(_02289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19473__A2 (.DIODE(_02289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19470__A2 (.DIODE(_02289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19467__A2 (.DIODE(_02289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19464__A2 (.DIODE(_02289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19461__A2 (.DIODE(_02289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19421__A (.DIODE(_02289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19409__B (.DIODE(_02289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19471__A2 (.DIODE(_02292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19468__A2 (.DIODE(_02292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19462__A2 (.DIODE(_02292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19449__A2 (.DIODE(_02292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19434__A2 (.DIODE(_02292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19422__A (.DIODE(_02292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19418__A2 (.DIODE(_02292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19503__A2 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19499__A2 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19495__A2 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19446__A2 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19443__A2 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19440__A2 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19437__A2 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19429__A2 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19425__A2 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19418__B1 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19466__A2 (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19459__A2 (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19456__A2 (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19453__A2 (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19447__A2 (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19444__A2 (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19441__A2 (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19438__A2 (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19430__A2 (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19426__A2 (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19455__B1 (.DIODE(_02303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19452__B1 (.DIODE(_02303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19449__B1 (.DIODE(_02303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19446__B1 (.DIODE(_02303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19443__B1 (.DIODE(_02303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19440__B1 (.DIODE(_02303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19437__B1 (.DIODE(_02303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19434__B1 (.DIODE(_02303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19429__B1 (.DIODE(_02303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19425__B1 (.DIODE(_02303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19503__B1 (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19499__B1 (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19495__B1 (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19491__B1 (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19487__B1 (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19483__B1 (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19479__B1 (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19475__B1 (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19429__C1 (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19425__C1 (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19491__A2 (.DIODE(_02310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19487__A2 (.DIODE(_02310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19483__A2 (.DIODE(_02310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19479__A2 (.DIODE(_02310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19475__A2 (.DIODE(_02310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19472__A2 (.DIODE(_02310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19469__A2 (.DIODE(_02310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19463__A2 (.DIODE(_02310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19450__A2 (.DIODE(_02310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19435__A2 (.DIODE(_02310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19462__C1 (.DIODE(_02311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19458__C1 (.DIODE(_02311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19455__C1 (.DIODE(_02311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19452__C1 (.DIODE(_02311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19449__C1 (.DIODE(_02311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19446__C1 (.DIODE(_02311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19443__C1 (.DIODE(_02311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19440__C1 (.DIODE(_02311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19437__C1 (.DIODE(_02311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19434__C1 (.DIODE(_02311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20050__C1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20048__C1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19919__C1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19777__C1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19775__C1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19473__C1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19470__C1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19467__C1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19464__C1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19461__C1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19616__C (.DIODE(_02363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19564__B (.DIODE(_02363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19511__C (.DIODE(_02363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19508__C (.DIODE(_02363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19507__A2 (.DIODE(_02363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19512__A (.DIODE(_02367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19542__S (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19539__S (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19536__S (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19533__S (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19530__S (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19527__S (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19524__S (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19521__S (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19518__S (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19514__S (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19583__A (.DIODE(_02393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19580__A (.DIODE(_02393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19577__A (.DIODE(_02393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19574__A (.DIODE(_02393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19571__A (.DIODE(_02393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19568__A (.DIODE(_02393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19562__A (.DIODE(_02393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19556__A (.DIODE(_02393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19553__A (.DIODE(_02393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19550__A (.DIODE(_02393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19613__S (.DIODE(_02405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19610__S (.DIODE(_02405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19607__S (.DIODE(_02405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19604__S (.DIODE(_02405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19601__S (.DIODE(_02405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19598__S (.DIODE(_02405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19566__A (.DIODE(_02405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19620__A (.DIODE(_02419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19614__A (.DIODE(_02419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19611__A (.DIODE(_02419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19608__A (.DIODE(_02419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19602__A (.DIODE(_02419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19599__A (.DIODE(_02419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19596__A (.DIODE(_02419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19593__A (.DIODE(_02419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19590__A (.DIODE(_02419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19587__A (.DIODE(_02419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19647__S (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19644__S (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19641__S (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19638__S (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19635__S (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19632__S (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19629__S (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19626__S (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19623__S (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19619__S (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19651__A (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19648__A (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19645__A (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19642__A (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19639__A (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19636__A (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19633__A (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19630__A (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19627__A (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19624__A (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19794__A (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19791__A (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19788__A (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19673__A (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19670__A (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19667__A (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19664__A (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19661__A (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19658__A (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19655__A (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19693__A (.DIODE(_02482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19692__A (.DIODE(_02482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19691__A (.DIODE(_02482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19690__A (.DIODE(_02482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19689__A (.DIODE(_02482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19688__A (.DIODE(_02482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19687__A (.DIODE(_02482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19686__A (.DIODE(_02482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19685__A (.DIODE(_02482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19684__A (.DIODE(_02482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19704__A (.DIODE(_02483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19703__A (.DIODE(_02483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19702__A (.DIODE(_02483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19701__A (.DIODE(_02483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19700__A (.DIODE(_02483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19699__A (.DIODE(_02483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19698__A (.DIODE(_02483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19697__A (.DIODE(_02483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19696__A (.DIODE(_02483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19695__A (.DIODE(_02483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19715__A (.DIODE(_02484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19714__A (.DIODE(_02484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19713__A (.DIODE(_02484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19712__A (.DIODE(_02484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19711__A (.DIODE(_02484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19710__A (.DIODE(_02484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19709__A (.DIODE(_02484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19708__A (.DIODE(_02484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19707__A (.DIODE(_02484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19706__A (.DIODE(_02484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19726__A (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19725__A (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19724__A (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19723__A (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19722__A (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19721__A (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19720__A (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19719__A (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19718__A (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19717__A (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20025__A (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20014__A (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20003__A (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19992__A (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19981__A (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19970__A (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19761__A (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19750__A (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19739__A (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19728__A (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19738__A (.DIODE(_02487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19737__A (.DIODE(_02487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19736__A (.DIODE(_02487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19735__A (.DIODE(_02487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19734__A (.DIODE(_02487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19733__A (.DIODE(_02487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19732__A (.DIODE(_02487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19731__A (.DIODE(_02487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19730__A (.DIODE(_02487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19729__A (.DIODE(_02487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19967__A (.DIODE(_02490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19966__A (.DIODE(_02490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19965__A (.DIODE(_02490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19964__A (.DIODE(_02490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19963__A (.DIODE(_02490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19766__A (.DIODE(_02490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19765__A (.DIODE(_02490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19764__A (.DIODE(_02490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19763__A (.DIODE(_02490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19762__A (.DIODE(_02490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19775__B1 (.DIODE(_02498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19777__B1 (.DIODE(_02499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19912__B (.DIODE(_02500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19859__B (.DIODE(_02500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19781__B (.DIODE(_02500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19780__A3 (.DIODE(_02500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19779__A2 (.DIODE(_02500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19856__S (.DIODE(_02503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19853__S (.DIODE(_02503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19835__S (.DIODE(_02503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19818__A (.DIODE(_02503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19786__A (.DIODE(_02503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19783__S (.DIODE(_02503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19785__A (.DIODE(_02505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19815__S (.DIODE(_02506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19812__S (.DIODE(_02506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19809__S (.DIODE(_02506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19806__S (.DIODE(_02506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19803__S (.DIODE(_02506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19800__S (.DIODE(_02506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19797__S (.DIODE(_02506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19793__S (.DIODE(_02506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19790__S (.DIODE(_02506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19787__S (.DIODE(_02506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19792__A (.DIODE(_02510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19814__A (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19816__B (.DIODE(_02526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19817__A (.DIODE(_02527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19850__S (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19847__S (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19844__S (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19841__S (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19838__S (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19832__S (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19829__S (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19825__S (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19822__S (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19819__S (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19820__B (.DIODE(_02529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19821__A (.DIODE(_02530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19823__B (.DIODE(_02531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19824__A (.DIODE(_02532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19826__B (.DIODE(_02533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19827__A (.DIODE(_02534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19863__A (.DIODE(_02535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19857__A (.DIODE(_02535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19854__A (.DIODE(_02535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19851__A (.DIODE(_02535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19848__A (.DIODE(_02535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19845__A (.DIODE(_02535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19842__A (.DIODE(_02535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19839__A (.DIODE(_02535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19833__A (.DIODE(_02535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19830__A (.DIODE(_02535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19830__B (.DIODE(_02536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19833__B (.DIODE(_02538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19909__S (.DIODE(_02557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19906__S (.DIODE(_02557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19903__S (.DIODE(_02557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19900__S (.DIODE(_02557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19897__S (.DIODE(_02557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19893__S (.DIODE(_02557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19861__A (.DIODE(_02557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19890__S (.DIODE(_02558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19887__S (.DIODE(_02558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19884__S (.DIODE(_02558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19881__S (.DIODE(_02558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19878__S (.DIODE(_02558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19875__S (.DIODE(_02558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19872__S (.DIODE(_02558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19869__S (.DIODE(_02558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19866__S (.DIODE(_02558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19862__S (.DIODE(_02558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19894__A (.DIODE(_02561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19891__A (.DIODE(_02561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19888__A (.DIODE(_02561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19885__A (.DIODE(_02561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19882__A (.DIODE(_02561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19879__A (.DIODE(_02561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19876__A (.DIODE(_02561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19873__A (.DIODE(_02561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19870__A (.DIODE(_02561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19867__A (.DIODE(_02561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19930__A (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19927__A (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19924__A (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19921__A (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19916__A (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19910__A (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19907__A (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19904__A (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19901__A (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19898__A (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19960__S (.DIODE(_02594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19957__S (.DIODE(_02594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19954__S (.DIODE(_02594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19951__S (.DIODE(_02594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19948__S (.DIODE(_02594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19945__S (.DIODE(_02594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19942__S (.DIODE(_02594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19914__A (.DIODE(_02594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19939__S (.DIODE(_02595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19936__S (.DIODE(_02595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19933__S (.DIODE(_02595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19929__S (.DIODE(_02595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19926__S (.DIODE(_02595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19923__S (.DIODE(_02595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19920__S (.DIODE(_02595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19919__A2 (.DIODE(_02595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19918__B (.DIODE(_02595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19915__S (.DIODE(_02595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19961__A (.DIODE(_02607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19958__A (.DIODE(_02607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19955__A (.DIODE(_02607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19952__A (.DIODE(_02607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19949__A (.DIODE(_02607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19946__A (.DIODE(_02607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19943__A (.DIODE(_02607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19940__A (.DIODE(_02607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19937__A (.DIODE(_02607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19934__A (.DIODE(_02607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19980__A (.DIODE(_02629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19979__A (.DIODE(_02629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19978__A (.DIODE(_02629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19977__A (.DIODE(_02629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19976__A (.DIODE(_02629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19975__A (.DIODE(_02629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19974__A (.DIODE(_02629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19973__A (.DIODE(_02629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19972__A (.DIODE(_02629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19971__A (.DIODE(_02629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19991__A (.DIODE(_02630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19990__A (.DIODE(_02630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19989__A (.DIODE(_02630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19988__A (.DIODE(_02630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19987__A (.DIODE(_02630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19986__A (.DIODE(_02630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19985__A (.DIODE(_02630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19984__A (.DIODE(_02630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19983__A (.DIODE(_02630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19982__A (.DIODE(_02630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20002__A (.DIODE(_02631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20001__A (.DIODE(_02631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20000__A (.DIODE(_02631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19999__A (.DIODE(_02631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19998__A (.DIODE(_02631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19997__A (.DIODE(_02631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19996__A (.DIODE(_02631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19995__A (.DIODE(_02631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19994__A (.DIODE(_02631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19993__A (.DIODE(_02631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20013__A (.DIODE(_02632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20012__A (.DIODE(_02632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20011__A (.DIODE(_02632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20010__A (.DIODE(_02632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20009__A (.DIODE(_02632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20008__A (.DIODE(_02632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20007__A (.DIODE(_02632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20006__A (.DIODE(_02632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20005__A (.DIODE(_02632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20004__A (.DIODE(_02632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20024__A (.DIODE(_02633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20023__A (.DIODE(_02633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20022__A (.DIODE(_02633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20021__A (.DIODE(_02633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20020__A (.DIODE(_02633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20019__A (.DIODE(_02633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20018__A (.DIODE(_02633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20017__A (.DIODE(_02633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20016__A (.DIODE(_02633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20015__A (.DIODE(_02633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20035__A (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20034__A (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20033__A (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20032__A (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20031__A (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20030__A (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20029__A (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20028__A (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20027__A (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20026__A (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20096__B1 (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20094__B1 (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20092__B1 (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20090__B1 (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20066__A (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20038__A (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20096__A2 (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20094__A2 (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20092__A2 (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20070__A (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20046__A (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20042__A2 (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20098__A2 (.DIODE(_02639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20095__A2 (.DIODE(_02639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20093__A2 (.DIODE(_02639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20069__A (.DIODE(_02639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20045__A (.DIODE(_02639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20042__C1 (.DIODE(_02639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20126__C1 (.DIODE(_02672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20124__C1 (.DIODE(_02672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20122__C1 (.DIODE(_02672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20117__C1 (.DIODE(_02672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20115__C1 (.DIODE(_02672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20113__C1 (.DIODE(_02672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20111__C1 (.DIODE(_02672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20109__C1 (.DIODE(_02672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20107__C1 (.DIODE(_02672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20098__C1 (.DIODE(_02672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20118__B (.DIODE(_02675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20103__B (.DIODE(_02675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10098__A1 (.DIODE(_02700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10091__A2 (.DIODE(_02700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10090__A (.DIODE(_02700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10071__A3 (.DIODE(_02700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10057__B (.DIODE(_02700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10177__B (.DIODE(_02704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10168__B (.DIODE(_02704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10164__B (.DIODE(_02704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10160__B (.DIODE(_02704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__B (.DIODE(_02704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10152__B (.DIODE(_02704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10146__B (.DIODE(_02704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10107__A (.DIODE(_02704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10061__A1 (.DIODE(_02704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10087__A1 (.DIODE(_02705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10061__B1 (.DIODE(_02705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19232__A1 (.DIODE(_02706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10105__C1 (.DIODE(_02706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10061__C1 (.DIODE(_02706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10250__A2 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10097__A (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10094__B1 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10092__A (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10066__B1 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10073__A (.DIODE(_02716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10269__S (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10267__S (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10265__S (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10263__S (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10261__S (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10087__S (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10085__S (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10082__S (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10080__S (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10078__S (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10247__A1 (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10138__S (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10134__S (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10130__S (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10126__S (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10122__S (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10118__S (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10112__S (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10103__A (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10085__A1 (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10243__A (.DIODE(_02729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10239__A (.DIODE(_02729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10235__A (.DIODE(_02729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10190__A (.DIODE(_02729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10172__A (.DIODE(_02729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10105__B1 (.DIODE(_02729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10093__B (.DIODE(_02729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10302__A2 (.DIODE(_02730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10301__B (.DIODE(_02730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10300__A2 (.DIODE(_02730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10299__A2 (.DIODE(_02730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10297__A2 (.DIODE(_02730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10294__A2 (.DIODE(_02730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10286__A2 (.DIODE(_02730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10094__A2 (.DIODE(_02730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10256__C (.DIODE(_02735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10254__D (.DIODE(_02735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10252__B1 (.DIODE(_02735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10249__B1 (.DIODE(_02735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10248__B1 (.DIODE(_02735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10245__B1 (.DIODE(_02735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10204__A (.DIODE(_02735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10150__A (.DIODE(_02735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10101__B (.DIODE(_02735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10100__A (.DIODE(_02735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10259__A2 (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10248__A1 (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10245__A1 (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10241__A1 (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10196__A (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10151__A (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10102__A (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10279__B (.DIODE(_02740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10170__B2 (.DIODE(_02740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10166__B2 (.DIODE(_02740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10162__B2 (.DIODE(_02740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10158__B2 (.DIODE(_02740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10154__B2 (.DIODE(_02740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10148__B2 (.DIODE(_02740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10144__B2 (.DIODE(_02740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10139__B2 (.DIODE(_02740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10109__A3 (.DIODE(_02740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10170__A1 (.DIODE(_02741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10166__A1 (.DIODE(_02741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10162__A1 (.DIODE(_02741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10158__A1 (.DIODE(_02741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10154__A1 (.DIODE(_02741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10106__A (.DIODE(_02741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19230__A1 (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10141__B (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10137__B (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10133__B (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10129__B (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10125__B (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10121__B (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10117__B (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10111__B (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10108__B (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10290__A1 (.DIODE(_02749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10283__A2 (.DIODE(_02749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10257__B1 (.DIODE(_02749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10251__B (.DIODE(_02749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10135__B2 (.DIODE(_02749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10131__B2 (.DIODE(_02749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10127__B2 (.DIODE(_02749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10123__B2 (.DIODE(_02749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10119__B2 (.DIODE(_02749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10115__B2 (.DIODE(_02749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10186__S (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10182__S (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10173__S (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10169__S (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10165__S (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10161__S (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10157__S (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10153__S (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10147__S (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10143__S (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10200__B1 (.DIODE(_02776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10195__B1 (.DIODE(_02776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10189__B1 (.DIODE(_02776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10185__B1 (.DIODE(_02776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10181__B1 (.DIODE(_02776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10171__A2 (.DIODE(_02776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10167__A2 (.DIODE(_02776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10163__A2 (.DIODE(_02776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10159__A2 (.DIODE(_02776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10155__A2 (.DIODE(_02776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10258__B2 (.DIODE(_02777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10195__A1 (.DIODE(_02777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10189__A1 (.DIODE(_02777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10185__A1 (.DIODE(_02777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10181__A1 (.DIODE(_02777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10171__B1 (.DIODE(_02777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10167__B1 (.DIODE(_02777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10163__B1 (.DIODE(_02777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10159__B1 (.DIODE(_02777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10155__B1 (.DIODE(_02777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10296__C1 (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10293__A (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10291__A2 (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10285__A (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10282__B1 (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10277__A2 (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10247__B1 (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10187__A (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10183__A (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10174__A (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13859__S (.DIODE(_02796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10246__A2 (.DIODE(_02796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10244__A2 (.DIODE(_02796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10240__A2 (.DIODE(_02796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10236__A2 (.DIODE(_02796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10232__A2 (.DIODE(_02796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10228__A2 (.DIODE(_02796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10224__A2 (.DIODE(_02796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10176__A (.DIODE(_02796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13396__S (.DIODE(_02798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10246__B1 (.DIODE(_02798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10244__B1 (.DIODE(_02798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10240__B1 (.DIODE(_02798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10236__B1 (.DIODE(_02798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10232__B1 (.DIODE(_02798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10228__B1 (.DIODE(_02798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10224__B1 (.DIODE(_02798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10178__A (.DIODE(_02798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10220__B1 (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10216__B1 (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10212__B1 (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10208__B1 (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10203__B1 (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10199__B1 (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10194__B1 (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10188__B1 (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10184__B1 (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10180__B1 (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10252__A2 (.DIODE(_02800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10249__A2 (.DIODE(_02800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10212__C1 (.DIODE(_02800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10208__C1 (.DIODE(_02800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10203__C1 (.DIODE(_02800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10199__C1 (.DIODE(_02800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10194__C1 (.DIODE(_02800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10188__C1 (.DIODE(_02800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10184__C1 (.DIODE(_02800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10180__C1 (.DIODE(_02800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10231__A (.DIODE(_02808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10227__A (.DIODE(_02808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10223__A (.DIODE(_02808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10219__A (.DIODE(_02808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10215__A (.DIODE(_02808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10211__A (.DIODE(_02808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10207__A (.DIODE(_02808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10202__A (.DIODE(_02808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10198__A (.DIODE(_02808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10193__A (.DIODE(_02808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10237__A1 (.DIODE(_02813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10233__A1 (.DIODE(_02813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10229__A1 (.DIODE(_02813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10225__A1 (.DIODE(_02813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10221__A1 (.DIODE(_02813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10217__A1 (.DIODE(_02813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10213__A1 (.DIODE(_02813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10209__A1 (.DIODE(_02813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10205__A1 (.DIODE(_02813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10200__A1 (.DIODE(_02813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10241__B1 (.DIODE(_02820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10237__B1 (.DIODE(_02820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10233__B1 (.DIODE(_02820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10229__B1 (.DIODE(_02820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10225__B1 (.DIODE(_02820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10221__B1 (.DIODE(_02820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10217__B1 (.DIODE(_02820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10213__B1 (.DIODE(_02820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10209__B1 (.DIODE(_02820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10205__B1 (.DIODE(_02820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13047__A1 (.DIODE(_02886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13035__B (.DIODE(_02886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13033__A1 (.DIODE(_02886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12996__A (.DIODE(_02886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12994__A (.DIODE(_02886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12968__A (.DIODE(_02886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12911__B1 (.DIODE(_02886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11744__A (.DIODE(_02886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11365__A (.DIODE(_02886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10304__A (.DIODE(_02886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12937__A (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12910__A1 (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12810__A (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12466__A (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12316__A (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11821__A (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11660__A (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11578__A (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11359__A (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10307__A (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10751__A2 (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__C (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10563__A2 (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10487__B (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10437__B (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10353__B (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10341__C (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10318__B (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10310__B (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10306__A (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10750__A2 (.DIODE(_02889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10488__B (.DIODE(_02889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10426__B (.DIODE(_02889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10421__A2 (.DIODE(_02889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10419__C (.DIODE(_02889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10346__B1 (.DIODE(_02889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10345__B (.DIODE(_02889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10327__A (.DIODE(_02889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10315__B1 (.DIODE(_02889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10307__B (.DIODE(_02889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13139__B1 (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13138__A (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__B1 (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11076__B1 (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10989__A (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10988__A (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10912__B1 (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10911__A (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10321__A (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10320__A (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12857__A (.DIODE(_02892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12448__A (.DIODE(_02892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12346__A (.DIODE(_02892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12298__A (.DIODE(_02892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11803__A (.DIODE(_02892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11726__A (.DIODE(_02892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11560__A (.DIODE(_02892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11286__A (.DIODE(_02892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11271__A (.DIODE(_02892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10310__A (.DIODE(_02892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11154__A (.DIODE(_02893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11135__A (.DIODE(_02893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11074__A (.DIODE(_02893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11057__A (.DIODE(_02893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10957__A (.DIODE(_02893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10894__A (.DIODE(_02893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10333__A (.DIODE(_02893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10319__A1_N (.DIODE(_02893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12858__B2 (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12603__A (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12503__A (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12449__B2 (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11978__B2 (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11977__A (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11561__B2 (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11424__A (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11345__A (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10312__A (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19800__A1 (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19465__A1 (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12615__B2 (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11132__B2 (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10955__B2 (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10906__A (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10892__A (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10332__A1 (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10319__B1 (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10315__A1 (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12603__B (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12503__B (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12449__A1 (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11978__A1 (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11977__B (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11727__A1 (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11561__A1 (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11424__B (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11345__B (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10314__A (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19797__A1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19463__A1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13011__B2 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12745__A1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12615__A1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11288__A1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11133__B (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11132__A1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10955__A1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10315__A2 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12965__A1 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12925__A1 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12896__B (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12895__A1 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12450__B (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__B (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11643__A1 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11562__B (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11485__B (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10317__A (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12993__A (.DIODE(_02900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12760__A1 (.DIODE(_02900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12732__A1 (.DIODE(_02900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12731__B (.DIODE(_02900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12616__B (.DIODE(_02900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12602__A1 (.DIODE(_02900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11423__A1 (.DIODE(_02900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11344__A1 (.DIODE(_02900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10954__A (.DIODE(_02900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10318__A (.DIODE(_02900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13047__B2 (.DIODE(_02906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13035__A (.DIODE(_02906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13033__B2 (.DIODE(_02906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13015__A (.DIODE(_02906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12997__A1 (.DIODE(_02906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12990__A (.DIODE(_02906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12934__A (.DIODE(_02906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12908__A (.DIODE(_02906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11364__A (.DIODE(_02906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10324__A (.DIODE(_02906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12318__A (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11826__A1 (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11823__A (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11749__A1 (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11746__A (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11662__A (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11580__A (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11376__A (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11371__A (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10325__A (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12905__A1 (.DIODE(_02908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12664__A1 (.DIODE(_02908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12652__A (.DIODE(_02908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12471__A1 (.DIODE(_02908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12321__A1 (.DIODE(_02908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12159__A (.DIODE(_02908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12052__A (.DIODE(_02908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12000__A1 (.DIODE(_02908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11583__A1 (.DIODE(_02908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10326__A (.DIODE(_02908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19793__A1 (.DIODE(_02909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19458__A1 (.DIODE(_02909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13154__A (.DIODE(_02909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13153__A1 (.DIODE(_02909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13140__A1 (.DIODE(_02909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13131__A (.DIODE(_02909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11157__A1 (.DIODE(_02909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11077__A1 (.DIODE(_02909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10913__A1 (.DIODE(_02909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10328__A (.DIODE(_02909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11077__A2 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10987__A2 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10913__A2 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10910__B (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10565__A2 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10480__A2 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10428__C (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10423__A2 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10408__A2 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10328__B (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11150__A (.DIODE(_02911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11070__A (.DIODE(_02911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10990__A1 (.DIODE(_02911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10982__A (.DIODE(_02911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10397__A2 (.DIODE(_02911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10329__B (.DIODE(_02911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13318__A (.DIODE(_02913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13302__A (.DIODE(_02913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13270__A (.DIODE(_02913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13213__A (.DIODE(_02913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13212__B1 (.DIODE(_02913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10840__A (.DIODE(_02913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10839__B1 (.DIODE(_02913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10584__A (.DIODE(_02913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10400__A (.DIODE(_02913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10331__A (.DIODE(_02913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13357__A1 (.DIODE(_02914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13316__A (.DIODE(_02914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13308__A (.DIODE(_02914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10685__A (.DIODE(_02914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10612__B1 (.DIODE(_02914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10611__A (.DIODE(_02914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10596__A1 (.DIODE(_02914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10592__A1 (.DIODE(_02914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10415__A (.DIODE(_02914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10402__A1 (.DIODE(_02914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13209__B (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10881__A (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10832__A1 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10827__A (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10755__A (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10681__A (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10643__A (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10642__A (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10392__A1 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10349__A (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12892__A1 (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12853__A1 (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12726__A1_N (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12725__C (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12721__A (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12136__A1 (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11414__A (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11339__A1 (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11044__A (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10335__A (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19803__A1 (.DIODE(_02918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19469__A1 (.DIODE(_02918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12957__A1 (.DIODE(_02918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12929__A (.DIODE(_02918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12754__A1 (.DIODE(_02918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10885__A1_N (.DIODE(_02918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10825__B2 (.DIODE(_02918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10750__A1 (.DIODE(_02918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10677__A1_N (.DIODE(_02918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10342__A (.DIODE(_02918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12293__A (.DIODE(_02919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12212__B2 (.DIODE(_02919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__B2 (.DIODE(_02919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11637__A (.DIODE(_02919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11554__B2 (.DIODE(_02919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11266__A (.DIODE(_02919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11262__B2 (.DIODE(_02919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10949__A (.DIODE(_02919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10625__A (.DIODE(_02919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10337__A (.DIODE(_02919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12590__A (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12292__B2 (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12213__A (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12133__B2 (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12019__B2 (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11797__B2 (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11721__A (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11260__A (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11046__A (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10338__A (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19809__A1 (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19475__A1 (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11970__A (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11128__A (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10887__B2 (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10751__B2 (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10674__B2 (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10638__B2 (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10346__A1 (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10341__A (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12595__B (.DIODE(_02922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12292__A1 (.DIODE(_02922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12213__B (.DIODE(_02922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12133__A1 (.DIODE(_02922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12019__A1 (.DIODE(_02922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11797__A1 (.DIODE(_02922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11721__B (.DIODE(_02922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11278__B (.DIODE(_02922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11046__B (.DIODE(_02922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10340__A (.DIODE(_02922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19806__A1 (.DIODE(_02923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19472__A1 (.DIODE(_02923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12892__B2 (.DIODE(_02923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11128__B (.DIODE(_02923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10887__A1 (.DIODE(_02923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10751__A1 (.DIODE(_02923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10674__A1 (.DIODE(_02923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10638__A1 (.DIODE(_02923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10346__A2 (.DIODE(_02923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10341__B (.DIODE(_02923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12854__B (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12445__A1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12295__A1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11967__A (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11800__A1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11336__A (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11279__A (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11268__A1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11126__A (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10344__A (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12755__A (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12737__A (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12610__A1 (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12596__A1 (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11973__A1 (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10943__A1_N (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10888__C (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10675__C (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10639__C (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10345__A (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12281__A1 (.DIODE(_02934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12117__A (.DIODE(_02934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11786__A1 (.DIODE(_02934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11781__A (.DIODE(_02934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11625__A1 (.DIODE(_02934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11246__A (.DIODE(_02934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11221__A1 (.DIODE(_02934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11215__A (.DIODE(_02934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10656__A (.DIODE(_02934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10352__A (.DIODE(_02934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12768__A (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12513__A1 (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12035__A (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11957__A1 (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11954__A (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11324__A1 (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11323__A (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11029__A (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10559__A (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10353__A (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12427__A1 (.DIODE(_02937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12425__B (.DIODE(_02937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12277__A1 (.DIODE(_02937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12116__B (.DIODE(_02937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11780__B (.DIODE(_02937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11621__A1 (.DIODE(_02937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11538__A1 (.DIODE(_02937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11247__A (.DIODE(_02937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11212__A1 (.DIODE(_02937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10355__A (.DIODE(_02937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12512__B (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12511__A1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12032__B (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11953__A1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11951__B (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11863__B (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11402__A1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11401__B (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11322__A1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10356__A (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11028__B (.DIODE(_02939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10936__B (.DIODE(_02939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10935__A1 (.DIODE(_02939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10872__B (.DIODE(_02939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10871__A1 (.DIODE(_02939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10763__B (.DIODE(_02939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10718__B (.DIODE(_02939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__A1 (.DIODE(_02939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10659__A1 (.DIODE(_02939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10363__A0 (.DIODE(_02939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12355__A1 (.DIODE(_02940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12196__A1 (.DIODE(_02940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12118__A1 (.DIODE(_02940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11782__A1 (.DIODE(_02940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11704__A1 (.DIODE(_02940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11537__B (.DIODE(_02940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11245__B (.DIODE(_02940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11218__A1 (.DIODE(_02940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11217__B (.DIODE(_02940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10358__A (.DIODE(_02940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11321__B (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11112__A1 (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11111__B (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11030__A1 (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10719__A (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10667__B (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10658__B (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__B (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10563__A1 (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__A (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12427__B2 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12355__B2 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12277__B2 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12196__B2 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11782__B2 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11704__B2 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11537__A (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11245__A (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11218__B2 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10361__A (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11951__A (.DIODE(_02944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11401__A (.DIODE(_02944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11321__A (.DIODE(_02944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11112__B2 (.DIODE(_02944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11111__A (.DIODE(_02944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11030__B2 (.DIODE(_02944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10667__A (.DIODE(_02944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10658__A (.DIODE(_02944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10386__A (.DIODE(_02944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10362__A (.DIODE(_02944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10388__B1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10364__B (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10573__A (.DIODE(_02947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10558__A (.DIODE(_02947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10482__A (.DIODE(_02947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10481__A (.DIODE(_02947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10477__A1 (.DIODE(_02947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10424__A (.DIODE(_02947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10411__A1 (.DIODE(_02947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10409__A (.DIODE(_02947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10391__A1 (.DIODE(_02947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10389__A (.DIODE(_02947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12515__B (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12106__A (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12038__A (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11938__A (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11850__A (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11387__A (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11310__A (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11228__A (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11185__A (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10366__A (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12563__A (.DIODE(_02949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12536__A1 (.DIODE(_02949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11100__A (.DIODE(_02949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11019__A (.DIODE(_02949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10928__A (.DIODE(_02949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10693__A1_N (.DIODE(_02949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10692__C (.DIODE(_02949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10652__A (.DIODE(_02949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10517__A (.DIODE(_02949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10367__A (.DIODE(_02949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19822__A1 (.DIODE(_02950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19491__A1 (.DIODE(_02950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13216__A1 (.DIODE(_02950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10809__A (.DIODE(_02950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10797__A1 (.DIODE(_02950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10480__A1 (.DIODE(_02950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10426__A (.DIODE(_02950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10423__A1 (.DIODE(_02950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10408__A1 (.DIODE(_02950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10385__A1 (.DIODE(_02950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11483__B (.DIODE(_02951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11016__A2 (.DIODE(_02951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10969__C (.DIODE(_02951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10751__B1 (.DIODE(_02951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10639__D (.DIODE(_02951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10631__A2 (.DIODE(_02951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__D (.DIODE(_02951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10563__B1 (.DIODE(_02951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10407__C (.DIODE(_02951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10369__A (.DIODE(_02951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13218__A2 (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13217__C (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10955__A2 (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10892__B (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10798__B (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10752__A1 (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10677__A2_N (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10518__B (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10406__A2 (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10370__A (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13131__B (.DIODE(_02953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11499__A2 (.DIODE(_02953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11441__B (.DIODE(_02953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11157__A2 (.DIODE(_02953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10906__B (.DIODE(_02953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10824__A (.DIODE(_02953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10434__B (.DIODE(_02953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10421__B1 (.DIODE(_02953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10420__A (.DIODE(_02953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10385__A2 (.DIODE(_02953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12360__A1 (.DIODE(_02954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12267__A1 (.DIODE(_02954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11772__B (.DIODE(_02954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11771__A1 (.DIODE(_02954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11693__A1 (.DIODE(_02954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11611__A1 (.DIODE(_02954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11201__B (.DIODE(_02954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11200__A1 (.DIODE(_02954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10382__A (.DIODE(_02954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10372__A (.DIODE(_02954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12536__B2 (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12515__A (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12040__B (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11942__B (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11940__A1 (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11313__B (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11312__A1 (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11104__A1 (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10726__B (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10373__A (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13225__A1 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13224__B (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11021__A1 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11020__B (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10929__B (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10772__A1 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10690__A1 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10654__B (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10649__A1 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10379__A1 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11093__C (.DIODE(_02957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11055__C (.DIODE(_02957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10954__B (.DIODE(_02957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10638__A2 (.DIODE(_02957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10636__C (.DIODE(_02957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10631__B1 (.DIODE(_02957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10628__D (.DIODE(_02957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10404__A (.DIODE(_02957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10384__C (.DIODE(_02957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10379__A2 (.DIODE(_02957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11385__C (.DIODE(_02958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11055__D (.DIODE(_02958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__C (.DIODE(_02958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10637__A (.DIODE(_02958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10636__D (.DIODE(_02958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10551__A2 (.DIODE(_02958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10550__C (.DIODE(_02958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10446__A (.DIODE(_02958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10384__D (.DIODE(_02958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10379__B1 (.DIODE(_02958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12267__B2 (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12266__A (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11772__A (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11771__B2 (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11611__B2 (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11610__A (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11201__A (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11200__B2 (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10380__A (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10377__A (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12040__A (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11942__A (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11940__B2 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11388__B2 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11313__A (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11312__B2 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11189__A (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11104__B2 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10726__A (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10378__A (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13225__B2 (.DIODE(_02961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13224__A (.DIODE(_02961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11021__B2 (.DIODE(_02961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11020__A (.DIODE(_02961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10929__A (.DIODE(_02961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10772__B2 (.DIODE(_02961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10690__B2 (.DIODE(_02961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10654__A (.DIODE(_02961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10649__B2 (.DIODE(_02961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10379__B2 (.DIODE(_02961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12418__A (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12185__A (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12107__B2 (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12039__B2 (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11852__A (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11692__A (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11527__A (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11389__A (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11230__B2 (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10381__A (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11103__A (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10860__B2 (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10859__A (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10771__A (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10727__B2 (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10689__A (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10551__B2 (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10550__A (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10405__A (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10384__A (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12418__B (.DIODE(_02965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12185__B (.DIODE(_02965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12039__A1 (.DIODE(_02965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11852__B (.DIODE(_02965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11527__B (.DIODE(_02965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11389__B (.DIODE(_02965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11388__A1 (.DIODE(_02965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11230__A1 (.DIODE(_02965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11189__B (.DIODE(_02965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10383__A (.DIODE(_02965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11103__B (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10860__A1 (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10859__B (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10771__B (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10727__A1 (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10689__B (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10551__A1 (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10550__B (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10403__A (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10384__B (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10391__A2 (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10389__B (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19819__A1 (.DIODE(_02969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19487__A1 (.DIODE(_02969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13218__B2 (.DIODE(_02969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13217__A (.DIODE(_02969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10800__B2 (.DIODE(_02969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10799__A (.DIODE(_02969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10764__B2 (.DIODE(_02969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10720__B2 (.DIODE(_02969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10718__A (.DIODE(_02969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10387__A (.DIODE(_02969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10598__A1 (.DIODE(_02971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10522__A (.DIODE(_02971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10484__A (.DIODE(_02971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10476__A (.DIODE(_02971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10465__A (.DIODE(_02971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10425__A (.DIODE(_02971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10410__A (.DIODE(_02971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10390__A (.DIODE(_02971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10794__A (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10398__A (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13320__A (.DIODE(_02981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13319__A (.DIODE(_02981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13303__A (.DIODE(_02981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13272__A (.DIODE(_02981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13271__A (.DIODE(_02981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13266__A (.DIODE(_02981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10842__A (.DIODE(_02981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10586__A (.DIODE(_02981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10585__A (.DIODE(_02981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10399__A (.DIODE(_02981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13383__A1 (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13337__A1 (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13309__A (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13215__A1 (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10687__A (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10614__A (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10504__A (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10417__A (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10416__A (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10401__A (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19825__A1 (.DIODE(_02986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19495__A1 (.DIODE(_02986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10927__A1 (.DIODE(_02986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10807__A1 (.DIODE(_02986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10806__B (.DIODE(_02986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10427__B (.DIODE(_02986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10421__A1 (.DIODE(_02986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10419__B (.DIODE(_02986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10407__B (.DIODE(_02986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10406__A1 (.DIODE(_02986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11422__B (.DIODE(_02987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10955__B1 (.DIODE(_02987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10885__A2_N (.DIODE(_02987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10800__A2 (.DIODE(_02987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10799__C (.DIODE(_02987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10675__D (.DIODE(_02987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10553__B (.DIODE(_02987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10439__A (.DIODE(_02987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10407__D (.DIODE(_02987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10406__B1 (.DIODE(_02987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19829__A1 (.DIODE(_02988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19499__A1 (.DIODE(_02988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10927__B2 (.DIODE(_02988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10807__B2 (.DIODE(_02988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10806__A (.DIODE(_02988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10427__A (.DIODE(_02988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10421__B2 (.DIODE(_02988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10419__A (.DIODE(_02988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10407__A (.DIODE(_02988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10406__B2 (.DIODE(_02988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12261__A (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12178__A (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12065__A (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11848__A (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11768__A (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11688__B2 (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11684__A (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11607__A (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11180__B2 (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10431__A (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12061__A (.DIODE(_03014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11930__A (.DIODE(_03014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11385__A (.DIODE(_03014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11308__A (.DIODE(_03014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11235__A (.DIODE(_03014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11094__B2 (.DIODE(_03014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11016__B2 (.DIODE(_03014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11015__A (.DIODE(_03014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10969__A (.DIODE(_03014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10432__A (.DIODE(_03014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11093__A (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10856__A (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10811__A (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10732__A (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10706__A (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10699__A (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10695__A (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10547__A (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10513__A (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10433__A (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19832__A1 (.DIODE(_03016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19503__A1 (.DIODE(_03016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10776__A (.DIODE(_03016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__A1 (.DIODE(_03016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10488__A (.DIODE(_03016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10485__A1 (.DIODE(_03016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10458__A (.DIODE(_03016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10447__A (.DIODE(_03016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10440__A (.DIODE(_03016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10434__A (.DIODE(_03016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12261__B (.DIODE(_03018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12178__B (.DIODE(_03018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12065__B (.DIODE(_03018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11848__B (.DIODE(_03018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11768__B (.DIODE(_03018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11688__A1 (.DIODE(_03018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11684__B (.DIODE(_03018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11520__B (.DIODE(_03018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11180__A1 (.DIODE(_03018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10436__A (.DIODE(_03018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12061__B (.DIODE(_03019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11930__B (.DIODE(_03019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11385__B (.DIODE(_03019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11308__B (.DIODE(_03019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11235__B (.DIODE(_03019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11094__A1 (.DIODE(_03019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11016__A1 (.DIODE(_03019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10969__B (.DIODE(_03019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10486__A (.DIODE(_03019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10437__A (.DIODE(_03019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10857__A (.DIODE(_03020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10733__A (.DIODE(_03020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10707__A (.DIODE(_03020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10700__A (.DIODE(_03020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10438__A (.DIODE(_03020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13229__A (.DIODE(_03021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10812__A (.DIODE(_03021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10777__A (.DIODE(_03021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10548__A (.DIODE(_03021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10514__A (.DIODE(_03021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__A3 (.DIODE(_03021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10485__A4 (.DIODE(_03021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10461__A (.DIODE(_03021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10448__A (.DIODE(_03021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10441__A (.DIODE(_03021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13218__B1 (.DIODE(_03022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13217__D (.DIODE(_03022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13154__B (.DIODE(_03022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13140__A2 (.DIODE(_03022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11438__A2 (.DIODE(_03022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11373__B (.DIODE(_03022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10762__B (.DIODE(_03022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10557__A2 (.DIODE(_03022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10485__A2 (.DIODE(_03022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10440__B (.DIODE(_03022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13227__B (.DIODE(_03029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13153__A2 (.DIODE(_03029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11502__B (.DIODE(_03029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11440__A2 (.DIODE(_03029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11369__A2 (.DIODE(_03029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11366__B (.DIODE(_03029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10800__B1 (.DIODE(_03029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10799__D (.DIODE(_03029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10717__B (.DIODE(_03029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10447__B (.DIODE(_03029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11485__C (.DIODE(_03038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11484__A2 (.DIODE(_03038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11308__C (.DIODE(_03038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10947__B (.DIODE(_03038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10887__A2 (.DIODE(_03038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10886__C (.DIODE(_03038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__D (.DIODE(_03038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10551__B1 (.DIODE(_03038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10550__D (.DIODE(_03038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10456__A (.DIODE(_03038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13225__A2 (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13224__C (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11133__D (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10764__B1 (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10763__D (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10720__A2 (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10718__C (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10674__B1 (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10657__B (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10457__A (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13216__A2 (.DIODE(_03040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11581__A2 (.DIODE(_03040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11578__B (.DIODE(_03040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11444__A2 (.DIODE(_03040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11443__B (.DIODE(_03040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11372__A2 (.DIODE(_03040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11287__B (.DIODE(_03040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11132__B1 (.DIODE(_03040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10809__B (.DIODE(_03040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10458__B (.DIODE(_03040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13051__A1 (.DIODE(_03069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13030__A (.DIODE(_03069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12577__A1_N (.DIODE(_03069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12563__B (.DIODE(_03069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12538__A1 (.DIODE(_03069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12537__C (.DIODE(_03069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12421__A (.DIODE(_03069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11093__B (.DIODE(_03069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10851__A (.DIODE(_03069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10487__A (.DIODE(_03069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10601__B (.DIODE(_03072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__B1 (.DIODE(_03072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11485__D (.DIODE(_03093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11484__B1 (.DIODE(_03093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11424__C (.DIODE(_03093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11235__C (.DIODE(_03093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11044__B (.DIODE(_03093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10950__A2 (.DIODE(_03093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10945__C (.DIODE(_03093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10886__D (.DIODE(_03093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10658__C (.DIODE(_03093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10511__A (.DIODE(_03093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13225__B1 (.DIODE(_03094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13224__D (.DIODE(_03094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11423__A2 (.DIODE(_03094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11271__B (.DIODE(_03094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10887__B1 (.DIODE(_03094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10807__A2 (.DIODE(_03094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10806__C (.DIODE(_03094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10718__D (.DIODE(_03094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10659__A2 (.DIODE(_03094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10512__A (.DIODE(_03094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11663__A2 (.DIODE(_03095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11660__B (.DIODE(_03095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11377__A2 (.DIODE(_03095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11375__B (.DIODE(_03095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11363__A2 (.DIODE(_03095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10797__A2 (.DIODE(_03095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10774__B (.DIODE(_03095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10720__B1 (.DIODE(_03095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10663__B (.DIODE(_03095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10513__B (.DIODE(_03095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10549__A (.DIODE(_03096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10520__A2_N (.DIODE(_03096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10514__B (.DIODE(_03096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13227__A (.DIODE(_03100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12565__B2 (.DIODE(_03100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10866__A1 (.DIODE(_03100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10862__A (.DIODE(_03100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10774__A (.DIODE(_03100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10761__A1 (.DIODE(_03100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10729__A (.DIODE(_03100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10557__A1 (.DIODE(_03100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10553__A (.DIODE(_03100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10518__A (.DIODE(_03100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11424__D (.DIODE(_03127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11345__C (.DIODE(_03127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11182__C (.DIODE(_03127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11126__B (.DIODE(_03127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11046__C (.DIODE(_03127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11045__A2 (.DIODE(_03127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10950__B1 (.DIODE(_03127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10945__D (.DIODE(_03127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10771__C (.DIODE(_03127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10545__A (.DIODE(_03127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11560__B (.DIODE(_03128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11423__B1 (.DIODE(_03128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11344__A2 (.DIODE(_03128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10806__D (.DIODE(_03128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10772__A2 (.DIODE(_03128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10667__C (.DIODE(_03128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__A2 (.DIODE(_03128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10659__B1 (.DIODE(_03128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10658__D (.DIODE(_03128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10546__A (.DIODE(_03128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11747__A2 (.DIODE(_03129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11744__B (.DIODE(_03129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11583__A2 (.DIODE(_03129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11577__A2 (.DIODE(_03129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11368__B (.DIODE(_03129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10870__B (.DIODE(_03129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10807__B1 (.DIODE(_03129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10761__A2 (.DIODE(_03129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10729__B (.DIODE(_03129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10547__B (.DIODE(_03129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13255__A (.DIODE(_03137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10555__B2 (.DIODE(_03137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10573__B (.DIODE(_03140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10558__B (.DIODE(_03140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19812__A1 (.DIODE(_03142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19479__A1 (.DIODE(_03142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12850__B2 (.DIODE(_03142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12715__A (.DIODE(_03142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12585__A1 (.DIODE(_03142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10870__A (.DIODE(_03142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10798__A (.DIODE(_03142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10762__A (.DIODE(_03142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10717__A (.DIODE(_03142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10565__A1 (.DIODE(_03142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12425__A (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12275__A (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12116__A (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11780__A (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11621__B2 (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11538__B2 (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11216__A (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11212__B2 (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11209__A (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10561__A (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12569__B2 (.DIODE(_03144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12512__A (.DIODE(_03144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12511__B2 (.DIODE(_03144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12354__A (.DIODE(_03144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12032__A (.DIODE(_03144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11953__B2 (.DIODE(_03144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11863__A (.DIODE(_03144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11402__B2 (.DIODE(_03144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11322__B2 (.DIODE(_03144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10562__A (.DIODE(_03144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11028__A (.DIODE(_03145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10936__A (.DIODE(_03145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10935__B2 (.DIODE(_03145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10872__A (.DIODE(_03145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10871__B2 (.DIODE(_03145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10763__A (.DIODE(_03145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__B2 (.DIODE(_03145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10659__B2 (.DIODE(_03145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__A (.DIODE(_03145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10563__B2 (.DIODE(_03145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12739__B2 (.DIODE(_03208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12719__A (.DIODE(_03208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12592__B2 (.DIODE(_03208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12493__B2 (.DIODE(_03208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12020__A (.DIODE(_03208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11415__A (.DIODE(_03208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11280__B2 (.DIODE(_03208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11127__B2 (.DIODE(_03208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10631__B2 (.DIODE(_03208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10628__A (.DIODE(_03208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12293__B (.DIODE(_03209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12212__A1 (.DIODE(_03209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11798__B (.DIODE(_03209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__A1 (.DIODE(_03209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11636__A1 (.DIODE(_03209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11554__A1 (.DIODE(_03209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11266__B (.DIODE(_03209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11262__A1 (.DIODE(_03209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10948__A (.DIODE(_03209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10627__A (.DIODE(_03209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12592__A1 (.DIODE(_03210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12493__A1 (.DIODE(_03210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12020__B (.DIODE(_03210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11883__B (.DIODE(_03210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11415__B (.DIODE(_03210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11335__B (.DIODE(_03210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11280__A1 (.DIODE(_03210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11127__A1 (.DIODE(_03210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10886__B (.DIODE(_03210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10628__B (.DIODE(_03210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10750__B1 (.DIODE(_03211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10632__A_N (.DIODE(_03211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12720__A1 (.DIODE(_03212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12590__B (.DIODE(_03212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12443__B (.DIODE(_03212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12340__A1 (.DIODE(_03212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12134__B (.DIODE(_03212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11555__B (.DIODE(_03212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11265__A1 (.DIODE(_03212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11260__B (.DIODE(_03212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10945__B (.DIODE(_03212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10630__A (.DIODE(_03212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12854__A (.DIODE(_03213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12724__A1 (.DIODE(_03213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12495__B (.DIODE(_03213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11970__B (.DIODE(_03213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11969__A1 (.DIODE(_03213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11416__A1 (.DIODE(_03213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11045__A1 (.DIODE(_03213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__B (.DIODE(_03213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10636__B (.DIODE(_03213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10631__A1 (.DIODE(_03213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10750__A3 (.DIODE(_03214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10632__B (.DIODE(_03214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12720__B2 (.DIODE(_03217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12443__A (.DIODE(_03217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12340__B2 (.DIODE(_03217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12134__A (.DIODE(_03217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11798__A (.DIODE(_03217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11636__B2 (.DIODE(_03217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11555__A (.DIODE(_03217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11265__B2 (.DIODE(_03217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10945__A (.DIODE(_03217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10635__A (.DIODE(_03217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12724__B2 (.DIODE(_03218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12495__A (.DIODE(_03218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11969__B2 (.DIODE(_03218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11883__A (.DIODE(_03218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11416__B2 (.DIODE(_03218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11335__A (.DIODE(_03218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11045__B2 (.DIODE(_03218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10886__A (.DIODE(_03218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__A (.DIODE(_03218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10636__A (.DIODE(_03218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11343__B (.DIODE(_03220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11133__C (.DIODE(_03220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11132__A2 (.DIODE(_03220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11052__B (.DIODE(_03220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10943__A2_N (.DIODE(_03220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10888__D (.DIODE(_03220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10764__A2 (.DIODE(_03220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10763__C (.DIODE(_03220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10674__A2 (.DIODE(_03220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10638__B1 (.DIODE(_03220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11562__C (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11561__A2 (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11415__D (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11337__A2 (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11335__C (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11279__B (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11273__D (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11272__B1 (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10689__D (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10646__A (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11803__B (.DIODE(_03229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11468__A2 (.DIODE(_03229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11416__B1 (.DIODE(_03229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11030__A2 (.DIODE(_03229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11028__C (.DIODE(_03229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10936__D (.DIODE(_03229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10731__A (.DIODE(_03229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10690__B1 (.DIODE(_03229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10654__C (.DIODE(_03229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10649__A2 (.DIODE(_03229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11688__A2 (.DIODE(_03230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11644__C (.DIODE(_03230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11643__A2 (.DIODE(_03230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11562__D (.DIODE(_03230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11337__B1 (.DIODE(_03230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11280__A2 (.DIODE(_03230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11278__C (.DIODE(_03230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11261__B (.DIODE(_03230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10653__A (.DIODE(_03230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10648__A (.DIODE(_03230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12053__A2 (.DIODE(_03231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12050__B (.DIODE(_03231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11911__A2 (.DIODE(_03231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11905__A2 (.DIODE(_03231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11888__B (.DIODE(_03231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11823__B (.DIODE(_03231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11028__D (.DIODE(_03231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10928__B (.DIODE(_03231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10695__B (.DIODE(_03231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10649__B1 (.DIODE(_03231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11520__C (.DIODE(_03233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11416__A2 (.DIODE(_03233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11415__C (.DIODE(_03233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11336__B (.DIODE(_03233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11273__C (.DIODE(_03233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11272__A2 (.DIODE(_03233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11127__B1 (.DIODE(_03233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10726__D (.DIODE(_03233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10688__A (.DIODE(_03233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10651__A (.DIODE(_03233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11909__A2 (.DIODE(_03234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11906__B (.DIODE(_03234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11749__A2 (.DIODE(_03234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11743__A2 (.DIODE(_03234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11662__B (.DIODE(_03234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11288__B1 (.DIODE(_03234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10935__A2 (.DIODE(_03234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10871__B1 (.DIODE(_03234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10776__B (.DIODE(_03234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10652__B (.DIODE(_03234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11561__B1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11400__B (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11335__D (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11268__A2 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11112__A2 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11111__C (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11030__B1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10860__A2 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10859__C (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10654__D (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12711__A1 (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12710__B (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12581__A (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12574__A1 (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12567__A (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11468__A1 (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11113__A (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10934__A (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10663__A (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10657__A (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10724__B1_N (.DIODE(_03241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10660__A (.DIODE(_03241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11345__D (.DIODE(_03247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11291__C (.DIODE(_03247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11178__C (.DIODE(_03247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11127__A2 (.DIODE(_03247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11046__D (.DIODE(_03247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10771__D (.DIODE(_03247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10727__A2 (.DIODE(_03247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10726__C (.DIODE(_03247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10691__A (.DIODE(_03247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10665__A (.DIODE(_03247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11642__B (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11414__B (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11344__B1 (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11288__A2 (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11128__C (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11045__B1 (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10872__C (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10772__B1 (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10667__D (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__B1 (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11726__B (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11339__A2 (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11291__D (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11128__D (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11029__B (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10936__C (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10872__D (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10727__B1 (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10690__A2 (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10689__C (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10716__A (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10693__B1 (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10692__A_N (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11824__A2 (.DIODE(_03274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11821__B (.DIODE(_03274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11665__A2 (.DIODE(_03274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11659__A2 (.DIODE(_03274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11580__B (.DIODE(_03274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10934__B (.DIODE(_03274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10871__A2 (.DIODE(_03274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10811__B (.DIODE(_03274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10693__A2_N (.DIODE(_03274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10692__D (.DIODE(_03274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11764__C (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__C (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11644__D (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11643__B1 (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11402__A2 (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11278__D (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11264__B (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11262__A2 (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11260__C (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10697__A (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11727__A2 (.DIODE(_03280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11401__C (.DIODE(_03280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11324__A2 (.DIODE(_03280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11280__B1 (.DIODE(_03280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11112__B1 (.DIODE(_03280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11111__D (.DIODE(_03280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10929__C (.DIODE(_03280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10860__B1 (.DIODE(_03280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10859__D (.DIODE(_03280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10698__A (.DIODE(_03280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12160__A2 (.DIODE(_03281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12157__B (.DIODE(_03281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12000__A2 (.DIODE(_03281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11993__A2 (.DIODE(_03281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11976__B (.DIODE(_03281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11908__B (.DIODE(_03281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11323__B (.DIODE(_03281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11019__B (.DIODE(_03281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10927__A2 (.DIODE(_03281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10699__B (.DIODE(_03281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10736__A2_N (.DIODE(_03282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10708__A (.DIODE(_03282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10700__B (.DIODE(_03282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11847__A2 (.DIODE(_03286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11805__C (.DIODE(_03286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__D (.DIODE(_03286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11553__B (.DIODE(_03286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11322__A2 (.DIODE(_03286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11265__A2 (.DIODE(_03286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11262__B1 (.DIODE(_03286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11260__D (.DIODE(_03286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11246__B (.DIODE(_03286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10704__A (.DIODE(_03286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11804__A2 (.DIODE(_03287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11727__B1 (.DIODE(_03287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11639__A2 (.DIODE(_03287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11402__B1 (.DIODE(_03287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11401__D (.DIODE(_03287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11321__C (.DIODE(_03287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11100__B (.DIODE(_03287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11021__A2 (.DIODE(_03287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10929__D (.DIODE(_03287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10705__A (.DIODE(_03287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12239__A2 (.DIODE(_03288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12236__B (.DIODE(_03288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12049__A2 (.DIODE(_03288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12048__A2 (.DIODE(_03288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12025__B (.DIODE(_03288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11997__B (.DIODE(_03288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11020__C (.DIODE(_03288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10927__B1 (.DIODE(_03288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10855__A (.DIODE(_03288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10706__B (.DIODE(_03288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10748__A (.DIODE(_03299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10723__A (.DIODE(_03299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19815__A1 (.DIODE(_03302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19483__A1 (.DIODE(_03302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13218__A1 (.DIODE(_03302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13217__B (.DIODE(_03302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12711__B2 (.DIODE(_03302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12710__A (.DIODE(_03302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10800__A1 (.DIODE(_03302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10799__B (.DIODE(_03302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10764__A1 (.DIODE(_03302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10720__A1 (.DIODE(_03302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10761__B1 (.DIODE(_03309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10728__A_N (.DIODE(_03309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10761__A3 (.DIODE(_03310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10728__B (.DIODE(_03310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11995__A2 (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11994__B (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11826__A2 (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11820__A2 (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11746__B (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11113__B (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10935__B1 (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10866__A2 (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10862__B (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10732__B (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10815__A2 (.DIODE(_03315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10777__B (.DIODE(_03315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10734__A (.DIODE(_03315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10797__B1 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10773__A (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13256__A2_N (.DIODE(_03394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13229__B (.DIODE(_03394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10813__A (.DIODE(_03394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13010__A (.DIODE(_03434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13009__A1 (.DIODE(_03434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12986__A (.DIODE(_03434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12983__A1 (.DIODE(_03434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12767__A (.DIODE(_03434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12715__B (.DIODE(_03434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12713__A1_N (.DIODE(_03434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12712__C (.DIODE(_03434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12565__A1 (.DIODE(_03434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10852__A (.DIODE(_03434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19790__A1 (.DIODE(_03435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19455__A1 (.DIODE(_03435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13059__B2 (.DIODE(_03435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13008__A (.DIODE(_03435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12958__A (.DIODE(_03435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12943__A (.DIODE(_03435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12942__A1 (.DIODE(_03435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12902__A (.DIODE(_03435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12850__A1 (.DIODE(_03435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10864__A1 (.DIODE(_03435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11933__A2 (.DIODE(_03436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11805__D (.DIODE(_03436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11635__B (.DIODE(_03436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11555__C (.DIODE(_03436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11554__A2 (.DIODE(_03436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11387__B (.DIODE(_03436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11265__B1 (.DIODE(_03436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11248__A2 (.DIODE(_03436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11245__C (.DIODE(_03436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10854__A (.DIODE(_03436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12319__A2 (.DIODE(_03437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12316__B (.DIODE(_03437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12162__A2 (.DIODE(_03437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12156__A2 (.DIODE(_03437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12139__B (.DIODE(_03437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12052__B (.DIODE(_03437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11021__B1 (.DIODE(_03437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11020__D (.DIODE(_03437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10864__A2 (.DIODE(_03437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10856__B (.DIODE(_03437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10879__A (.DIODE(_03449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10869__A (.DIODE(_03449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13050__A (.DIODE(_03490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12600__A (.DIODE(_03490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12500__A (.DIODE(_03490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12218__A (.DIODE(_03490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12139__A (.DIODE(_03490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11976__A (.DIODE(_03490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11888__A (.DIODE(_03490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11483__A (.DIODE(_03490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11343__A (.DIODE(_03490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10908__A (.DIODE(_03490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12868__A1 (.DIODE(_03491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12809__A1 (.DIODE(_03491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12743__A (.DIODE(_03491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12730__A (.DIODE(_03491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12613__A (.DIODE(_03491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12465__A1 (.DIODE(_03491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12315__A1 (.DIODE(_03491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11905__A1 (.DIODE(_03491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11820__A1 (.DIODE(_03491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10909__A (.DIODE(_03491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19787__A1 (.DIODE(_03492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19452__A1 (.DIODE(_03492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13065__A (.DIODE(_03492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13059__A1 (.DIODE(_03492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13031__A1 (.DIODE(_03492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12649__A1 (.DIODE(_03492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12156__A1 (.DIODE(_03492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12049__A1 (.DIODE(_03492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10987__A1 (.DIODE(_03492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10910__A (.DIODE(_03492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12591__A (.DIODE(_03529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12492__A (.DIODE(_03529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12441__A (.DIODE(_03529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12291__A (.DIODE(_03529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12132__A (.DIODE(_03529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12018__A (.DIODE(_03529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11881__A (.DIODE(_03529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11796__A (.DIODE(_03529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11639__A1 (.DIODE(_03529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10947__A (.DIODE(_03529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12739__A1 (.DIODE(_03531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12738__B (.DIODE(_03531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12723__B (.DIODE(_03531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12719__B (.DIODE(_03531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12594__A1 (.DIODE(_03531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12442__A1 (.DIODE(_03531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12341__B (.DIODE(_03531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11882__A1 (.DIODE(_03531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11337__A1 (.DIODE(_03531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10950__A1 (.DIODE(_03531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12738__A (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12723__A (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12595__A (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12594__B2 (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12442__B2 (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12341__A (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11882__B2 (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11337__B2 (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11278__A (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10950__B2 (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10959__A2 (.DIODE(_03535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10953__B (.DIODE(_03535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12061__C (.DIODE(_03551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11978__A2 (.DIODE(_03551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11890__D (.DIODE(_03551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11800__A2 (.DIODE(_03551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11310__B (.DIODE(_03551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11248__B1 (.DIODE(_03551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11104__B1 (.DIODE(_03551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11102__A (.DIODE(_03551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11016__B1 (.DIODE(_03551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10969__D (.DIODE(_03551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11018__A1 (.DIODE(_03552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11017__B (.DIODE(_03552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10972__A (.DIODE(_03552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10971__A (.DIODE(_03552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12385__A1 (.DIODE(_03596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12104__B (.DIODE(_03596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12099__B (.DIODE(_03596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11933__A1 (.DIODE(_03596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11383__A1 (.DIODE(_03596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11306__A1 (.DIODE(_03596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11305__B (.DIODE(_03596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11233__A1 (.DIODE(_03596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11182__B (.DIODE(_03596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11015__B (.DIODE(_03596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11977__C (.DIODE(_03597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11796__B (.DIODE(_03597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11721__C (.DIODE(_03597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11625__A2 (.DIODE(_03597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11388__B1 (.DIODE(_03597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11313__C (.DIODE(_03597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11312__A2 (.DIODE(_03597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11228__B (.DIODE(_03597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11094__B1 (.DIODE(_03597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11015__D (.DIODE(_03597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11090__B1 (.DIODE(_03605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11033__B (.DIODE(_03605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11024__C_N (.DIODE(_03605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11090__B2 (.DIODE(_03606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11024__D_N (.DIODE(_03606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11027__B (.DIODE(_03608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11026__B_N (.DIODE(_03608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11118__A1 (.DIODE(_03614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11117__B (.DIODE(_03614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11032__B (.DIODE(_03614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12965__B2 (.DIODE(_03633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12925__B2 (.DIODE(_03633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12895__B2 (.DIODE(_03633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12859__A (.DIODE(_03633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12450__A (.DIODE(_03633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__A (.DIODE(_03633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11643__B2 (.DIODE(_03633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11562__A (.DIODE(_03633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11485__A (.DIODE(_03633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11051__A (.DIODE(_03633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12760__B2 (.DIODE(_03634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12745__B2 (.DIODE(_03634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12732__B2 (.DIODE(_03634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12731__A (.DIODE(_03634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12616__A (.DIODE(_03634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12602__B2 (.DIODE(_03634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11423__B2 (.DIODE(_03634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11288__B2 (.DIODE(_03634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11133__A (.DIODE(_03634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11052__A (.DIODE(_03634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12966__A (.DIODE(_03636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12348__A (.DIODE(_03636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12299__B2 (.DIODE(_03636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12220__A (.DIODE(_03636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12141__A (.DIODE(_03636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11890__A (.DIODE(_03636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11804__B2 (.DIODE(_03636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11727__B2 (.DIODE(_03636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11272__B2 (.DIODE(_03636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11055__A (.DIODE(_03636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12966__B (.DIODE(_03637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12859__B (.DIODE(_03637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12348__B (.DIODE(_03637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12299__A1 (.DIODE(_03637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12220__B (.DIODE(_03637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12141__B (.DIODE(_03637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11890__B (.DIODE(_03637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11804__A1 (.DIODE(_03637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11272__A1 (.DIODE(_03637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11055__B (.DIODE(_03637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12102__A2 (.DIODE(_03674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12099__C (.DIODE(_03674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__A2 (.DIODE(_03674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11637__D (.DIODE(_03674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11636__B1 (.DIODE(_03674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11389__D (.DIODE(_03674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11218__B1 (.DIODE(_03674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11217__D (.DIODE(_03674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11212__A2 (.DIODE(_03674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11092__A (.DIODE(_03674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12469__A2 (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12466__B (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12321__A2 (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12315__A2 (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12298__B (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12238__B (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12026__A2 (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11978__B1 (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11539__B (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11093__D (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12102__B2 (.DIODE(_03678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12064__B2 (.DIODE(_03678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11935__A (.DIODE(_03678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11847__B2 (.DIODE(_03678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11844__A (.DIODE(_03678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11603__A (.DIODE(_03678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11520__A (.DIODE(_03678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11233__B2 (.DIODE(_03678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11232__A (.DIODE(_03678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11098__A (.DIODE(_03678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12102__A1 (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12064__A1 (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11935__B (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11847__A1 (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11844__B (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11764__B (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11603__B (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11232__B (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11178__B (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11098__B (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12104__C (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11798__C (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__B1 (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11620__B (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11538__A2 (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11537__C (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11230__A2 (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11212__B1 (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11185__B (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11098__D (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11384__B (.DIODE(_03681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11107__A (.DIODE(_03681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11099__B1 (.DIODE(_03681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11930__C (.DIODE(_03684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11890__C (.DIODE(_03684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11889__A2 (.DIODE(_03684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11804__B1 (.DIODE(_03684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11322__B1 (.DIODE(_03684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11321__D (.DIODE(_03684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11221__A2 (.DIODE(_03684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11219__B (.DIODE(_03684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11104__A2 (.DIODE(_03684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11103__C (.DIODE(_03684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12375__A2 (.DIODE(_03685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12372__B (.DIODE(_03685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12241__A2 (.DIODE(_03685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12235__A2 (.DIODE(_03685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12218__B (.DIODE(_03685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12159__B (.DIODE(_03685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11993__B2 (.DIODE(_03685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11979__A1 (.DIODE(_03685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11889__B1 (.DIODE(_03685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11103__D (.DIODE(_03685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11118__A2 (.DIODE(_03699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11117__C (.DIODE(_03699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11144__B (.DIODE(_03705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11123__B (.DIODE(_03705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11131__B1 (.DIODE(_03712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11130__C (.DIODE(_03712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11141__B1 (.DIODE(_03721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11140__A (.DIODE(_03721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13417__A (.DIODE(_03755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13409__A1 (.DIODE(_03755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13353__A1 (.DIODE(_03755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12181__B2 (.DIODE(_03756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11767__B2 (.DIODE(_03756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11689__A (.DIODE(_03756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11606__B2 (.DIODE(_03756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11523__B2 (.DIODE(_03756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11197__A (.DIODE(_03756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11196__B2 (.DIODE(_03756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11183__A (.DIODE(_03756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11176__A (.DIODE(_03756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11175__A (.DIODE(_03756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12181__A1 (.DIODE(_03757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11767__A1 (.DIODE(_03757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11689__B (.DIODE(_03757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11607__B (.DIODE(_03757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11606__A1 (.DIODE(_03757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11523__A1 (.DIODE(_03757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11197__B (.DIODE(_03757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11196__A1 (.DIODE(_03757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11183__B (.DIODE(_03757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11175__B (.DIODE(_03757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12385__B2 (.DIODE(_03759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12104__A (.DIODE(_03759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12099__A (.DIODE(_03759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11933__B2 (.DIODE(_03759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11764__A (.DIODE(_03759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11383__B2 (.DIODE(_03759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11306__B2 (.DIODE(_03759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11305__A (.DIODE(_03759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11182__A (.DIODE(_03759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11178__A (.DIODE(_03759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12134__C (.DIODE(_03760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12133__A2 (.DIODE(_03760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11866__A2 (.DIODE(_03760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11861__A (.DIODE(_03760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11782__B1 (.DIODE(_03760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11691__B (.DIODE(_03760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11528__B1 (.DIODE(_03760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11527__D (.DIODE(_03760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11196__B1 (.DIODE(_03760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11178__D (.DIODE(_03760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11864__A (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11782__A2 (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11704__B1 (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11702__D (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11609__B (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11528__A2 (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11527__C (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11200__B1 (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11182__D (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11180__B1 (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12261__C (.DIODE(_03769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11798__D (.DIODE(_03769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11621__A2 (.DIODE(_03769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11538__B1 (.DIODE(_03769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11537__D (.DIODE(_03769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11305__D (.DIODE(_03769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11227__D (.DIODE(_03769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11199__B (.DIODE(_03769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11192__A2 (.DIODE(_03769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11189__C (.DIODE(_03769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11968__A (.DIODE(_03770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11781__B (.DIODE(_03770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11704__A2 (.DIODE(_03770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11621__B1 (.DIODE(_03770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11526__B (.DIODE(_03770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11233__B1 (.DIODE(_03770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11232__D (.DIODE(_03770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11200__A2 (.DIODE(_03770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11192__B1 (.DIODE(_03770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11188__A (.DIODE(_03770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12385__A2 (.DIODE(_03771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12300__C (.DIODE(_03771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12299__A2 (.DIODE(_03771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12220__D (.DIODE(_03771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12018__B (.DIODE(_03771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11883__D (.DIODE(_03771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11882__B1 (.DIODE(_03771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11702__C (.DIODE(_03771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11235__D (.DIODE(_03771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11189__D (.DIODE(_03771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12417__A1 (.DIODE(_03773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12362__B (.DIODE(_03773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12186__A1 (.DIODE(_03773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12108__B (.DIODE(_03773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12107__A1 (.DIODE(_03773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11851__A1 (.DIODE(_03773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11692__B (.DIODE(_03773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11528__A1 (.DIODE(_03773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11227__B (.DIODE(_03773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11192__A1 (.DIODE(_03773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12417__B2 (.DIODE(_03774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12362__A (.DIODE(_03774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12360__B2 (.DIODE(_03774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12186__B2 (.DIODE(_03774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12108__A (.DIODE(_03774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11851__B2 (.DIODE(_03774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11693__B2 (.DIODE(_03774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11528__B2 (.DIODE(_03774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11227__A (.DIODE(_03774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11192__B2 (.DIODE(_03774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12064__A2 (.DIODE(_03793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11719__B (.DIODE(_03793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11636__A2 (.DIODE(_03793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11555__D (.DIODE(_03793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11554__B1 (.DIODE(_03793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11389__C (.DIODE(_03793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11388__A2 (.DIODE(_03793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11218__A2 (.DIODE(_03793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11217__C (.DIODE(_03793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11211__B (.DIODE(_03793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12431__A1 (.DIODE(_03798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12356__A (.DIODE(_03798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12197__A (.DIODE(_03798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12122__A1 (.DIODE(_03798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12037__A1 (.DIODE(_03798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11867__A (.DIODE(_03798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11705__A (.DIODE(_03798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11539__A (.DIODE(_03798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11400__A (.DIODE(_03798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11219__A (.DIODE(_03798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12573__A (.DIODE(_03799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12572__B2 (.DIODE(_03799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12568__A (.DIODE(_03799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12195__A (.DIODE(_03799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12118__B2 (.DIODE(_03799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12034__B2 (.DIODE(_03799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11866__B2 (.DIODE(_03799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11702__A (.DIODE(_03799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11248__B2 (.DIODE(_03799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11217__A (.DIODE(_03799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12220__C (.DIODE(_03812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12141__D (.DIODE(_03812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11883__C (.DIODE(_03812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11882__A2 (.DIODE(_03812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11797__B1 (.DIODE(_03812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11786__A2 (.DIODE(_03812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11703__A (.DIODE(_03812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11308__D (.DIODE(_03812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11306__B1 (.DIODE(_03812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11230__B1 (.DIODE(_03812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12573__B (.DIODE(_03830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12572__A1 (.DIODE(_03830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12569__A1 (.DIODE(_03830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12568__B (.DIODE(_03830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12354__B (.DIODE(_03830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12195__B (.DIODE(_03830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12034__A1 (.DIODE(_03830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11866__A1 (.DIODE(_03830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11702__B (.DIODE(_03830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11248__A1 (.DIODE(_03830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11568__B1 (.DIODE(_03858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11276__C (.DIODE(_03858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13051__B1 (.DIODE(_03869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13011__A1 (.DIODE(_03869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12025__A (.DIODE(_03869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11993__A1 (.DIODE(_03869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11743__A1 (.DIODE(_03869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11659__A1 (.DIODE(_03869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11577__A1 (.DIODE(_03869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11422__A (.DIODE(_03869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11362__A (.DIODE(_03869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11287__A (.DIODE(_03869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12761__A (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12502__B2 (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12347__B2 (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12219__B2 (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12140__B2 (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12026__B2 (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11889__B2 (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11484__B2 (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11344__B2 (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11291__A (.DIODE(_03872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12858__A1 (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12761__B (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12502__A1 (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12347__A1 (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12219__A1 (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12140__A1 (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12026__A1 (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11889__A1 (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11484__A1 (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11291__B (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__B1 (.DIODE(_03876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11294__C (.DIODE(_03876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12141__C (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12140__A2 (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11972__A (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11881__B (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11797__A2 (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11721__D (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11385__D (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11383__B1 (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11313__D (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11312__B1 (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11350__B1 (.DIODE(_03930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11348__C (.DIODE(_03930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11589__A (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11588__A1 (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11454__C1 (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11450__A1 (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11381__A (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11589__B (.DIODE(_03941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11588__A2 (.DIODE(_03941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11381__B (.DIODE(_03941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13060__A (.DIODE(_03942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12970__A (.DIODE(_03942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12784__A (.DIODE(_03942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12779__A (.DIODE(_03942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12650__A (.DIODE(_03942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12157__A (.DIODE(_03942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12050__A (.DIODE(_03942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11995__A1 (.DIODE(_03942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11441__A (.DIODE(_03942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11360__A (.DIODE(_03942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13065__B (.DIODE(_03943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13064__A1 (.DIODE(_03943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12528__A1 (.DIODE(_03943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12375__A1 (.DIODE(_03943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11909__A1 (.DIODE(_03943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11824__A1 (.DIODE(_03943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11747__A1 (.DIODE(_03943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11663__A1 (.DIODE(_03943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11498__A (.DIODE(_03943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11361__A (.DIODE(_03943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13063__A (.DIODE(_03944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12833__A1 (.DIODE(_03944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12808__A1 (.DIODE(_03944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12662__A1 (.DIODE(_03944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12469__A1 (.DIODE(_03944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12319__A1 (.DIODE(_03944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12053__A1 (.DIODE(_03944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11581__A1 (.DIODE(_03944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11438__A1 (.DIODE(_03944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11369__A1 (.DIODE(_03944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12783__A1 (.DIODE(_03945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12778__A1 (.DIODE(_03945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12759__A (.DIODE(_03945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12643__A1 (.DIODE(_03945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12524__A1 (.DIODE(_03945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12371__A1 (.DIODE(_03945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12235__A1 (.DIODE(_03945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11440__A1 (.DIODE(_03945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11372__A1 (.DIODE(_03945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11363__A1 (.DIODE(_03945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12971__A1 (.DIODE(_03947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12871__A (.DIODE(_03947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12812__A (.DIODE(_03947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12527__A (.DIODE(_03947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12468__A (.DIODE(_03947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12374__A (.DIODE(_03947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12238__A (.DIODE(_03947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11908__A (.DIODE(_03947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11665__A1 (.DIODE(_03947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11368__A (.DIODE(_03947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12936__A1 (.DIODE(_03948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12869__A (.DIODE(_03948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12644__A (.DIODE(_03948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12525__A (.DIODE(_03948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12372__A (.DIODE(_03948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12236__A (.DIODE(_03948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11994__A (.DIODE(_03948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11906__A (.DIODE(_03948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11373__A (.DIODE(_03948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11366__A (.DIODE(_03948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11452__B (.DIODE(_03953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11379__A (.DIODE(_03953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12813__A1 (.DIODE(_03954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12786__A (.DIODE(_03954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12781__A (.DIODE(_03954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12646__A (.DIODE(_03954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12522__A1 (.DIODE(_03954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12370__A1 (.DIODE(_03954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11997__A (.DIODE(_03954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11911__A1 (.DIODE(_03954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11443__A (.DIODE(_03954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11375__A (.DIODE(_03954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12874__A1 (.DIODE(_03959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12835__A1 (.DIODE(_03959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12787__A1 (.DIODE(_03959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12653__A1 (.DIODE(_03959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12241__A1 (.DIODE(_03959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12162__A1 (.DIODE(_03959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12048__A1 (.DIODE(_03959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11502__A (.DIODE(_03959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11444__A1 (.DIODE(_03959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11377__A1 (.DIODE(_03959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11428__B1 (.DIODE(_04009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11427__C (.DIODE(_04009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11513__C1 (.DIODE(_04019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11512__A1 (.DIODE(_04019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11458__A (.DIODE(_04019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11449__A (.DIODE(_04019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11448__A1 (.DIODE(_04019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11456__B (.DIODE(_04022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11446__A (.DIODE(_04022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11489__B1 (.DIODE(_04070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11488__C (.DIODE(_04070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19783__A1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19450__A1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13591__A1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13588__A1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12872__A1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12782__A1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12647__A1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12239__A1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12160__A1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11499__A1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13175__A (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11508__A (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13175__B_N (.DIODE(_04090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11508__B (.DIODE(_04090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12213__C (.DIODE(_04102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12212__A2 (.DIODE(_04102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12134__D (.DIODE(_04102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11866__B1 (.DIODE(_04102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11862__A (.DIODE(_04102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11770__B (.DIODE(_04102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11693__A2 (.DIODE(_04102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11692__C (.DIODE(_04102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11611__B1 (.DIODE(_04102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11520__D (.DIODE(_04102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11650__B1 (.DIODE(_04147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11565__C (.DIODE(_04147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11570__B1 (.DIODE(_04150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11569__B (.DIODE(_04150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11671__A (.DIODE(_04158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11670__A1 (.DIODE(_04158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11593__C1 (.DIODE(_04158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11590__A1 (.DIODE(_04158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11587__A (.DIODE(_04158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11671__B (.DIODE(_04159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11670__A2 (.DIODE(_04159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11587__B (.DIODE(_04159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11591__A_N (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11585__A (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12293__C (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12212__B1 (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12034__A2 (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11950__A (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11850__B (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11771__A2 (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11693__B1 (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11692__D (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11606__B1 (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11603__D (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11740__A1 (.DIODE(_04215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11658__C1 (.DIODE(_04215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11657__A1 (.DIODE(_04215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11655__A (.DIODE(_04215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11734__B1 (.DIODE(_04229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11647__C (.DIODE(_04229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11674__A_N (.DIODE(_04247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11667__A (.DIODE(_04247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12340__A2 (.DIODE(_04270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12293__D (.DIODE(_04270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12118__A2 (.DIODE(_04270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12116__C (.DIODE(_04270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12034__B1 (.DIODE(_04270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11937__A (.DIODE(_04270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11852__C (.DIODE(_04270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11851__A2 (.DIODE(_04270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11771__B1 (.DIODE(_04270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11688__B1 (.DIODE(_04270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12662__A2 (.DIODE(_04286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12650__B (.DIODE(_04286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12471__A2 (.DIODE(_04286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12465__A2 (.DIODE(_04286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12448__B (.DIODE(_04286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12374__B (.DIODE(_04286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12219__A2 (.DIODE(_04286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12140__B1 (.DIODE(_04286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11967__B (.DIODE(_04286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11705__B (.DIODE(_04286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11757__B (.DIODE(_04331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11751__A (.DIODE(_04331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12443__C (.DIODE(_04346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12340__B1 (.DIODE(_04346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12276__B (.DIODE(_04346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12196__A2 (.DIODE(_04346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12195__C (.DIODE(_04346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12118__B1 (.DIODE(_04346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12116__D (.DIODE(_04346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11852__D (.DIODE(_04346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11851__B1 (.DIODE(_04346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11764__D (.DIODE(_04346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12450__C (.DIODE(_04444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12449__A2 (.DIODE(_04444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12348__D (.DIODE(_04444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12347__B1 (.DIODE(_04444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12295__A2 (.DIODE(_04444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12211__B (.DIODE(_04444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12020__D (.DIODE(_04444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12019__B1 (.DIODE(_04444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11952__A (.DIODE(_04444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11863__C (.DIODE(_04444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12503__C (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12502__A2 (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12450__D (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12449__B1 (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12291__B (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12133__B1 (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12033__A (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11953__A2 (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11951__C (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11863__D (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12348__C (.DIODE(_04447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12347__A2 (.DIODE(_04447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12300__D (.DIODE(_04447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12299__B1 (.DIODE(_04447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12132__B (.DIODE(_04447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12020__C (.DIODE(_04447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12019__A2 (.DIODE(_04447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11970__D (.DIODE(_04447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11969__B1 (.DIODE(_04447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11865__A (.DIODE(_04447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12833__A2 (.DIODE(_04448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12810__B (.DIODE(_04448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12664__A2 (.DIODE(_04448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12649__A2 (.DIODE(_04448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12613__B (.DIODE(_04448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12538__A2 (.DIODE(_04448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12527__B (.DIODE(_04448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12421__B (.DIODE(_04448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11957__A2 (.DIODE(_04448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11867__B (.DIODE(_04448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12924__B (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12592__A2 (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12590__C (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12494__A (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12493__B1 (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12354__C (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12040__D (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12039__B1 (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11933__B1 (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11930__D (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12590__D (.DIODE(_04517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12427__A2 (.DIODE(_04517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12355__B1 (.DIODE(_04517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12354__D (.DIODE(_04517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12185__C (.DIODE(_04517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12108__D (.DIODE(_04517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12107__B1 (.DIODE(_04517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12064__B1 (.DIODE(_04517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12060__A (.DIODE(_04517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11935__D (.DIODE(_04517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12614__A (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12603__C (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12602__A2 (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12441__B (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12341__C (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12292__B1 (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12281__A2 (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12197__B (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12032__D (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11938__B (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12761__C (.DIODE(_04522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12760__A2 (.DIODE(_04522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12603__D (.DIODE(_04522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12601__A (.DIODE(_04522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12492__B (.DIODE(_04522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12442__A2 (.DIODE(_04522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12341__D (.DIODE(_04522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12038__B (.DIODE(_04522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11942__C (.DIODE(_04522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11940__A2 (.DIODE(_04522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12894__B (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12761__D (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12744__A (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12591__B (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12495__C (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12493__A2 (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12442__B1 (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12431__A2 (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12356__B (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11942__D (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12503__D (.DIODE(_04533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12501__A (.DIODE(_04533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12445__A2 (.DIODE(_04533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12339__B (.DIODE(_04533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12292__A2 (.DIODE(_04533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12213__D (.DIODE(_04533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12117__B (.DIODE(_04533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12032__C (.DIODE(_04533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11953__B1 (.DIODE(_04533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11951__D (.DIODE(_04533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12808__A2 (.DIODE(_04535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12784__B (.DIODE(_04535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12653__A2 (.DIODE(_04535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12652__B (.DIODE(_04535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12643__A2 (.DIODE(_04535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12600__B (.DIODE(_04535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12577__A2_N (.DIODE(_04535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12537__D (.DIODE(_04535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12037__A2 (.DIODE(_04535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11954__B (.DIODE(_04535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12647__A2 (.DIODE(_04551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12644__B (.DIODE(_04551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12524__A2 (.DIODE(_04551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12522__A2 (.DIODE(_04551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12500__B (.DIODE(_04551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12468__B (.DIODE(_04551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12219__B1 (.DIODE(_04551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12136__A2 (.DIODE(_04551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11970__C (.DIODE(_04551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11969__A2 (.DIODE(_04551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12528__A2 (.DIODE(_04555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12525__B (.DIODE(_04555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12371__A2 (.DIODE(_04555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12370__A2 (.DIODE(_04555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12346__B (.DIODE(_04555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12318__B (.DIODE(_04555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12049__B2 (.DIODE(_04555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12027__A1 (.DIODE(_04555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12026__B1 (.DIODE(_04555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11973__A2 (.DIODE(_04555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12009__A_N (.DIODE(_04582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12002__A (.DIODE(_04582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12835__A2 (.DIODE(_04616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12809__A2 (.DIODE(_04616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12782__A2 (.DIODE(_04616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12779__B (.DIODE(_04616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12759__B (.DIODE(_04616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12646__B (.DIODE(_04616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12565__A2 (.DIODE(_04616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12563__C (.DIODE(_04616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12122__A2 (.DIODE(_04616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12035__B (.DIODE(_04616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12964__B (.DIODE(_04643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12859__C (.DIODE(_04643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12858__A2 (.DIODE(_04643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12732__B1 (.DIODE(_04643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12595__C (.DIODE(_04643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12594__A2 (.DIODE(_04643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12592__B1 (.DIODE(_04643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12580__A (.DIODE(_04643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12513__A2 (.DIODE(_04643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12061__D (.DIODE(_04643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12896__C (.DIODE(_04681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12738__C (.DIODE(_04681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12595__D (.DIODE(_04681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12512__C (.DIODE(_04681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12509__A (.DIODE(_04681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12427__B1 (.DIODE(_04681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12186__B1 (.DIODE(_04681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12185__D (.DIODE(_04681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12102__B1 (.DIODE(_04681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12099__D (.DIODE(_04681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12926__C (.DIODE(_04686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12896__D (.DIODE(_04686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12738__D (.DIODE(_04686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12723__C (.DIODE(_04686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12569__A2 (.DIODE(_04686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12568__C (.DIODE(_04686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12512__D (.DIODE(_04686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12510__A (.DIODE(_04686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12362__C (.DIODE(_04686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12104__D (.DIODE(_04686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12306__B1 (.DIODE(_04805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12223__C (.DIODE(_04805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12228__B1 (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12227__B (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12353__B1 (.DIODE(_04885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12303__C (.DIODE(_04885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12926__D (.DIODE(_04944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12720__A2 (.DIODE(_04944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12573__C (.DIODE(_04944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12572__A2 (.DIODE(_04944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12569__B1 (.DIODE(_04944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12568__D (.DIODE(_04944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12535__A (.DIODE(_04944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12515__C (.DIODE(_04944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12418__C (.DIODE(_04944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12362__D (.DIODE(_04944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12966__D (.DIODE(_04967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12965__B1 (.DIODE(_04967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12854__D (.DIODE(_04967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12720__B1 (.DIODE(_04967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12719__D (.DIODE(_04967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12573__D (.DIODE(_04967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12572__B1 (.DIODE(_04967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12562__A (.DIODE(_04967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12536__B1 (.DIODE(_04967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12385__B1 (.DIODE(_04967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12497__A1 (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12491__A (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12444__B1_N (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12447__B1 (.DIODE(_05027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12446__B (.DIODE(_05027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12508__B1 (.DIODE(_05035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12453__C (.DIODE(_05035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12553__A1 (.DIODE(_05044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12552__C1 (.DIODE(_05044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12464__B1 (.DIODE(_05044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12463__A2 (.DIODE(_05044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12996__B (.DIODE(_05077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12994__B (.DIODE(_05077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12943__B (.DIODE(_05077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12908__B (.DIODE(_05077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12755__B (.DIODE(_05077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12745__B1 (.DIODE(_05077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12732__A2 (.DIODE(_05077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12731__C (.DIODE(_05077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12596__A2 (.DIODE(_05077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12495__D (.DIODE(_05077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12872__A2 (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12869__B (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12813__A2 (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12812__B (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12783__A2 (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12767__B (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12743__B (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12616__C (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12615__A2 (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12502__B1 (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12549__B1 (.DIODE(_05090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12548__A (.DIODE(_05090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12521__A1 (.DIODE(_05090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12542__B1 (.DIODE(_05096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12541__A (.DIODE(_05096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12518__A1 (.DIODE(_05096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13030__C (.DIODE(_05118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12966__C (.DIODE(_05118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12965__A2 (.DIODE(_05118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12925__B1 (.DIODE(_05118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12854__C (.DIODE(_05118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12724__B1 (.DIODE(_05118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12723__D (.DIODE(_05118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12719__C (.DIODE(_05118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12709__A (.DIODE(_05118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12536__A2 (.DIODE(_05118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12631__A1 (.DIODE(_05126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12630__C1 (.DIODE(_05126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12547__B1 (.DIODE(_05126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12546__A2 (.DIODE(_05126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12545__A2 (.DIODE(_05126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12553__C1 (.DIODE(_05128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12552__A1 (.DIODE(_05128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12661__A1 (.DIODE(_05133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12660__C1 (.DIODE(_05133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12553__B1 (.DIODE(_05133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12552__A2 (.DIODE(_05133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13050__B (.DIODE(_05145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13049__A_N (.DIODE(_05145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13035__D (.DIODE(_05145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13011__B1 (.DIODE(_05145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12993__D (.DIODE(_05145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12892__B1 (.DIODE(_05145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12711__B1 (.DIODE(_05145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12710__D (.DIODE(_05145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12564__A (.DIODE(_05145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12563__D (.DIODE(_05145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12627__A (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12579__A (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12566__A (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13591__A2 (.DIODE(_05147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13065__D (.DIODE(_05147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13059__B1 (.DIODE(_05147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13047__B1 (.DIODE(_05147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13046__A (.DIODE(_05147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12957__A2 (.DIODE(_05147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12929__B (.DIODE(_05147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12850__B1 (.DIODE(_05147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12715__D (.DIODE(_05147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12565__B1 (.DIODE(_05147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12627__B (.DIODE(_05161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12579__B (.DIODE(_05161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13033__A2 (.DIODE(_05163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13017__C (.DIODE(_05163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12983__A2 (.DIODE(_05163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12958__B (.DIODE(_05163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12934__B (.DIODE(_05163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12778__B2 (.DIODE(_05163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12754__A2 (.DIODE(_05163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12737__B (.DIODE(_05163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12733__A1 (.DIODE(_05163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12581__B (.DIODE(_05163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13047__A2 (.DIODE(_05167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13035__C (.DIODE(_05167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13011__A2 (.DIODE(_05167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13009__A2 (.DIODE(_05167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13008__B (.DIODE(_05167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12990__B (.DIODE(_05167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12986__B (.DIODE(_05167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12971__A2 (.DIODE(_05167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12726__A2_N (.DIODE(_05167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12585__A2 (.DIODE(_05167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12609__B1_N (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12597__A1 (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12593__A (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12937__B (.DIODE(_05184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12936__A2 (.DIODE(_05184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12874__A2 (.DIODE(_05184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12868__A2 (.DIODE(_05184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12857__B (.DIODE(_05184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12850__A2 (.DIODE(_05184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12781__B (.DIODE(_05184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12715__C (.DIODE(_05184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12610__A2 (.DIODE(_05184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12602__B1 (.DIODE(_05184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12911__C1 (.DIODE(_05197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12910__A2 (.DIODE(_05197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12787__A2 (.DIODE(_05197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12786__B (.DIODE(_05197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12778__A2 (.DIODE(_05197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12730__B (.DIODE(_05197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12713__A2_N (.DIODE(_05197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12712__D (.DIODE(_05197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12616__D (.DIODE(_05197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12615__B1 (.DIODE(_05197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12631__A2 (.DIODE(_05212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12630__B1 (.DIODE(_05212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12661__A2 (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12660__B1 (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13458__B1 (.DIODE(_05280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12708__A2 (.DIODE(_05280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13588__A2 (.DIODE(_05292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13065__C (.DIODE(_05292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13059__A2 (.DIODE(_05292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13051__A2 (.DIODE(_05292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13033__B1 (.DIODE(_05292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13031__A2 (.DIODE(_05292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13017__D (.DIODE(_05292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12892__A2 (.DIODE(_05292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12711__A2 (.DIODE(_05292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12710__C (.DIODE(_05292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12970__B (.DIODE(_05327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12968__B (.DIODE(_05327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12942__A2 (.DIODE(_05327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12905__A2 (.DIODE(_05327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12902__B (.DIODE(_05327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12871__B (.DIODE(_05327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12783__B2 (.DIODE(_05327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12760__B1 (.DIODE(_05327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12746__A1 (.DIODE(_05327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12745__A2 (.DIODE(_05327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12911__A1 (.DIODE(_05479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12910__B1 (.DIODE(_05479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12909__C (.DIODE(_05479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12898__A2 (.DIODE(_05479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12897__C (.DIODE(_05479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13549__A (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13539__A (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13083__C (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13081__A (.DIODE(_05506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12954__A (.DIODE(_05506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12957__B1 (.DIODE(_05510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12929__C (.DIODE(_05510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12957__B2 (.DIODE(_05511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12929__D (.DIODE(_05511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12955__B (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12952__B (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12951__B (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12985__B1 (.DIODE(_05547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12984__B (.DIODE(_05547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12967__A1 (.DIODE(_05547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12985__A2 (.DIODE(_05548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12984__C (.DIODE(_05548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12967__A2 (.DIODE(_05548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12985__A1 (.DIODE(_05549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12984__A (.DIODE(_05549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12967__B1_N (.DIODE(_05549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13064__A2 (.DIODE(_05575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13063__B (.DIODE(_05575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13060__B (.DIODE(_05575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13054__A1 (.DIODE(_05575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13051__B2 (.DIODE(_05575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13049__C (.DIODE(_05575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13037__A1 (.DIODE(_05575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13015__B (.DIODE(_05575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13010__B (.DIODE(_05575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12997__A2 (.DIODE(_05575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13012__A (.DIODE(_05576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12996__C (.DIODE(_05576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12995__A (.DIODE(_05576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13034__A (.DIODE(_05600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13023__B (.DIODE(_05600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13018__B (.DIODE(_05600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13049__B (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13046__B (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13037__A3 (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13549__B (.DIODE(_05662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13080__A (.DIODE(_05662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13539__B (.DIODE(_05665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13083__D (.DIODE(_05665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13531__B (.DIODE(_05666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13456__A1 (.DIODE(_05666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13115__A1 (.DIODE(_05666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13111__A (.DIODE(_05668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13099__A (.DIODE(_05668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13095__A (.DIODE(_05668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13456__A2 (.DIODE(_05685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13115__A2 (.DIODE(_05685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13456__B1 (.DIODE(_05697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13115__C1 (.DIODE(_05697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13435__B (.DIODE(_05698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13419__A2 (.DIODE(_05698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13191__A2 (.DIODE(_05698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13124__B1 (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13123__A (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13135__A (.DIODE(_05706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13134__A1 (.DIODE(_05706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13130__B1 (.DIODE(_05706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13126__A1 (.DIODE(_05706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13125__B1 (.DIODE(_05706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13130__C1 (.DIODE(_05707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13126__A2 (.DIODE(_05707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13125__C1 (.DIODE(_05707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13142__B_N (.DIODE(_05711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13129__B (.DIODE(_05711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13135__B (.DIODE(_05713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13134__A2 (.DIODE(_05713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13166__A (.DIODE(_05736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13160__A1 (.DIODE(_05736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13158__C (.DIODE(_05739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13157__B1 (.DIODE(_05739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13170__C (.DIODE(_05751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13169__B1 (.DIODE(_05751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13193__B (.DIODE(_05755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13173__B (.DIODE(_05755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13429__A1 (.DIODE(_05774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13425__A1 (.DIODE(_05774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13412__A1 (.DIODE(_05774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13203__A1 (.DIODE(_05774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13429__A2 (.DIODE(_05781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13425__A2 (.DIODE(_05781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13412__A2 (.DIODE(_05781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13203__A2 (.DIODE(_05781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13417__B (.DIODE(_05786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13409__A2 (.DIODE(_05786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13353__A2 (.DIODE(_05786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13418__A (.DIODE(_05929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13409__B1_N (.DIODE(_05929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13352__A (.DIODE(_05929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13403__A1 (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13402__A1 (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13403__A2 (.DIODE(_05974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13402__A2 (.DIODE(_05974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17916__A2 (.DIODE(_05976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13397__A (.DIODE(_05976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17916__A3 (.DIODE(_05978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13397__B (.DIODE(_05978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13400__A (.DIODE(_05980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13592__A2 (.DIODE(_05981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13554__A (.DIODE(_05981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13510__A (.DIODE(_05981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13466__A (.DIODE(_05981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13401__A (.DIODE(_05981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13592__B1 (.DIODE(_05984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13590__B1 (.DIODE(_05984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13547__A (.DIODE(_05984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13504__A (.DIODE(_05984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13404__A (.DIODE(_05984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13424__A1 (.DIODE(_06002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13424__A2 (.DIODE(_06003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13439__D (.DIODE(_06019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13445__C1 (.DIODE(_06021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13591__B1_N (.DIODE(_06035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13552__C_N (.DIODE(_06035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13489__A (.DIODE(_06035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13475__A (.DIODE(_06035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13455__A (.DIODE(_06035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13476__A1 (.DIODE(_06041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13470__B (.DIODE(_06041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13461__A3 (.DIODE(_06041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13464__B (.DIODE(_06044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13468__B (.DIODE(_06047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13472__B (.DIODE(_06050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13476__A2 (.DIODE(_06052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13575__A (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13567__A (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13563__A (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13559__A (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13542__A (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13537__A (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13534__A (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13529__A (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13526__A (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13476__B1 (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13493__A1 (.DIODE(_06055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13488__A2 (.DIODE(_06055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13487__C (.DIODE(_06055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13479__A2_N (.DIODE(_06055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13482__B (.DIODE(_06058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13485__B (.DIODE(_06060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13490__A1 (.DIODE(_06062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13490__A2 (.DIODE(_06063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13589__B1 (.DIODE(_06064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13586__B1 (.DIODE(_06064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13583__B1_N (.DIODE(_06064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13579__B1 (.DIODE(_06064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13571__B1_N (.DIODE(_06064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13556__B1_N (.DIODE(_06064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13545__B_N (.DIODE(_06064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13499__B_N (.DIODE(_06064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13493__B1 (.DIODE(_06064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13490__B1_N (.DIODE(_06064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13493__A2 (.DIODE(_06066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13499__A (.DIODE(_06071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13502__B (.DIODE(_06073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13508__B (.DIODE(_06078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13512__B (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13519__B (.DIODE(_06087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13522__B (.DIODE(_06089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13526__B (.DIODE(_06092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13529__B (.DIODE(_06094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13534__B (.DIODE(_06098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13537__B (.DIODE(_06100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13542__B (.DIODE(_06104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13545__A (.DIODE(_06106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13587__B1 (.DIODE(_06108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13584__B1 (.DIODE(_06108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13580__B1 (.DIODE(_06108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13576__B1 (.DIODE(_06108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13572__B1 (.DIODE(_06108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13568__B1 (.DIODE(_06108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13564__B1 (.DIODE(_06108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13560__B1 (.DIODE(_06108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13557__B1 (.DIODE(_06108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13553__B1 (.DIODE(_06108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13633__S (.DIODE(_06153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13631__S (.DIODE(_06153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13629__S (.DIODE(_06153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13627__S (.DIODE(_06153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13625__S (.DIODE(_06153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13623__S (.DIODE(_06153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13621__S (.DIODE(_06153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13619__S (.DIODE(_06153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13617__S (.DIODE(_06153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13615__S (.DIODE(_06153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13798__S (.DIODE(_06255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13794__S (.DIODE(_06255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13790__S (.DIODE(_06255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13786__S (.DIODE(_06255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13782__S (.DIODE(_06255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13778__S (.DIODE(_06255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13774__S (.DIODE(_06255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13746__A (.DIODE(_06255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13739__A (.DIODE(_06255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13804__S (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13800__S (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13795__S (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13791__S (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13787__S (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13783__S (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13779__S (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13742__A (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13775__S (.DIODE(_06259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13771__S (.DIODE(_06259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13767__S (.DIODE(_06259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13763__S (.DIODE(_06259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13759__S (.DIODE(_06259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13756__A2 (.DIODE(_06259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13755__B1 (.DIODE(_06259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13752__S (.DIODE(_06259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13748__S (.DIODE(_06259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13743__S (.DIODE(_06259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13803__A2 (.DIODE(_06262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13802__B (.DIODE(_06262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13770__S (.DIODE(_06262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13766__S (.DIODE(_06262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13762__S (.DIODE(_06262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13758__S (.DIODE(_06262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13755__A2 (.DIODE(_06262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13754__B (.DIODE(_06262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13751__S (.DIODE(_06262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13747__S (.DIODE(_06262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13865__B (.DIODE(_06354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13854__B_N (.DIODE(_06354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17231__A (.DIODE(_06356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17112__A2 (.DIODE(_06356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17110__A2 (.DIODE(_06356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17108__A2 (.DIODE(_06356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17106__A2 (.DIODE(_06356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17104__A2 (.DIODE(_06356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17102__A2 (.DIODE(_06356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17100__A2 (.DIODE(_06356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17073__A (.DIODE(_06356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13856__A (.DIODE(_06356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17775__A2 (.DIODE(_06357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17772__A2 (.DIODE(_06357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17769__A2 (.DIODE(_06357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17766__A2 (.DIODE(_06357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17762__A2 (.DIODE(_06357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17723__A (.DIODE(_06357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13860__A2 (.DIODE(_06357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17231__B (.DIODE(_06360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13916__C (.DIODE(_06360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13902__A3 (.DIODE(_06360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13861__B (.DIODE(_06360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13914__S (.DIODE(_06361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13911__S (.DIODE(_06361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13907__S (.DIODE(_06361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13901__B (.DIODE(_06361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13896__S (.DIODE(_06361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13892__S (.DIODE(_06361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13883__S (.DIODE(_06361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13866__A (.DIODE(_06361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13863__B1 (.DIODE(_06361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13899__B1 (.DIODE(_06365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13898__B1 (.DIODE(_06365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13889__A2 (.DIODE(_06365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13888__A (.DIODE(_06365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13886__B1 (.DIODE(_06365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13885__B1 (.DIODE(_06365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13879__S (.DIODE(_06365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13875__S (.DIODE(_06365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13871__S (.DIODE(_06365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13867__S (.DIODE(_06365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16416__S (.DIODE(_06403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16408__S (.DIODE(_06403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16403__S (.DIODE(_06403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16394__S (.DIODE(_06403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16290__A (.DIODE(_06403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13920__A (.DIODE(_06403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16427__A2 (.DIODE(_06404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16426__C1 (.DIODE(_06404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16369__A2 (.DIODE(_06404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16368__C1 (.DIODE(_06404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16355__A2 (.DIODE(_06404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16354__C1 (.DIODE(_06404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16326__A2 (.DIODE(_06404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16325__B1 (.DIODE(_06404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15601__A2 (.DIODE(_06404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13927__B1 (.DIODE(_06404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14588__A (.DIODE(_06405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14301__B2 (.DIODE(_06405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14280__B2 (.DIODE(_06405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14022__A (.DIODE(_06405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13977__B2 (.DIODE(_06405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13947__B2 (.DIODE(_06405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13945__A (.DIODE(_06405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13934__B2 (.DIODE(_06405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13933__A (.DIODE(_06405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13922__A (.DIODE(_06405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16305__A (.DIODE(_06406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15597__A (.DIODE(_06406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15583__A1 (.DIODE(_06406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14189__A (.DIODE(_06406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14142__B2 (.DIODE(_06406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14141__A (.DIODE(_06406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14086__B2 (.DIODE(_06406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14085__A (.DIODE(_06406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14023__B2 (.DIODE(_06406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13923__A (.DIODE(_06406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16406__B1 (.DIODE(_06407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16401__B1 (.DIODE(_06407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16392__A (.DIODE(_06407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16333__B1 (.DIODE(_06407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16330__B1 (.DIODE(_06407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16316__B1 (.DIODE(_06407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16295__B1 (.DIODE(_06407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15580__C1 (.DIODE(_06407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13924__A (.DIODE(_06407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16425__B1 (.DIODE(_06408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16415__A1 (.DIODE(_06408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16407__A1 (.DIODE(_06408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16372__B1 (.DIODE(_06408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16367__B (.DIODE(_06408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16359__A1 (.DIODE(_06408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16342__A1 (.DIODE(_06408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16303__B1 (.DIODE(_06408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16299__B2 (.DIODE(_06408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13927__A1 (.DIODE(_06408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14693__C (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14692__A2 (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14222__A2 (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14068__C (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14061__B (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14056__B1 (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14007__B1 (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14005__C (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13985__A (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13926__A (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16283__A1 (.DIODE(_06410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16235__A (.DIODE(_06410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15705__A1 (.DIODE(_06410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15699__A1 (.DIODE(_06410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15676__A1 (.DIODE(_06410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15651__A (.DIODE(_06410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15629__B1 (.DIODE(_06410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15628__A (.DIODE(_06410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13927__A2 (.DIODE(_06410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14518__B2 (.DIODE(_06412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14301__A1 (.DIODE(_06412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14280__A1 (.DIODE(_06412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14190__A (.DIODE(_06412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14021__A (.DIODE(_06412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13977__A1 (.DIODE(_06412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13947__A1 (.DIODE(_06412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13945__B (.DIODE(_06412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13934__A1 (.DIODE(_06412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13933__B (.DIODE(_06412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15659__A1 (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15610__A2 (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15027__A (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14950__C (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14686__A2 (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14624__B (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14308__D (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13977__B1 (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13976__D (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13930__A (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14951__A2 (.DIODE(_06414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14884__A2 (.DIODE(_06414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14824__B1 (.DIODE(_06414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14556__B (.DIODE(_06414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14431__B1 (.DIODE(_06414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14430__D (.DIODE(_06414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14307__B1 (.DIODE(_06414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13948__A (.DIODE(_06414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13934__A2 (.DIODE(_06414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13933__C (.DIODE(_06414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15683__A1 (.DIODE(_06415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15028__B1 (.DIODE(_06415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15027__B (.DIODE(_06415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14882__A2 (.DIODE(_06415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14767__B (.DIODE(_06415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14686__B1 (.DIODE(_06415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14623__A2 (.DIODE(_06415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14622__C (.DIODE(_06415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14567__B (.DIODE(_06415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13932__A (.DIODE(_06415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14951__B1 (.DIODE(_06416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14950__D (.DIODE(_06416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14881__C (.DIODE(_06416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14286__A (.DIODE(_06416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14236__C (.DIODE(_06416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14235__A2 (.DIODE(_06416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13947__A2 (.DIODE(_06416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13945__C (.DIODE(_06416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13934__B1 (.DIODE(_06416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13933__D (.DIODE(_06416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14506__A (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14333__A1_N (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14303__A1_N (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14282__A1_N (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14025__A (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14024__C (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13980__A (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13949__C (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13941__A1_N (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13940__C (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15610__A1 (.DIODE(_06421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14894__B1 (.DIODE(_06421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14824__A2 (.DIODE(_06421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14687__B (.DIODE(_06421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14561__B1 (.DIODE(_06421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14308__C (.DIODE(_06421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14240__D (.DIODE(_06421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13977__A2 (.DIODE(_06421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13976__C (.DIODE(_06421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13938__A (.DIODE(_06421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15641__A1 (.DIODE(_06422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14952__B (.DIODE(_06422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14893__D (.DIODE(_06422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14431__A2 (.DIODE(_06422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14430__C (.DIODE(_06422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14338__D (.DIODE(_06422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14307__A2 (.DIODE(_06422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14242__B1 (.DIODE(_06422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14022__D (.DIODE(_06422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13939__A (.DIODE(_06422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17183__A1 (.DIODE(_06423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15691__A2 (.DIODE(_06423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14723__B (.DIODE(_06423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14649__B (.DIODE(_06423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14575__B (.DIODE(_06423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14337__B1 (.DIODE(_06423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14290__B (.DIODE(_06423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14023__B1 (.DIODE(_06423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13941__A2_N (.DIODE(_06423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13940__D (.DIODE(_06423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15118__A2 (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15083__B1 (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14882__B1 (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14766__A2 (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14765__C (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14622__D (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14566__A2 (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14546__B (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14421__C (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13944__A (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15026__B (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14881__D (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14674__B (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14623__B1 (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14565__C (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14301__A2 (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14300__C (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14236__D (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13946__A (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13945__D (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17195__A1 (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15383__A2 (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15104__B (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15096__B (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14942__B (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14420__A2 (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14282__A2_N (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14281__D (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14235__B1 (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13947__B1 (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17187__A1 (.DIODE(_06432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14883__B (.DIODE(_06432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14851__A2 (.DIODE(_06432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14843__B (.DIODE(_06432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14333__A2_N (.DIODE(_06432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14288__C (.DIODE(_06432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14287__A2 (.DIODE(_06432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14276__B (.DIODE(_06432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14238__A2 (.DIODE(_06432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13949__D (.DIODE(_06432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15010__B2 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14800__A (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14420__A1 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14338__B (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14337__A1 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14307__A1 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14236__B (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14235__A1 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13987__A (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13961__A1 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15627__B (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14967__A2 (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14966__C (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14629__B1 (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14573__A2 (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14572__C (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14448__B1 (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14228__C (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13964__C (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13957__A (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14896__A2 (.DIODE(_06441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14895__B (.DIODE(_06441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14695__B (.DIODE(_06441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14319__B1 (.DIODE(_06441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14318__D (.DIODE(_06441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14243__D (.DIODE(_06441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14231__A2 (.DIODE(_06441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14085__C (.DIODE(_06441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13989__A (.DIODE(_06441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13961__A2 (.DIODE(_06441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15637__B1 (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14967__B1 (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14966__D (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14894__A2 (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14730__B (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14573__B1 (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14561__A2 (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14240__C (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13964__D (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13959__A (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14893__C (.DIODE(_06443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14574__A1 (.DIODE(_06443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14338__C (.DIODE(_06443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14242__A2 (.DIODE(_06443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14231__B1 (.DIODE(_06443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14228__D (.DIODE(_06443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14085__D (.DIODE(_06443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14022__C (.DIODE(_06443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13979__A (.DIODE(_06443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13961__B1 (.DIODE(_06443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14661__B2 (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14420__B2 (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14338__A (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14337__B2 (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14307__B2 (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14236__A (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14235__B2 (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13992__A (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13990__A (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13961__B2 (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14940__B2 (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14939__A (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14870__A (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14869__B2 (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14754__B2 (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14493__A (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14492__B2 (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14421__A (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14308__A (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13964__A (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14940__A1 (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14939__B (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14870__B (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14869__A1 (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14754__A1 (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14661__A1 (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14492__A1 (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14421__B (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14308__B (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13964__B (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14012__B1 (.DIODE(_06448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13965__B (.DIODE(_06448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15010__A1 (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14880__A1 (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14872__A (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14757__A (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14676__A1 (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14664__A (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14599__A (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14494__A1 (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13984__A (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13967__A (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19545__A1 (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19107__A1 (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14341__A (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14340__A1 (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14290__A (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14238__A1 (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14131__A1 (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14097__A1 (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14042__A1 (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13971__A (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15627__A (.DIODE(_06452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14693__D (.DIODE(_06452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14692__B1 (.DIODE(_06452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14630__A1 (.DIODE(_06452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14629__A2 (.DIODE(_06452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14448__A2 (.DIODE(_06452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14447__C (.DIODE(_06452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14318__C (.DIODE(_06452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14222__B1 (.DIODE(_06452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13969__A (.DIODE(_06452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15646__A (.DIODE(_06453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15396__A2 (.DIODE(_06453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14969__B (.DIODE(_06453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14735__B (.DIODE(_06453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14451__A1 (.DIODE(_06453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14349__B1 (.DIODE(_06453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14319__A2 (.DIODE(_06453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13992__C (.DIODE(_06453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13988__A (.DIODE(_06453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13970__A (.DIODE(_06453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15828__A2 (.DIODE(_06454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15827__A2 (.DIODE(_06454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15727__B (.DIODE(_06454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15726__A_N (.DIODE(_06454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15624__B1 (.DIODE(_06454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15613__A1 (.DIODE(_06454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14188__A (.DIODE(_06454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14088__A2_N (.DIODE(_06454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14087__D (.DIODE(_06454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13971__B (.DIODE(_06454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15855__A1 (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15624__A2 (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14631__B (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14432__B (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14337__A2 (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14310__B (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14086__B1 (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14029__A (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14023__A2 (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13980__B (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15383__A1 (.DIODE(_06468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15057__A (.DIODE(_06468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14942__A (.DIODE(_06468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14809__A (.DIODE(_06468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14435__A1 (.DIODE(_06468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14424__A (.DIODE(_06468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14310__A (.DIODE(_06468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14276__A (.DIODE(_06468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14012__A1 (.DIODE(_06468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13986__A (.DIODE(_06468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14450__A2 (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14349__A2 (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14081__C (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14066__B1 (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14058__B (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14041__A (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14033__A2 (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14032__B (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14010__B (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13986__B (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19549__A1 (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19111__A1 (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14288__B (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14287__A1 (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14082__A2 (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14081__B (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14033__A1 (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14032__A (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13992__B (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13991__A1 (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15636__A (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14348__A (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14233__B (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14223__A (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14142__A2 (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14141__C (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14033__B1 (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14032__C (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14012__A2 (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13991__A2 (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15646__B (.DIODE(_06473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15624__A1 (.DIODE(_06473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14436__A2_N (.DIODE(_06473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14142__B1 (.DIODE(_06473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14141__D (.DIODE(_06473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14086__A2 (.DIODE(_06473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14026__A (.DIODE(_06473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14024__D (.DIODE(_06473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13992__D (.DIODE(_06473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13991__B1 (.DIODE(_06473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19552__A1 (.DIODE(_06474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19114__A1 (.DIODE(_06474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14288__A (.DIODE(_06474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14287__B2 (.DIODE(_06474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14096__A (.DIODE(_06474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14082__A1 (.DIODE(_06474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14081__A (.DIODE(_06474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14034__A1 (.DIODE(_06474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14033__B2 (.DIODE(_06474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13991__B2 (.DIODE(_06474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15145__A1_N (.DIODE(_06484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15062__C (.DIODE(_06484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15058__A1_N (.DIODE(_06484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15006__C (.DIODE(_06484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15002__A (.DIODE(_06484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14767__A (.DIODE(_06484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14674__A (.DIODE(_06484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14609__A (.DIODE(_06484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14483__A (.DIODE(_06484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14001__A (.DIODE(_06484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15147__B (.DIODE(_06485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14952__A (.DIODE(_06485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14884__A1 (.DIODE(_06485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14883__A (.DIODE(_06485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14799__A1 (.DIODE(_06485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14501__A (.DIODE(_06485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14432__A (.DIODE(_06485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14243__C (.DIODE(_06485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14010__A (.DIODE(_06485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14002__A (.DIODE(_06485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19536__A1 (.DIODE(_06486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19099__A1 (.DIODE(_06486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15242__A (.DIODE(_06486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15206__A1 (.DIODE(_06486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14806__A1 (.DIODE(_06486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14436__A1_N (.DIODE(_06486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14346__A1 (.DIODE(_06486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14316__A1 (.DIODE(_06486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14233__A (.DIODE(_06486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14009__A1 (.DIODE(_06486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14950__A (.DIODE(_06487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14882__B2 (.DIODE(_06487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14881__A (.DIODE(_06487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14766__B2 (.DIODE(_06487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14499__A (.DIODE(_06487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14484__B2 (.DIODE(_06487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14240__A (.DIODE(_06487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14228__A (.DIODE(_06487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14007__A1 (.DIODE(_06487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14005__A (.DIODE(_06487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15061__A1 (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14765__B (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14673__A1 (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14672__B (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14608__A1 (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14500__A1 (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14499__B (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14484__A1 (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14482__B (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14005__B (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14378__A2 (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14348__B (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14009__B1 (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14008__A (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14950__B (.DIODE(_06490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14882__A1 (.DIODE(_06490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14881__B (.DIODE(_06490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14766__A1 (.DIODE(_06490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14430__B (.DIODE(_06490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14241__A (.DIODE(_06490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14240__B (.DIODE(_06490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14231__A1 (.DIODE(_06490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14228__B (.DIODE(_06490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14007__A2 (.DIODE(_06490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14136__A (.DIODE(_06493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14135__A (.DIODE(_06493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14102__A (.DIODE(_06493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14101__A (.DIODE(_06493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14045__A (.DIODE(_06493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14044__A (.DIODE(_06493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14017__A (.DIODE(_06493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14016__A (.DIODE(_06493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15501__B1 (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14380__A (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14133__A (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14132__A (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14107__A1 (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14099__A (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14098__A (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14043__A (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14014__A (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14013__A (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19558__A1 (.DIODE(_06505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19121__A1 (.DIODE(_06505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15579__A (.DIODE(_06505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14191__A (.DIODE(_06505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14142__A1 (.DIODE(_06505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14141__B (.DIODE(_06505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14086__A1 (.DIODE(_06505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14085__B (.DIODE(_06505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14023__A1 (.DIODE(_06505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14022__B (.DIODE(_06505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19555__A1 (.DIODE(_06509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19118__A1 (.DIODE(_06509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15579__B (.DIODE(_06509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14191__B (.DIODE(_06509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14187__A1 (.DIODE(_06509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14140__A (.DIODE(_06509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14088__A1_N (.DIODE(_06509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14087__C (.DIODE(_06509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14030__A1 (.DIODE(_06509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14027__A1_N (.DIODE(_06509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17173__A1 (.DIODE(_06510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15827__B1_N (.DIODE(_06510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15706__A1 (.DIODE(_06510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15625__A1 (.DIODE(_06510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14923__B (.DIODE(_06510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14788__B (.DIODE(_06510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14785__B (.DIODE(_06510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14341__B (.DIODE(_06510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14340__A2 (.DIODE(_06510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14027__A2_N (.DIODE(_06510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17179__A1 (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15824__A1 (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15706__A2 (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15691__A1 (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15625__A2 (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14726__B (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14717__B (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14712__A2 (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14645__A1_N (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14030__A2 (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15828__A1 (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15827__A1 (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15623__A1 (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14346__A2 (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14192__A (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14140__B (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14116__A (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14097__A2 (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14082__B1 (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14042__A2 (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15228__B2 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15185__B2 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15126__B2 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15118__B2 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15081__A (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15028__B2 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14693__A (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14573__B2 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14572__A (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14056__A1 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15228__A1 (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15185__A1 (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15126__A1 (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15118__A1 (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15081__B (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15028__A1 (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14693__B (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14573__A1 (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14572__B (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14056__A2 (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15398__A (.DIODE(_06543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14973__A (.DIODE(_06543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14455__A1 (.DIODE(_06543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14227__A1 (.DIODE(_06543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14073__A (.DIODE(_06543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14071__A1 (.DIODE(_06543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15261__A1 (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15224__B (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15131__A1 (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14815__A1 (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14687__A (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14624__A (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14567__A (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14550__A (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14067__A (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14061__A (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15192__B2 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15133__B2 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15114__A (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15113__B2 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15076__A (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15075__B2 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14729__B2 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14685__A (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14545__A (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14063__A (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19533__A1 (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19095__A1 (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14894__B2 (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14893__A (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14565__A (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14552__A (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14448__B2 (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14222__B2 (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14068__A (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14066__A1 (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15193__B (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15192__A1 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15114__B (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15113__A1 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15075__A1 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14729__A1 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14685__B (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14547__A1 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14545__B (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14065__A (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19530__A1 (.DIODE(_06549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19093__A1 (.DIODE(_06549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15261__B2 (.DIODE(_06549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15224__A (.DIODE(_06549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14894__A1 (.DIODE(_06549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14893__B (.DIODE(_06549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14565__B (.DIODE(_06549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14222__A1 (.DIODE(_06549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14068__B (.DIODE(_06549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14066__A2 (.DIODE(_06549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19527__A1 (.DIODE(_06551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19090__A1 (.DIODE(_06551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15396__A1 (.DIODE(_06551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15320__A1 (.DIODE(_06551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15285__A (.DIODE(_06551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14969__A (.DIODE(_06551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14896__A1 (.DIODE(_06551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14895__A (.DIODE(_06551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14450__A1 (.DIODE(_06551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14069__A (.DIODE(_06551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15510__A1 (.DIODE(_06555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15504__A (.DIODE(_06555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14395__A1 (.DIODE(_06555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14362__A (.DIODE(_06555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14072__A (.DIODE(_06555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15574__A1 (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15527__A1 (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14389__A (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14210__A1 (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14185__A (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14167__A1 (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14159__A (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14124__A1 (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14109__A (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14077__A (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15503__A (.DIODE(_06557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14388__A (.DIODE(_06557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14361__A (.DIODE(_06557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14183__A (.DIODE(_06557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14182__B1 (.DIODE(_06557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14157__A (.DIODE(_06557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14156__B1 (.DIODE(_06557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14108__A (.DIODE(_06557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14075__A (.DIODE(_06557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14074__B1 (.DIODE(_06557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15308__A (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15211__A (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15173__A (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15163__A (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15096__A (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15042__A (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14843__A (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14716__A (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14649__A (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14117__A (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15976__A (.DIODE(_06600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15974__A1 (.DIODE(_06600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15943__A (.DIODE(_06600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15805__A (.DIODE(_06600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15672__A1 (.DIODE(_06600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15621__A1 (.DIODE(_06600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15581__A (.DIODE(_06600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14187__A2 (.DIODE(_06600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14131__A2 (.DIODE(_06600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14117__B (.DIODE(_06600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15512__A (.DIODE(_06601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15460__A (.DIODE(_06601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15427__A (.DIODE(_06601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15406__A (.DIODE(_06601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14983__A (.DIODE(_06601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14469__A (.DIODE(_06601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14118__A (.DIODE(_06601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15532__A (.DIODE(_06602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15531__A (.DIODE(_06602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15513__A (.DIODE(_06602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15439__A (.DIODE(_06602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15378__A (.DIODE(_06602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14400__A (.DIODE(_06602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14399__A (.DIODE(_06602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14368__A (.DIODE(_06602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14251__A (.DIODE(_06602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14119__A (.DIODE(_06602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15593__A (.DIODE(_06603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15589__A1 (.DIODE(_06603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15469__A (.DIODE(_06603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15465__A (.DIODE(_06603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14476__A1 (.DIODE(_06603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14219__A1 (.DIODE(_06603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14214__A (.DIODE(_06603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14176__A1 (.DIODE(_06603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14172__A (.DIODE(_06603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14128__A (.DIODE(_06603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15329__A1 (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15317__A1 (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15283__A (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15259__A (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14822__A (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14735__A (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14695__A (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14631__A (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14575__A (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14121__A (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19521__A1 (.DIODE(_06605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19084__A1 (.DIODE(_06605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15341__A (.DIODE(_06605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15333__A (.DIODE(_06605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15307__A1 (.DIODE(_06605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15140__A1 (.DIODE(_06605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14912__A (.DIODE(_06605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14785__A (.DIODE(_06605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14712__A1 (.DIODE(_06605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14122__A1 (.DIODE(_06605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15459__A (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15426__A (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15377__A (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14982__A (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14397__A (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14396__A (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14123__A (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15529__A (.DIODE(_06607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15528__A (.DIODE(_06607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15511__A (.DIODE(_06607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15376__A (.DIODE(_06607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14468__A (.DIODE(_06607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14250__A (.DIODE(_06607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14169__A (.DIODE(_06607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14168__A (.DIODE(_06607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14126__A (.DIODE(_06607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14125__A (.DIODE(_06607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15417__A (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15415__A (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15393__A (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14964__A (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14902__B1 (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14900__A (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14458__A (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14165__A (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15526__A (.DIODE(_06649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15509__A (.DIODE(_06649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14394__A (.DIODE(_06649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14247__B1 (.DIODE(_06649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14246__A (.DIODE(_06649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14166__A (.DIODE(_06649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15593__B (.DIODE(_06653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15520__A (.DIODE(_06653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15468__A (.DIODE(_06653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15464__A (.DIODE(_06653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15438__A (.DIODE(_06653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14475__A (.DIODE(_06653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14249__A (.DIODE(_06653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14212__A (.DIODE(_06653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14211__A (.DIODE(_06653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14170__A (.DIODE(_06653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17166__A1 (.DIODE(_06672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15706__B1 (.DIODE(_06672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15580__A1 (.DIODE(_06672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14930__B (.DIODE(_06672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14915__B (.DIODE(_06672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14912__B (.DIODE(_06672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14712__B2 (.DIODE(_06672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14378__A1 (.DIODE(_06672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14316__A2 (.DIODE(_06672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14189__B (.DIODE(_06672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15580__A2 (.DIODE(_06674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14593__A (.DIODE(_06674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14519__A1 (.DIODE(_06674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14192__B (.DIODE(_06674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19542__A1 (.DIODE(_06714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19105__A1 (.DIODE(_06714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14951__B2 (.DIODE(_06714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14431__B2 (.DIODE(_06714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14430__A (.DIODE(_06714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14349__B2 (.DIODE(_06714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14319__B2 (.DIODE(_06714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14318__A (.DIODE(_06714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14242__B2 (.DIODE(_06714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14231__B2 (.DIODE(_06714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19539__A1 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19101__A1 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15206__B2 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15147__A (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14951__A1 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14431__A1 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14349__A1 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14319__A1 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14318__B (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14242__A1 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15788__A (.DIODE(_06736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15738__A (.DIODE(_06736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15718__B (.DIODE(_06736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15184__A (.DIODE(_06736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15125__B (.DIODE(_06736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14545__D (.DIODE(_06736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14257__A (.DIODE(_06736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14253__A (.DIODE(_06736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15780__A1 (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15185__A2 (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15126__B1 (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14816__B (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14672__D (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14608__A2 (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14607__C (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14547__B1 (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14532__B (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14256__C (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15790__A1 (.DIODE(_06738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15227__A (.DIODE(_06738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15185__B1 (.DIODE(_06738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15020__B (.DIODE(_06738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14818__C (.DIODE(_06738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14817__A2 (.DIODE(_06738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14607__D (.DIODE(_06738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14531__A2 (.DIODE(_06738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14258__A (.DIODE(_06738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14255__A (.DIODE(_06738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15228__A2 (.DIODE(_06739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14870__D (.DIODE(_06739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14755__C (.DIODE(_06739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14754__A2 (.DIODE(_06739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14608__B1 (.DIODE(_06739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14552__D (.DIODE(_06739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14551__B1 (.DIODE(_06739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14269__A2 (.DIODE(_06739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14267__C (.DIODE(_06739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14256__D (.DIODE(_06739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14940__B1 (.DIODE(_06741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14939__C (.DIODE(_06741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14870__C (.DIODE(_06741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14869__A2 (.DIODE(_06741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14673__B1 (.DIODE(_06741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14552__C (.DIODE(_06741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14551__A2 (.DIODE(_06741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14279__D (.DIODE(_06741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14270__A (.DIODE(_06741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14259__A2 (.DIODE(_06741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17207__A1 (.DIODE(_06742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15211__B (.DIODE(_06742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15202__A2 (.DIODE(_06742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15128__B (.DIODE(_06742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14935__A2 (.DIODE(_06742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14869__B1 (.DIODE(_06742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14664__B (.DIODE(_06742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14483__B (.DIODE(_06742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14415__B (.DIODE(_06742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14259__B1 (.DIODE(_06742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15778__A (.DIODE(_06744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15718__A (.DIODE(_06744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15682__B (.DIODE(_06744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15125__A (.DIODE(_06744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15117__B (.DIODE(_06744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14545__C (.DIODE(_06744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14263__A (.DIODE(_06744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14261__A (.DIODE(_06744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15080__B (.DIODE(_06745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14940__A2 (.DIODE(_06745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14766__B1 (.DIODE(_06745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14609__B (.DIODE(_06745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14566__B1 (.DIODE(_06745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14565__D (.DIODE(_06745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14300__D (.DIODE(_06745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14280__A2 (.DIODE(_06745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14279__C (.DIODE(_06745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14262__D (.DIODE(_06745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15739__A1 (.DIODE(_06747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15126__A2 (.DIODE(_06747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15118__B1 (.DIODE(_06747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14765__D (.DIODE(_06747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14673__A2 (.DIODE(_06747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14672__C (.DIODE(_06747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14550__B (.DIODE(_06747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14547__A2 (.DIODE(_06747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14421__D (.DIODE(_06747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14264__A (.DIODE(_06747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17199__A1 (.DIODE(_06748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15383__B2 (.DIODE(_06748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15352__A2 (.DIODE(_06748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15173__B (.DIODE(_06748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14941__A1 (.DIODE(_06748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14872__B (.DIODE(_06748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14815__A2 (.DIODE(_06748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14420__B1 (.DIODE(_06748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14301__B1 (.DIODE(_06748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14265__A2_N (.DIODE(_06748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15840__A (.DIODE(_06750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15812__A1 (.DIODE(_06750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15022__C (.DIODE(_06750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15021__A2 (.DIODE(_06750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14817__B1 (.DIODE(_06750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14531__B1 (.DIODE(_06750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14482__C (.DIODE(_06750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14410__A (.DIODE(_06750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14268__A (.DIODE(_06750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14267__D (.DIODE(_06750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17211__A1 (.DIODE(_06752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15246__B (.DIODE(_06752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15237__A2 (.DIODE(_06752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15187__B (.DIODE(_06752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14799__A2 (.DIODE(_06752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14676__A2 (.DIODE(_06752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14661__A2 (.DIODE(_06752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14599__B (.DIODE(_06752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14501__B (.DIODE(_06752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14269__B1 (.DIODE(_06752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17203__A1 (.DIODE(_06754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15163__B (.DIODE(_06754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15144__A2 (.DIODE(_06754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15140__A2 (.DIODE(_06754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15120__B (.DIODE(_06754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14880__A2 (.DIODE(_06754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14757__B (.DIODE(_06754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14409__A2_N (.DIODE(_06754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14280__B1 (.DIODE(_06754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14271__D (.DIODE(_06754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17191__A1 (.DIODE(_06770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15050__B (.DIODE(_06770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15042__B (.DIODE(_06770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14822__B (.DIODE(_06770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14435__A2 (.DIODE(_06770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14424__B (.DIODE(_06770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14303__A2_N (.DIODE(_06770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14302__D (.DIODE(_06770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14288__D (.DIODE(_06770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14287__B1 (.DIODE(_06770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15257__A2 (.DIODE(_06894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15228__B1 (.DIODE(_06894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15074__B (.DIODE(_06894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14863__B (.DIODE(_06894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14755__D (.DIODE(_06894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14754__B1 (.DIODE(_06894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14662__C (.DIODE(_06894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14484__A2 (.DIODE(_06894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14414__A2 (.DIODE(_06894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14413__C (.DIODE(_06894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15877__A (.DIODE(_06895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15811__A (.DIODE(_06895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15789__B (.DIODE(_06895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15280__A (.DIODE(_06895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15256__B (.DIODE(_06895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15022__D (.DIODE(_06895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14481__A (.DIODE(_06895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14412__A (.DIODE(_06895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15257__B1 (.DIODE(_06896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15131__A2 (.DIODE(_06896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15002__B (.DIODE(_06896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14748__B (.DIODE(_06896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14662__D (.DIODE(_06896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14597__A2 (.DIODE(_06896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14499__C (.DIODE(_06896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14484__B1 (.DIODE(_06896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14414__B1 (.DIODE(_06896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14413__D (.DIODE(_06896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15193__A (.DIODE(_06929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14967__B2 (.DIODE(_06929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14966__A (.DIODE(_06929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14686__B2 (.DIODE(_06929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14623__B2 (.DIODE(_06929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14622__A (.DIODE(_06929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14566__B2 (.DIODE(_06929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14551__B2 (.DIODE(_06929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14547__B2 (.DIODE(_06929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14447__A (.DIODE(_06929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14967__A1 (.DIODE(_06930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14966__B (.DIODE(_06930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14686__A1 (.DIODE(_06930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14623__A1 (.DIODE(_06930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14622__B (.DIODE(_06930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14566__A1 (.DIODE(_06930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14552__B (.DIODE(_06930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14551__A1 (.DIODE(_06930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14448__A1 (.DIODE(_06930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14447__B (.DIODE(_06930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15842__A1 (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15112__B (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15076__C (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15075__A2 (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15021__B1 (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14862__A2 (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14861__C (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14523__A (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14500__A2 (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14482__D (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15950__A (.DIODE(_06970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15875__A (.DIODE(_06970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15841__B (.DIODE(_06970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15328__A (.DIODE(_06970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15316__B (.DIODE(_06970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15134__C (.DIODE(_06970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15004__C (.DIODE(_06970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14803__D (.DIODE(_06970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14507__A (.DIODE(_06970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14487__A (.DIODE(_06970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15145__A2_N (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15062__D (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14747__B1 (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14746__D (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14654__A2 (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14653__C (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14592__A2 (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14590__B (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14520__B1 (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14488__A (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17223__A1 (.DIODE(_06972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15341__B (.DIODE(_06972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15327__A2 (.DIODE(_06972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15326__A2 (.DIODE(_06972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15315__B1 (.DIODE(_06972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15308__B (.DIODE(_06972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15307__A2 (.DIODE(_06972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15283__B (.DIODE(_06972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14809__B (.DIODE(_06972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14494__A2 (.DIODE(_06972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15193__C (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15192__A2 (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15133__B1 (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15061__A2 (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15005__B1 (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14653__D (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14589__A2 (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14517__A (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14509__B1 (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14490__A (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15224__C (.DIODE(_06974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15009__A (.DIODE(_06974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14800__C (.DIODE(_06974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14654__B1 (.DIODE(_06974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14588__C (.DIODE(_06974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14534__B2 (.DIODE(_06974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14518__A2 (.DIODE(_06974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14510__A1 (.DIODE(_06974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14493__C (.DIODE(_06974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14492__A2 (.DIODE(_06974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15193__D (.DIODE(_06975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15192__B1 (.DIODE(_06975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15061__B1 (.DIODE(_06975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14589__B1 (.DIODE(_06975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14588__D (.DIODE(_06975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14518__B1 (.DIODE(_06975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14517__B (.DIODE(_06975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14505__A (.DIODE(_06975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14493__D (.DIODE(_06975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14492__B1 (.DIODE(_06975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15114__C (.DIODE(_06982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15075__B1 (.DIODE(_06982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15006__D (.DIODE(_06982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14862__B1 (.DIODE(_06982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14747__A2 (.DIODE(_06982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14597__B1 (.DIODE(_06982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14596__C (.DIODE(_06982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14534__A2 (.DIODE(_06982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14500__B1 (.DIODE(_06982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14499__D (.DIODE(_06982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16120__A (.DIODE(_06989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15329__A2 (.DIODE(_06989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15261__B1 (.DIODE(_06989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15224__D (.DIODE(_06989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15205__A (.DIODE(_06989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15147__D (.DIODE(_06989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15057__B (.DIODE(_06989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15010__B1 (.DIODE(_06989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14800__D (.DIODE(_06989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14506__B (.DIODE(_06989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15918__A1 (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15191__B (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15133__A2 (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15114__D (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15113__B1 (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15005__A2 (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14804__B1 (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14521__D (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14509__A2 (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14508__C (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15919__A (.DIODE(_06995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15876__A1 (.DIODE(_06995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15132__B (.DIODE(_06995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15113__A2 (.DIODE(_06995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15076__D (.DIODE(_06995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14861__D (.DIODE(_06995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14804__A2 (.DIODE(_06995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14521__C (.DIODE(_06995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14520__A2 (.DIODE(_06995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14512__A (.DIODE(_06995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17219__A1 (.DIODE(_06996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15315__A2 (.DIODE(_06996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15293__B (.DIODE(_06996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15291__A2 (.DIODE(_06996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15281__B1 (.DIODE(_06996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15259__B (.DIODE(_06996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15058__A2_N (.DIODE(_06996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14746__C (.DIODE(_06996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14655__B (.DIODE(_06996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14513__B (.DIODE(_06996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14834__A1 (.DIODE(_07000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14813__A (.DIODE(_07000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14544__B1_N (.DIODE(_07000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14542__A_N (.DIODE(_07000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16074__A (.DIODE(_07001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16071__A (.DIODE(_07001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15952__A (.DIODE(_07001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15342__C1 (.DIODE(_07001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14593__B (.DIODE(_07001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14519__A2 (.DIODE(_07001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17215__A1 (.DIODE(_07007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15281__A2 (.DIODE(_07007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15268__B (.DIODE(_07007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15226__B (.DIODE(_07007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14806__A2 (.DIODE(_07007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14750__A2 (.DIODE(_07007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14676__B2 (.DIODE(_07007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14661__B1 (.DIODE(_07007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14598__A1 (.DIODE(_07007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14524__B (.DIODE(_07007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14587__A (.DIODE(_07010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14528__A (.DIODE(_07010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15258__A1 (.DIODE(_07041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15229__A1 (.DIODE(_07041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15186__A1 (.DIODE(_07041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15127__A1 (.DIODE(_07041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15029__A1 (.DIODE(_07041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14840__A (.DIODE(_07041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14825__A1 (.DIODE(_07041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14562__A1 (.DIODE(_07041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15617__B1_N (.DIODE(_07042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15605__A1 (.DIODE(_07042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15604__B (.DIODE(_07042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14841__A2 (.DIODE(_07042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14562__A2 (.DIODE(_07042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19514__A1 (.DIODE(_07043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19066__A (.DIODE(_07043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15327__A1 (.DIODE(_07043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15315__A1 (.DIODE(_07043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15281__A1 (.DIODE(_07043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15257__A1 (.DIODE(_07043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14824__A1 (.DIODE(_07043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14692__A1 (.DIODE(_07043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14629__A1 (.DIODE(_07043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14561__A1 (.DIODE(_07043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19518__A1 (.DIODE(_07044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19078__A1 (.DIODE(_07044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15327__B2 (.DIODE(_07044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15315__B2 (.DIODE(_07044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15281__B2 (.DIODE(_07044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15257__B2 (.DIODE(_07044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14824__B2 (.DIODE(_07044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14692__B2 (.DIODE(_07044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14629__B2 (.DIODE(_07044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14561__B2 (.DIODE(_07044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14708__A1 (.DIODE(_07088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14706__B1 (.DIODE(_07088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14684__A1 (.DIODE(_07088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14652__A (.DIODE(_07088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14619__A1 (.DIODE(_07088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14618__A (.DIODE(_07088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14652__B (.DIODE(_07089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14619__A2 (.DIODE(_07089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14618__B (.DIODE(_07089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15352__A1 (.DIODE(_07200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15326__A1 (.DIODE(_07200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15323__A1 (.DIODE(_07200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15291__A1 (.DIODE(_07200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15237__A1 (.DIODE(_07200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15104__A (.DIODE(_07200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14915__A (.DIODE(_07200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14788__A (.DIODE(_07200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14722__A (.DIODE(_07200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14717__A (.DIODE(_07200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19524__A1 (.DIODE(_07206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19086__A1 (.DIODE(_07206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15202__A1 (.DIODE(_07206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15144__A1 (.DIODE(_07206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15050__A (.DIODE(_07206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14930__A (.DIODE(_07206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14923__A (.DIODE(_07206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14851__A1 (.DIODE(_07206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14726__A (.DIODE(_07206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14723__A (.DIODE(_07206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15001__B1 (.DIODE(_07295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15000__C (.DIODE(_07295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14812__C (.DIODE(_07295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15637__A1 (.DIODE(_07307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15609__B (.DIODE(_07307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15040__A2 (.DIODE(_07307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14825__A2 (.DIODE(_07307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15343__A (.DIODE(_07324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15306__A (.DIODE(_07324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15288__A1 (.DIODE(_07324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15282__A1 (.DIODE(_07324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15266__B2 (.DIODE(_07324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15234__A1 (.DIODE(_07324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15199__A1 (.DIODE(_07324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15094__A1 (.DIODE(_07324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15040__A1 (.DIODE(_07324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14841__A1 (.DIODE(_07324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17227__A1 (.DIODE(_07493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15333__B (.DIODE(_07493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15327__B1 (.DIODE(_07493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15323__A2 (.DIODE(_07493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15318__B (.DIODE(_07493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15317__A2 (.DIODE(_07493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15261__A2 (.DIODE(_07493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15206__A2 (.DIODE(_07493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15147__C (.DIODE(_07493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15010__A2 (.DIODE(_07493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15056__B (.DIODE(_07495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15012__B (.DIODE(_07495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15641__B1_N (.DIODE(_07511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15094__A2 (.DIODE(_07511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15029__A2 (.DIODE(_07511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15334__A1 (.DIODE(_07565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15329__B2 (.DIODE(_07565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15317__B2 (.DIODE(_07565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15171__A1_N (.DIODE(_07565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15140__B2 (.DIODE(_07565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15119__A1 (.DIODE(_07565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15084__A1 (.DIODE(_07565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15659__B1 (.DIODE(_07566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15171__A2_N (.DIODE(_07566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15084__A2 (.DIODE(_07566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15103__B1 (.DIODE(_07578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15095__B (.DIODE(_07578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15683__B1 (.DIODE(_07601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15140__B1 (.DIODE(_07601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15119__A2 (.DIODE(_07601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15719__B1_N (.DIODE(_07609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15199__A2 (.DIODE(_07609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15127__A2 (.DIODE(_07609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16193__A (.DIODE(_07668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16191__A (.DIODE(_07668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15739__B1_N (.DIODE(_07668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15234__A2 (.DIODE(_07668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15186__A2 (.DIODE(_07668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17229__A0 (.DIODE(_07689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16178__A (.DIODE(_07689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16171__A1 (.DIODE(_07689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16137__A (.DIODE(_07689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15331__A2 (.DIODE(_07689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15330__B (.DIODE(_07689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15320__A2 (.DIODE(_07689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15285__B (.DIODE(_07689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15242__B (.DIODE(_07689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15206__B1 (.DIODE(_07689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15780__B1_N (.DIODE(_07711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15266__B1 (.DIODE(_07711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15229__A2 (.DIODE(_07711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15790__B1_N (.DIODE(_07740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15288__A2 (.DIODE(_07740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15258__A2 (.DIODE(_07740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15812__B1_N (.DIODE(_07764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15306__B (.DIODE(_07764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15282__A2 (.DIODE(_07764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15842__B1 (.DIODE(_07800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15334__A2 (.DIODE(_07800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15317__B1 (.DIODE(_07800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15331__B1 (.DIODE(_07813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15330__C (.DIODE(_07813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16357__A (.DIODE(_07934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16345__A1 (.DIODE(_07934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15486__A1 (.DIODE(_07934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15490__B (.DIODE(_07958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15489__A2 (.DIODE(_07958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15480__A1 (.DIODE(_07958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15476__B1 (.DIODE(_07958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16340__A (.DIODE(_07970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16339__A (.DIODE(_07970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16332__A1 (.DIODE(_07970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15492__B (.DIODE(_07970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16264__A0 (.DIODE(_08066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16262__A (.DIODE(_08066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16257__A0 (.DIODE(_08066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16248__A (.DIODE(_08066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16245__A (.DIODE(_08066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15772__A (.DIODE(_08066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15771__A (.DIODE(_08066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15704__A1 (.DIODE(_08066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15602__A (.DIODE(_08066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15583__C1 (.DIODE(_08066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15600__A2 (.DIODE(_08080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15599__A2 (.DIODE(_08080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19123__A1 (.DIODE(_08081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16414__B1 (.DIODE(_08081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16387__S (.DIODE(_08081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16370__B1 (.DIODE(_08081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16358__A (.DIODE(_08081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16352__B1 (.DIODE(_08081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16341__A (.DIODE(_08081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16324__A (.DIODE(_08081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16288__A (.DIODE(_08081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15598__A (.DIODE(_08081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19561__A1 (.DIODE(_08082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16426__A1 (.DIODE(_08082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16402__A1 (.DIODE(_08082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16393__A1_N (.DIODE(_08082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16368__A1 (.DIODE(_08082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16354__A1 (.DIODE(_08082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16322__A (.DIODE(_08082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16317__A1 (.DIODE(_08082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16289__A1 (.DIODE(_08082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15599__B1 (.DIODE(_08082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15601__B2 (.DIODE(_08084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17155__A0 (.DIODE(_08085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16282__A1 (.DIODE(_08085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16281__A (.DIODE(_08085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16280__A0 (.DIODE(_08085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15765__A (.DIODE(_08085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15712__A0 (.DIODE(_08085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15702__A1 (.DIODE(_08085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15701__A0 (.DIODE(_08085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15681__A (.DIODE(_08085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15680__A (.DIODE(_08085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15803__A (.DIODE(_08090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15796__A (.DIODE(_08090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15724__A (.DIODE(_08090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15687__A (.DIODE(_08090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15612__A (.DIODE(_08090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15611__A (.DIODE(_08090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16111__A (.DIODE(_08093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16089__A (.DIODE(_08093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15804__A1 (.DIODE(_08093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15797__A (.DIODE(_08093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15727__A_N (.DIODE(_08093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15726__B (.DIODE(_08093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15612__B (.DIODE(_08093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15611__B (.DIODE(_08093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15689__A (.DIODE(_08099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15663__A1 (.DIODE(_08099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15622__A (.DIODE(_08099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15619__A (.DIODE(_08099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15618__A (.DIODE(_08099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15825__A (.DIODE(_08122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15817__A (.DIODE(_08122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15743__A (.DIODE(_08122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15722__A (.DIODE(_08122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15643__A (.DIODE(_08122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15642__A (.DIODE(_08122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16114__A (.DIODE(_08124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16110__A (.DIODE(_08124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15826__A (.DIODE(_08124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15818__A (.DIODE(_08124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15751__A2 (.DIODE(_08124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15745__B (.DIODE(_08124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15643__B (.DIODE(_08124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15642__B (.DIODE(_08124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15939__A1 (.DIODE(_08127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15934__A (.DIODE(_08127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15649__A2 (.DIODE(_08127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15645__B (.DIODE(_08127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15856__A1 (.DIODE(_08142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15847__A (.DIODE(_08142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15786__B (.DIODE(_08142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15662__A (.DIODE(_08142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15661__A (.DIODE(_08142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15849__A (.DIODE(_08143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15848__A (.DIODE(_08143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15784__A (.DIODE(_08143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15742__A1 (.DIODE(_08143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15662__B (.DIODE(_08143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15661__B (.DIODE(_08143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16151__A (.DIODE(_08166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15890__A1 (.DIODE(_08166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15882__A (.DIODE(_08166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15803__B (.DIODE(_08166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15796__B (.DIODE(_08166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15686__A (.DIODE(_08166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15685__A (.DIODE(_08166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15884__A (.DIODE(_08167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15883__A (.DIODE(_08167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15794__A (.DIODE(_08167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15783__A1 (.DIODE(_08167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15686__B (.DIODE(_08167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15685__B (.DIODE(_08167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15926__A (.DIODE(_08200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15925__A (.DIODE(_08200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15809__A (.DIODE(_08200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15793__A1 (.DIODE(_08200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15721__A (.DIODE(_08200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15720__A (.DIODE(_08200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16159__A (.DIODE(_08202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15932__A1 (.DIODE(_08202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15924__A (.DIODE(_08202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15825__B (.DIODE(_08202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15817__B (.DIODE(_08202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15721__B (.DIODE(_08202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15720__B (.DIODE(_08202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15956__A (.DIODE(_08220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15955__A (.DIODE(_08220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15839__A (.DIODE(_08220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15815__A1 (.DIODE(_08220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15741__A (.DIODE(_08220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15740__A (.DIODE(_08220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16168__A (.DIODE(_08222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16166__A1 (.DIODE(_08222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15962__A1 (.DIODE(_08222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15958__A (.DIODE(_08222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15849__B (.DIODE(_08222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15848__B (.DIODE(_08222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15741__B (.DIODE(_08222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15740__B (.DIODE(_08222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15991__A (.DIODE(_08261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15985__A (.DIODE(_08261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15873__A (.DIODE(_08261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15845__A1 (.DIODE(_08261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15782__A (.DIODE(_08261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15781__A (.DIODE(_08261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16177__A (.DIODE(_08263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16174__A (.DIODE(_08263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15987__A (.DIODE(_08263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15986__A (.DIODE(_08263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15884__B (.DIODE(_08263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15883__B (.DIODE(_08263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15782__B (.DIODE(_08263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15781__B (.DIODE(_08263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16021__A (.DIODE(_08271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16016__A (.DIODE(_08271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15914__A (.DIODE(_08271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15874__A (.DIODE(_08271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15792__A (.DIODE(_08271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15791__A (.DIODE(_08271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16192__A (.DIODE(_08273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16185__A (.DIODE(_08273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16183__A1 (.DIODE(_08273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16022__A (.DIODE(_08273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16017__A (.DIODE(_08273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15926__B (.DIODE(_08273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15925__B (.DIODE(_08273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15792__B (.DIODE(_08273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15791__B (.DIODE(_08273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16123__A (.DIODE(_08298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16118__A1 (.DIODE(_08298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15819__A_N (.DIODE(_08298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15816__B (.DIODE(_08298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16075__A1 (.DIODE(_08325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16072__A (.DIODE(_08325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15991__B (.DIODE(_08325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15985__B (.DIODE(_08325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15872__B (.DIODE(_08325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15844__B (.DIODE(_08325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15843__B (.DIODE(_08325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16223__A2 (.DIODE(_08330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16132__A (.DIODE(_08330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16131__A1 (.DIODE(_08330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15851__A (.DIODE(_08330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16160__A (.DIODE(_08364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16153__A1 (.DIODE(_08364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15913__A (.DIODE(_08364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15888__A1 (.DIODE(_08364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16170__A (.DIODE(_08399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16161__A1 (.DIODE(_08399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16121__B (.DIODE(_08399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16100__B (.DIODE(_08399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16014__B (.DIODE(_08399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15982__B (.DIODE(_08399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15950__B (.DIODE(_08399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15918__A2 (.DIODE(_08399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16117__B (.DIODE(_08404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16116__B (.DIODE(_08404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15922__B1 (.DIODE(_08404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16211__A2 (.DIODE(_08425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15943__B (.DIODE(_08425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15978__B (.DIODE(_08443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15965__B (.DIODE(_08443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15961__B (.DIODE(_08443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15968__A_N (.DIODE(_08445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15963__B (.DIODE(_08445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16425__A1 (.DIODE(_08683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16424__A (.DIODE(_08683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16202__A2 (.DIODE(_08683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16370__A4 (.DIODE(_08695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16213__B1 (.DIODE(_08695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16372__A2_N (.DIODE(_08696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16366__C (.DIODE(_08696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16365__A2 (.DIODE(_08696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16214__B (.DIODE(_08696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16291__A1 (.DIODE(_08772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17235__A (.DIODE(_08773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16388__S (.DIODE(_08773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16373__S (.DIODE(_08773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16360__S (.DIODE(_08773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16343__S (.DIODE(_08773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16336__S (.DIODE(_08773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16318__S (.DIODE(_08773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16308__S (.DIODE(_08773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16300__S (.DIODE(_08773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16291__S (.DIODE(_08773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16300__A1 (.DIODE(_08781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16308__A1 (.DIODE(_08788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16318__A1 (.DIODE(_08797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16326__B1_N (.DIODE(_08804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16335__A1_N (.DIODE(_08808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16335__A2_N (.DIODE(_08809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16336__A1 (.DIODE(_08813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16342__B1 (.DIODE(_08818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16343__A1 (.DIODE(_08819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16354__B1 (.DIODE(_08829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16355__B1_N (.DIODE(_08830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16359__B1 (.DIODE(_08833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16360__A1 (.DIODE(_08834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16368__B1 (.DIODE(_08841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16372__B2 (.DIODE(_08844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16373__A1 (.DIODE(_08845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16407__B2 (.DIODE(_08853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16382__B_N (.DIODE(_08853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16387__A1 (.DIODE(_08858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16393__B1 (.DIODE(_08862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16393__B2 (.DIODE(_08863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16402__A2 (.DIODE(_08867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16402__A3 (.DIODE(_08868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16407__B1 (.DIODE(_08875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16415__A2 (.DIODE(_08880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16416__A1 (.DIODE(_08883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16426__A2 (.DIODE(_08888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16427__B1_N (.DIODE(_08893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16853__A (.DIODE(_08895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16641__A2 (.DIODE(_08895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16631__A2 (.DIODE(_08895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16609__A2 (.DIODE(_08895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16598__A (.DIODE(_08895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16596__A (.DIODE(_08895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16462__B (.DIODE(_08895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16460__A1 (.DIODE(_08895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16458__A (.DIODE(_08895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16430__A (.DIODE(_08895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17024__B2 (.DIODE(_08896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16831__A2 (.DIODE(_08896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16828__A2 (.DIODE(_08896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16825__A2 (.DIODE(_08896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16819__A2 (.DIODE(_08896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16817__A2 (.DIODE(_08896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16813__B2 (.DIODE(_08896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16590__A2 (.DIODE(_08896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16453__B2 (.DIODE(_08896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16449__A1 (.DIODE(_08896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16882__S (.DIODE(_08902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16880__S (.DIODE(_08902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16879__S (.DIODE(_08902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16687__S (.DIODE(_08902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16685__S (.DIODE(_08902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16676__B (.DIODE(_08902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16665__S (.DIODE(_08902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16490__A (.DIODE(_08902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16445__A (.DIODE(_08902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16437__B (.DIODE(_08902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16900__A1 (.DIODE(_08904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16899__B_N (.DIODE(_08904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16693__B_N (.DIODE(_08904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16684__S (.DIODE(_08904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16674__S (.DIODE(_08904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16648__B_N (.DIODE(_08904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16500__B (.DIODE(_08904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16452__A (.DIODE(_08904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16442__A (.DIODE(_08904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16439__B (.DIODE(_08904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17238__C1 (.DIODE(_08907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16449__A2 (.DIODE(_08907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16910__A1 (.DIODE(_08908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16905__S (.DIODE(_08908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16859__B_N (.DIODE(_08908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16704__A1 (.DIODE(_08908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16700__S (.DIODE(_08908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16694__A1 (.DIODE(_08908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16659__A1 (.DIODE(_08908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16529__B (.DIODE(_08908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16524__A1 (.DIODE(_08908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16443__A (.DIODE(_08908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16917__A1 (.DIODE(_08909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16913__A1 (.DIODE(_08909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16860__A1 (.DIODE(_08909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16655__A1 (.DIODE(_08909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16649__A1 (.DIODE(_08909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16538__A1 (.DIODE(_08909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16533__B (.DIODE(_08909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16504__A2 (.DIODE(_08909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16453__B1 (.DIODE(_08909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16448__A1 (.DIODE(_08909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16906__A (.DIODE(_08910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16866__S (.DIODE(_08910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16701__A (.DIODE(_08910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16696__A (.DIODE(_08910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16692__S (.DIODE(_08910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16663__S (.DIODE(_08910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16503__A (.DIODE(_08910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16501__A (.DIODE(_08910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16459__B2 (.DIODE(_08910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16448__A2 (.DIODE(_08910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16923__A1 (.DIODE(_08912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16921__A1 (.DIODE(_08912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16914__A (.DIODE(_08912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16908__A1 (.DIODE(_08912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16714__A1 (.DIODE(_08912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16709__A1 (.DIODE(_08912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16703__A1 (.DIODE(_08912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16690__A1 (.DIODE(_08912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16526__A1 (.DIODE(_08912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16447__A (.DIODE(_08912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16931__A1 (.DIODE(_08913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16928__A1 (.DIODE(_08913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16926__A1 (.DIODE(_08913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16863__A1 (.DIODE(_08913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16719__A1 (.DIODE(_08913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16718__A1 (.DIODE(_08913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16715__A1 (.DIODE(_08913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16656__A1 (.DIODE(_08913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16652__A1 (.DIODE(_08913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16448__B1 (.DIODE(_08913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17023__B1 (.DIODE(_08915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16823__A (.DIODE(_08915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16812__B1 (.DIODE(_08915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16639__A (.DIODE(_08915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16630__A (.DIODE(_08915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16623__A (.DIODE(_08915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16620__A (.DIODE(_08915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16617__A (.DIODE(_08915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16608__A (.DIODE(_08915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16451__A (.DIODE(_08915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17239__A1 (.DIODE(_08916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17062__B1 (.DIODE(_08916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17057__B1 (.DIODE(_08916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17054__B1 (.DIODE(_08916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17051__B1 (.DIODE(_08916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17046__B1 (.DIODE(_08916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17043__B1 (.DIODE(_08916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17037__B1 (.DIODE(_08916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17034__B1 (.DIODE(_08916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16453__A1_N (.DIODE(_08916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16637__C (.DIODE(_08918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16634__A (.DIODE(_08918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16615__A (.DIODE(_08918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16612__B (.DIODE(_08918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16605__A (.DIODE(_08918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16591__A (.DIODE(_08918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16455__A (.DIODE(_08918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17064__A1 (.DIODE(_08919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17059__A1 (.DIODE(_08919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17048__A1 (.DIODE(_08919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17032__A1 (.DIODE(_08919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16852__A1 (.DIODE(_08919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16644__B1 (.DIODE(_08919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16602__C1 (.DIODE(_08919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16589__C1 (.DIODE(_08919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16460__A0 (.DIODE(_08919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16459__A2 (.DIODE(_08919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16891__A2 (.DIODE(_08921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16883__A2 (.DIODE(_08921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16688__A2 (.DIODE(_08921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16529__C (.DIODE(_08921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16478__A (.DIODE(_08921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16459__A3 (.DIODE(_08921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17067__A2 (.DIODE(_08922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17040__A2 (.DIODE(_08922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17030__A2 (.DIODE(_08922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17027__A2 (.DIODE(_08922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16848__A2 (.DIODE(_08922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16844__A2 (.DIODE(_08922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16841__A2 (.DIODE(_08922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16834__A2 (.DIODE(_08922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16594__B1 (.DIODE(_08922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16459__B1 (.DIODE(_08922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16960__A (.DIODE(_08927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16760__A (.DIODE(_08927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16756__B1 (.DIODE(_08927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16753__B1 (.DIODE(_08927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16750__A (.DIODE(_08927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16536__A (.DIODE(_08927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16535__A (.DIODE(_08927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16527__B1 (.DIODE(_08927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16483__A (.DIODE(_08927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16468__A (.DIODE(_08927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16957__B1 (.DIODE(_08928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16954__A (.DIODE(_08928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16951__A (.DIODE(_08928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16747__B1 (.DIODE(_08928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16744__A (.DIODE(_08928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16741__B1 (.DIODE(_08928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16531__A0 (.DIODE(_08928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16518__A1 (.DIODE(_08928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16513__A0 (.DIODE(_08928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16469__A (.DIODE(_08928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16948__B1 (.DIODE(_08929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16946__A (.DIODE(_08929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16738__B1 (.DIODE(_08929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16735__A (.DIODE(_08929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16733__B1 (.DIODE(_08929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16505__B2 (.DIODE(_08929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16497__A0 (.DIODE(_08929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16492__A (.DIODE(_08929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16491__A (.DIODE(_08929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16470__A (.DIODE(_08929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16935__A (.DIODE(_08930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16932__B1 (.DIODE(_08930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16809__A1 (.DIODE(_08930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16722__A1 (.DIODE(_08930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16721__A1 (.DIODE(_08930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16720__B1 (.DIODE(_08930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16590__A1 (.DIODE(_08930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16589__A1 (.DIODE(_08930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16482__A (.DIODE(_08930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16471__A (.DIODE(_08930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16918__B2 (.DIODE(_08937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16915__B2 (.DIODE(_08937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16911__A (.DIODE(_08937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16870__A (.DIODE(_08937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16711__B2 (.DIODE(_08937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16667__A (.DIODE(_08937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16511__A (.DIODE(_08937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16496__B (.DIODE(_08937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16481__A (.DIODE(_08937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16478__B (.DIODE(_08937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16891__B1 (.DIODE(_08940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16883__B1 (.DIODE(_08940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16688__B1 (.DIODE(_08940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16677__A2 (.DIODE(_08940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16533__C (.DIODE(_08940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16508__A1 (.DIODE(_08940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16481__B (.DIODE(_08940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16907__A1 (.DIODE(_08944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16903__A1 (.DIODE(_08944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16702__A1 (.DIODE(_08944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16697__A1 (.DIODE(_08944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16485__B (.DIODE(_08944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16906__B (.DIODE(_08948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16902__B (.DIODE(_08948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16894__A1 (.DIODE(_08948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16883__C1 (.DIODE(_08948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16701__B (.DIODE(_08948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16696__B (.DIODE(_08948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16688__C1 (.DIODE(_08948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16681__A1 (.DIODE(_08948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16489__B (.DIODE(_08948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16912__B2 (.DIODE(_08959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16904__A1 (.DIODE(_08959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16706__B2 (.DIODE(_08959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16698__A1 (.DIODE(_08959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16668__A1 (.DIODE(_08959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16533__A (.DIODE(_08959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16529__A (.DIODE(_08959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16515__A (.DIODE(_08959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16502__A (.DIODE(_08959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16500__A (.DIODE(_08959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16929__A1 (.DIODE(_08962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16924__A1 (.DIODE(_08962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16919__A1 (.DIODE(_08962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16871__A1 (.DIODE(_08962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16861__A (.DIODE(_08962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16716__A1 (.DIODE(_08962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16712__A1 (.DIODE(_08962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16660__A1 (.DIODE(_08962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16650__A (.DIODE(_08962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16504__A1 (.DIODE(_08962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16918__A1 (.DIODE(_08967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16915__A1 (.DIODE(_08967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16912__A1 (.DIODE(_08967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16871__B2 (.DIODE(_08967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16711__A1 (.DIODE(_08967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16668__B2 (.DIODE(_08967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16534__A2 (.DIODE(_08967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16530__A3 (.DIODE(_08967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16512__A2 (.DIODE(_08967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16508__A2 (.DIODE(_08967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16907__B2 (.DIODE(_08976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16903__B2 (.DIODE(_08976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16894__B2 (.DIODE(_08976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16885__B2 (.DIODE(_08976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16702__B2 (.DIODE(_08976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16697__B2 (.DIODE(_08976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16690__B2 (.DIODE(_08976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16681__B2 (.DIODE(_08976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16517__A2 (.DIODE(_08976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16869__S (.DIODE(_08982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16858__S (.DIODE(_08982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16695__S (.DIODE(_08982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16689__A1 (.DIODE(_08982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16666__S (.DIODE(_08982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16647__S (.DIODE(_08982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16538__A2 (.DIODE(_08982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16530__A1 (.DIODE(_08982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16526__A2 (.DIODE(_08982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16523__A (.DIODE(_08982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17020__A1 (.DIODE(_09004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16966__A (.DIODE(_09004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16963__B1 (.DIODE(_09004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16941__A (.DIODE(_09004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16938__B1 (.DIODE(_09004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16545__A (.DIODE(_09004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17040__B1 (.DIODE(_09050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17030__B1 (.DIODE(_09050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16838__A1 (.DIODE(_09050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16836__A1 (.DIODE(_09050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16821__A1 (.DIODE(_09050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16819__B1 (.DIODE(_09050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16817__B1 (.DIODE(_09050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16815__A1 (.DIODE(_09050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16597__A1 (.DIODE(_09050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16594__A1 (.DIODE(_09050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17064__B1 (.DIODE(_09054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17059__B1 (.DIODE(_09054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17048__B1 (.DIODE(_09054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17032__B1 (.DIODE(_09054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16852__B1 (.DIODE(_09054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16838__B1 (.DIODE(_09054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16836__B1 (.DIODE(_09054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16821__B1 (.DIODE(_09054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16815__B1 (.DIODE(_09054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16597__B1 (.DIODE(_09054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16638__A2 (.DIODE(_09055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16635__A2 (.DIODE(_09055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16628__A2 (.DIODE(_09055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16625__A2 (.DIODE(_09055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16622__A2 (.DIODE(_09055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16619__A2 (.DIODE(_09055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16616__A2 (.DIODE(_09055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16613__A2 (.DIODE(_09055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16606__A2 (.DIODE(_09055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16603__A2 (.DIODE(_09055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17238__A2 (.DIODE(_09056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16854__B1 (.DIODE(_09056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16641__B1 (.DIODE(_09056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16631__B1 (.DIODE(_09056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16609__B1 (.DIODE(_09056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16600__A (.DIODE(_09056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16638__B1 (.DIODE(_09057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16635__B1 (.DIODE(_09057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16628__B1 (.DIODE(_09057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16625__B1 (.DIODE(_09057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16622__B1 (.DIODE(_09057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16619__B1 (.DIODE(_09057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16616__B1 (.DIODE(_09057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16613__B1 (.DIODE(_09057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16606__B1 (.DIODE(_09057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16603__B1 (.DIODE(_09057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17062__A2 (.DIODE(_09086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17057__A2 (.DIODE(_09086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17054__A2 (.DIODE(_09086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17051__A2 (.DIODE(_09086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17046__A2 (.DIODE(_09086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17043__A2 (.DIODE(_09086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17037__A2 (.DIODE(_09086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17034__A2 (.DIODE(_09086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16850__B1 (.DIODE(_09086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16645__A2 (.DIODE(_09086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17066__A (.DIODE(_09261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17026__B1 (.DIODE(_09261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16850__A1 (.DIODE(_09261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16847__A (.DIODE(_09261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16843__A (.DIODE(_09261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16840__A (.DIODE(_09261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16833__A (.DIODE(_09261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16830__A (.DIODE(_09261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16827__A (.DIODE(_09261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16824__A (.DIODE(_09261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17161__A2 (.DIODE(_09282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17027__A1 (.DIODE(_09282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17017__A (.DIODE(_09282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16934__A (.DIODE(_09282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17155__A1 (.DIODE(_09544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17229__S (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17226__C1 (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17222__C1 (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17218__C1 (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17214__C1 (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17210__C1 (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17164__A (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17155__S (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17239__A2 (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17227__A2 (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17223__A2 (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17219__A2 (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17215__A2 (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17211__A2 (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17159__A (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17166__B1 (.DIODE(_09555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17173__B1 (.DIODE(_09560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17173__B2 (.DIODE(_09561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17179__B1 (.DIODE(_09563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17179__B2 (.DIODE(_09566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17183__B1 (.DIODE(_09568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17183__B2 (.DIODE(_09569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17187__B1 (.DIODE(_09571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17187__B2 (.DIODE(_09572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17191__B1 (.DIODE(_09574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17191__B2 (.DIODE(_09575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17195__B1 (.DIODE(_09577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17195__B2 (.DIODE(_09578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17199__B1 (.DIODE(_09580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17199__B2 (.DIODE(_09581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17203__B1 (.DIODE(_09583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17203__B2 (.DIODE(_09584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17207__B1 (.DIODE(_09586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17207__B2 (.DIODE(_09587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17211__B1 (.DIODE(_09589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17211__B2 (.DIODE(_09590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17215__B1 (.DIODE(_09592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17215__B2 (.DIODE(_09593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17223__B1 (.DIODE(_09598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17223__B2 (.DIODE(_09599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17229__A1 (.DIODE(_09603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17238__B1 (.DIODE(_09605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17235__B (.DIODE(_09605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17356__S (.DIODE(_09607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17352__S (.DIODE(_09607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17348__S (.DIODE(_09607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17344__S (.DIODE(_09607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17340__S (.DIODE(_09607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17336__S (.DIODE(_09607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17332__S (.DIODE(_09607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17328__S (.DIODE(_09607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17324__S (.DIODE(_09607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17234__A (.DIODE(_09607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17320__S (.DIODE(_09608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17316__S (.DIODE(_09608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17312__S (.DIODE(_09608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17308__S (.DIODE(_09608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17304__S (.DIODE(_09608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17300__S (.DIODE(_09608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17296__S (.DIODE(_09608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17292__S (.DIODE(_09608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17288__S (.DIODE(_09608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17235__C_N (.DIODE(_09608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18157__A2 (.DIODE(_09754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17439__B1 (.DIODE(_09754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17437__B1 (.DIODE(_09754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17433__B1 (.DIODE(_09754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17430__B1 (.DIODE(_09754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17427__A1 (.DIODE(_09754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17424__B1 (.DIODE(_09754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17421__B1 (.DIODE(_09754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17418__B1 (.DIODE(_09754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17413__A0 (.DIODE(_09754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17439__A2 (.DIODE(_09756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17437__A2 (.DIODE(_09756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17433__A2 (.DIODE(_09756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17430__A2 (.DIODE(_09756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17427__B1 (.DIODE(_09756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17424__A2 (.DIODE(_09756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17421__A2 (.DIODE(_09756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17418__A2 (.DIODE(_09756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17413__A1 (.DIODE(_09756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18757__A1 (.DIODE(_09782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18577__A1 (.DIODE(_09782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17729__S (.DIODE(_09782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17463__S (.DIODE(_09782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17460__A1 (.DIODE(_09782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17459__B_N (.DIODE(_09782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17457__S (.DIODE(_09782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17453__A1 (.DIODE(_09782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17452__B_N (.DIODE(_09782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17449__A1 (.DIODE(_09782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17717__C1 (.DIODE(_09791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17710__C1 (.DIODE(_09791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17638__A (.DIODE(_09791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17563__A (.DIODE(_09791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17473__A (.DIODE(_09791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17467__A (.DIODE(_09791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17717__B1 (.DIODE(_09801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17710__B1 (.DIODE(_09801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17637__A (.DIODE(_09801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17562__A (.DIODE(_09801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17472__A (.DIODE(_09801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17467__B (.DIODE(_09801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17719__B (.DIODE(_09803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17712__B (.DIODE(_09803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17705__B (.DIODE(_09803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17698__B (.DIODE(_09803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17691__B (.DIODE(_09803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17684__B (.DIODE(_09803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17677__B (.DIODE(_09803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17527__A (.DIODE(_09803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17490__B1 (.DIODE(_09803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17469__A (.DIODE(_09803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17718__A2 (.DIODE(_09804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17711__A2 (.DIODE(_09804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17635__A (.DIODE(_09804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17560__A (.DIODE(_09804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17520__B (.DIODE(_09804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17513__B (.DIODE(_09804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17506__B (.DIODE(_09804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17499__B (.DIODE(_09804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17492__B (.DIODE(_09804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17470__A (.DIODE(_09804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17555__A2 (.DIODE(_09805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17548__A2 (.DIODE(_09805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17541__A2 (.DIODE(_09805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17534__A2 (.DIODE(_09805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17526__A2 (.DIODE(_09805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17519__A2 (.DIODE(_09805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17512__A2 (.DIODE(_09805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17505__A2 (.DIODE(_09805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17498__A2 (.DIODE(_09805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17475__A2 (.DIODE(_09805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17554__B1 (.DIODE(_09807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17547__B1 (.DIODE(_09807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17540__B1 (.DIODE(_09807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17533__B1 (.DIODE(_09807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17525__B1 (.DIODE(_09807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17518__B1 (.DIODE(_09807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17511__B1 (.DIODE(_09807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17504__B1 (.DIODE(_09807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17497__B1 (.DIODE(_09807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17474__B1 (.DIODE(_09807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17554__C1 (.DIODE(_09808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17547__C1 (.DIODE(_09808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17540__C1 (.DIODE(_09808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17533__C1 (.DIODE(_09808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17525__C1 (.DIODE(_09808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17518__C1 (.DIODE(_09808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17511__C1 (.DIODE(_09808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17504__C1 (.DIODE(_09808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17497__C1 (.DIODE(_09808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17474__C1 (.DIODE(_09808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17720__A1 (.DIODE(_09825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17713__A1 (.DIODE(_09825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17641__A (.DIODE(_09825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17566__A (.DIODE(_09825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17491__A (.DIODE(_09825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17557__A1 (.DIODE(_09826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17550__A1 (.DIODE(_09826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17543__A1 (.DIODE(_09826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17536__A1 (.DIODE(_09826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17529__A1 (.DIODE(_09826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17521__A1 (.DIODE(_09826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17514__A1 (.DIODE(_09826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17507__A1 (.DIODE(_09826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17500__A1 (.DIODE(_09826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17493__A1 (.DIODE(_09826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17595__B (.DIODE(_09857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17588__B (.DIODE(_09857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17581__B (.DIODE(_09857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17574__B (.DIODE(_09857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17567__B (.DIODE(_09857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17556__B (.DIODE(_09857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17549__B (.DIODE(_09857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17542__B (.DIODE(_09857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17535__B (.DIODE(_09857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17528__B (.DIODE(_09857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17630__A2 (.DIODE(_09885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17623__A2 (.DIODE(_09885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17616__A2 (.DIODE(_09885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17609__A2 (.DIODE(_09885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17601__A2 (.DIODE(_09885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17594__A2 (.DIODE(_09885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17587__A2 (.DIODE(_09885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17580__A2 (.DIODE(_09885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17573__A2 (.DIODE(_09885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17565__A2 (.DIODE(_09885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17629__B1 (.DIODE(_09887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17622__B1 (.DIODE(_09887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17615__B1 (.DIODE(_09887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17608__B1 (.DIODE(_09887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17600__B1 (.DIODE(_09887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17593__B1 (.DIODE(_09887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17586__B1 (.DIODE(_09887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17579__B1 (.DIODE(_09887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17572__B1 (.DIODE(_09887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17564__B1 (.DIODE(_09887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17629__C1 (.DIODE(_09888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17622__C1 (.DIODE(_09888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17615__C1 (.DIODE(_09888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17608__C1 (.DIODE(_09888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17600__C1 (.DIODE(_09888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17593__C1 (.DIODE(_09888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17586__C1 (.DIODE(_09888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17579__C1 (.DIODE(_09888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17572__C1 (.DIODE(_09888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17564__C1 (.DIODE(_09888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17632__A1 (.DIODE(_09891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17625__A1 (.DIODE(_09891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17618__A1 (.DIODE(_09891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17611__A1 (.DIODE(_09891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17604__A1 (.DIODE(_09891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17596__A1 (.DIODE(_09891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17589__A1 (.DIODE(_09891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17582__A1 (.DIODE(_09891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17575__A1 (.DIODE(_09891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17568__A1 (.DIODE(_09891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17670__B (.DIODE(_09922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17663__B (.DIODE(_09922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17656__B (.DIODE(_09922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17649__B (.DIODE(_09922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17642__B (.DIODE(_09922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17631__B (.DIODE(_09922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17624__B (.DIODE(_09922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17617__B (.DIODE(_09922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17610__B (.DIODE(_09922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17603__B (.DIODE(_09922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17704__A2 (.DIODE(_09950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17697__A2 (.DIODE(_09950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17690__A2 (.DIODE(_09950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17683__A2 (.DIODE(_09950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17676__A2 (.DIODE(_09950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17669__A2 (.DIODE(_09950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17662__A2 (.DIODE(_09950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17655__A2 (.DIODE(_09950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17648__A2 (.DIODE(_09950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17640__A2 (.DIODE(_09950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17703__B1 (.DIODE(_09952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17696__B1 (.DIODE(_09952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17689__B1 (.DIODE(_09952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17682__B1 (.DIODE(_09952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17675__B1 (.DIODE(_09952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17668__B1 (.DIODE(_09952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17661__B1 (.DIODE(_09952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17654__B1 (.DIODE(_09952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17647__B1 (.DIODE(_09952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17639__B1 (.DIODE(_09952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17703__C1 (.DIODE(_09953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17696__C1 (.DIODE(_09953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17689__C1 (.DIODE(_09953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17682__C1 (.DIODE(_09953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17675__C1 (.DIODE(_09953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17668__C1 (.DIODE(_09953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17661__C1 (.DIODE(_09953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17654__C1 (.DIODE(_09953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17647__C1 (.DIODE(_09953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17639__C1 (.DIODE(_09953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17706__A1 (.DIODE(_09956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17699__A1 (.DIODE(_09956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17692__A1 (.DIODE(_09956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17685__A1 (.DIODE(_09956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17678__A1 (.DIODE(_09956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17671__A1 (.DIODE(_09956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17664__A1 (.DIODE(_09956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17657__A1 (.DIODE(_09956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17650__A1 (.DIODE(_09956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17643__A1 (.DIODE(_09956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17828__S (.DIODE(_10027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17825__S (.DIODE(_10027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17822__S (.DIODE(_10027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17819__S (.DIODE(_10027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17816__S (.DIODE(_10027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17813__S (.DIODE(_10027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17810__S (.DIODE(_10027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17778__A (.DIODE(_10027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17728__B1 (.DIODE(_10027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17725__B (.DIODE(_10027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17775__B1 (.DIODE(_10028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17772__B1 (.DIODE(_10028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17769__B1 (.DIODE(_10028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17766__B1 (.DIODE(_10028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17762__B1 (.DIODE(_10028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17726__A (.DIODE(_10028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17829__S (.DIODE(_10033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17826__S (.DIODE(_10033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17795__A (.DIODE(_10033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17763__A (.DIODE(_10033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17732__A (.DIODE(_10033_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(dout1[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(dout1[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(dout1[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(dout1[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(dout1[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(dout1[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(dout1[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(dout1[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(dout1[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(dout1[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(dout1[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(dout1[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(dout1[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(dout1[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(dout1[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(dout1[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(dout1[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(dout1[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(dout1[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(dout1[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(dout1[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(dout1[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(dout1[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(dout1[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(dout1[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(dout1[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(dout1[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(dout1[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(dout1[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(dout1[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(dout1[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(dout1[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(io_wbs_adr[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(io_wbs_adr[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(io_wbs_adr[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(io_wbs_adr[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(io_wbs_adr[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(io_wbs_adr[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(io_wbs_adr[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(io_wbs_adr[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(io_wbs_adr[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(io_wbs_adr[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(io_wbs_adr[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(io_wbs_adr[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(io_wbs_adr[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(io_wbs_adr[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(io_wbs_adr[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(io_wbs_adr[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(io_wbs_adr[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(io_wbs_adr[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(io_wbs_adr[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(io_wbs_adr[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(io_wbs_adr[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(io_wbs_adr[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(io_wbs_adr[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(io_wbs_adr[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(io_wbs_adr[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(io_wbs_adr[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(io_wbs_adr[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(io_wbs_adr[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(io_wbs_adr[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(io_wbs_adr[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(io_wbs_adr[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(io_wbs_adr[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_io_wbs_clk_A (.DIODE(io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(io_wbs_cyc));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(io_wbs_datwr[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(io_wbs_datwr[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(io_wbs_datwr[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(io_wbs_datwr[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(io_wbs_datwr[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(io_wbs_datwr[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(io_wbs_datwr[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(io_wbs_datwr[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(io_wbs_datwr[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(io_wbs_datwr[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(io_wbs_datwr[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(io_wbs_datwr[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(io_wbs_datwr[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(io_wbs_datwr[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(io_wbs_datwr[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(io_wbs_datwr[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(io_wbs_datwr[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(io_wbs_datwr[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(io_wbs_datwr[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(io_wbs_datwr[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(io_wbs_datwr[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(io_wbs_datwr[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(io_wbs_datwr[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(io_wbs_datwr[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(io_wbs_datwr[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(io_wbs_datwr[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(io_wbs_datwr[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(io_wbs_datwr[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(io_wbs_datwr[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(io_wbs_datwr[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(io_wbs_datwr[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(io_wbs_datwr[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_A (.DIODE(io_wbs_rst));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_A (.DIODE(io_wbs_stb));
 sky130_fd_sc_hd__diode_2 ANTENNA_input100_A (.DIODE(io_wbs_we));
 sky130_fd_sc_hd__diode_2 ANTENNA__20042__A1 (.DIODE(\wfg_core_top.active_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18108__A (.DIODE(\wfg_core_top.active_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18098__C1 (.DIODE(\wfg_core_top.active_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18095__C1 (.DIODE(\wfg_core_top.active_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18064__A (.DIODE(\wfg_core_top.active_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17896__A1 (.DIODE(\wfg_core_top.active_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17884__A (.DIODE(\wfg_core_top.active_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17881__B1 (.DIODE(\wfg_core_top.active_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17838__A (.DIODE(\wfg_core_top.active_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17836__C (.DIODE(\wfg_core_top.active_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20073__A1 (.DIODE(\wfg_core_top.cfg_subcycle_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18246__A1 (.DIODE(\wfg_core_top.cfg_subcycle_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18077__A1 (.DIODE(\wfg_core_top.cfg_subcycle_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20075__A1 (.DIODE(\wfg_core_top.cfg_subcycle_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18250__A1 (.DIODE(\wfg_core_top.cfg_subcycle_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18080__A1 (.DIODE(\wfg_core_top.cfg_subcycle_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20078__A1 (.DIODE(\wfg_core_top.cfg_subcycle_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18254__A1 (.DIODE(\wfg_core_top.cfg_subcycle_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18083__A1 (.DIODE(\wfg_core_top.cfg_subcycle_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20047__A1 (.DIODE(\wfg_core_top.cfg_sync_q[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18292__A1 (.DIODE(\wfg_core_top.cfg_sync_q[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17911__A1 (.DIODE(\wfg_core_top.cfg_sync_q[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20049__A1 (.DIODE(\wfg_core_top.cfg_sync_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18296__A1 (.DIODE(\wfg_core_top.cfg_sync_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17907__B2 (.DIODE(\wfg_core_top.cfg_sync_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20051__A1 (.DIODE(\wfg_core_top.cfg_sync_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18300__A1 (.DIODE(\wfg_core_top.cfg_sync_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17904__B2 (.DIODE(\wfg_core_top.cfg_sync_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20056__A1 (.DIODE(\wfg_core_top.cfg_sync_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18308__A1 (.DIODE(\wfg_core_top.cfg_sync_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17898__B2 (.DIODE(\wfg_core_top.cfg_sync_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20058__A1 (.DIODE(\wfg_core_top.cfg_sync_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18313__A1 (.DIODE(\wfg_core_top.cfg_sync_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17895__A1 (.DIODE(\wfg_core_top.cfg_sync_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20068__A1 (.DIODE(\wfg_core_top.wbs_dat_o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17998__A1 (.DIODE(\wfg_core_top.wbs_dat_o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20074__A1 (.DIODE(\wfg_core_top.wbs_dat_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18004__A1 (.DIODE(\wfg_core_top.wbs_dat_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18196__A0 (.DIODE(\wfg_core_top.wfg_core.temp_subcycle ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17886__S (.DIODE(\wfg_core_top.wfg_core.temp_subcycle ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17834__B (.DIODE(\wfg_core_top.wfg_core.temp_subcycle ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18198__A0 (.DIODE(\wfg_core_top.wfg_core.temp_sync ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17882__A1 (.DIODE(\wfg_core_top.wfg_core.temp_sync ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17881__A1 (.DIODE(\wfg_core_top.wfg_core.temp_sync ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10062__B (.DIODE(\wfg_core_top.wfg_core.temp_sync ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18769__A1 (.DIODE(\wfg_drive_pat_top.cfg_begin_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18520__A1 (.DIODE(\wfg_drive_pat_top.cfg_begin_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17478__B2 (.DIODE(\wfg_drive_pat_top.cfg_begin_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17477__A2_N (.DIODE(\wfg_drive_pat_top.cfg_begin_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18854__A1 (.DIODE(\wfg_drive_pat_top.patsel0_low_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18573__B2 (.DIODE(\wfg_drive_pat_top.patsel0_low_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17610__A_N (.DIODE(\wfg_drive_pat_top.patsel0_low_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17608__A1 (.DIODE(\wfg_drive_pat_top.patsel0_low_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18812__A1 (.DIODE(\wfg_drive_pat_top.patsel0_low_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18516__B2 (.DIODE(\wfg_drive_pat_top.patsel0_low_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17506__A_N (.DIODE(\wfg_drive_pat_top.patsel0_low_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17504__A1 (.DIODE(\wfg_drive_pat_top.patsel0_low_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18834__A1 (.DIODE(\wfg_drive_pat_top.patsel0_low_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18547__B2 (.DIODE(\wfg_drive_pat_top.patsel0_low_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17492__A_N (.DIODE(\wfg_drive_pat_top.patsel0_low_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17474__A1 (.DIODE(\wfg_drive_pat_top.patsel0_low_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18916__A1 (.DIODE(\wfg_drive_pat_top.patsel1_high_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18515__B2 (.DIODE(\wfg_drive_pat_top.patsel1_high_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17506__C (.DIODE(\wfg_drive_pat_top.patsel1_high_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17503__A (.DIODE(\wfg_drive_pat_top.patsel1_high_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18938__A1 (.DIODE(\wfg_drive_pat_top.patsel1_high_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18548__A1 (.DIODE(\wfg_drive_pat_top.patsel1_high_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17492__C (.DIODE(\wfg_drive_pat_top.patsel1_high_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17471__A (.DIODE(\wfg_drive_pat_top.patsel1_high_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18504__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17943__B2 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18566__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18006__A (.DIODE(\wfg_drive_pat_top.wbs_dat_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18570__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18009__A (.DIODE(\wfg_drive_pat_top.wbs_dat_o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18579__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18015__A (.DIODE(\wfg_drive_pat_top.wbs_dat_o[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18587__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18018__A (.DIODE(\wfg_drive_pat_top.wbs_dat_o[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18592__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18021__B2 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18597__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18025__B2 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18602__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18029__B2 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18605__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18033__B2 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18610__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18037__B2 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18613__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18041__B2 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18617__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18047__A (.DIODE(\wfg_drive_pat_top.wbs_dat_o[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18620__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18049__A (.DIODE(\wfg_drive_pat_top.wbs_dat_o[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18625__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18051__A (.DIODE(\wfg_drive_pat_top.wbs_dat_o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18628__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18053__A (.DIODE(\wfg_drive_pat_top.wbs_dat_o[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18631__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18055__A (.DIODE(\wfg_drive_pat_top.wbs_dat_o[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18636__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18057__A (.DIODE(\wfg_drive_pat_top.wbs_dat_o[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18641__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18059__A (.DIODE(\wfg_drive_pat_top.wbs_dat_o[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18646__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18061__A (.DIODE(\wfg_drive_pat_top.wbs_dat_o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18522__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17968__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18526__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17973__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18535__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17981__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18540__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17984__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18545__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17989__A (.DIODE(\wfg_drive_pat_top.wbs_dat_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18549__A1 (.DIODE(\wfg_drive_pat_top.wbs_dat_o[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17992__A (.DIODE(\wfg_drive_pat_top.wbs_dat_o[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17799__A0 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[10].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17648__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[10].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17646__B (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[10].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17796__A0 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[11].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17640__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[11].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17636__B (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[11].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17792__A0 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[12].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17630__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[12].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17628__B (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[12].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17789__A0 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[13].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17623__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[13].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17621__B (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[13].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17786__A0 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[14].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17616__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[14].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17614__B (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[14].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17783__A0 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[15].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17609__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[15].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17607__B (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[15].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17780__A0 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[16].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17601__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[16].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17599__B (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[16].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17776__A0 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[17].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17594__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[17].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17592__B (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[17].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17773__A0 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[18].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17587__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[18].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17585__B (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[18].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17770__A0 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[19].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17718__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[19].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17716__B (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[19].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17767__A0 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[20].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17573__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[20].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17571__B (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[20].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17764__A0 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[21].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17565__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[21].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17561__B (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[21].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17760__A0 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[22].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17555__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[22].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17553__B (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[22].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17757__A0 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[23].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17548__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[23].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17546__B (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[23].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17748__A0 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[26].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17526__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[26].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17524__B (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[26].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17739__A0 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[29].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17711__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[29].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17709__B (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[29].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18659__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[2].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18515__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[2].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17507__B1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[2].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17505__C1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[2].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17733__A0 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[31].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17704__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[31].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17702__B (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[31].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17820__A0 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[3].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17697__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[3].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17695__B (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[3].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17817__A0 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[4].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17690__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[4].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17688__B (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[4].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17814__A0 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[5].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17683__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[5].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17681__B (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[5].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18668__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[5].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18528__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[5].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17685__B1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[5].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17683__C1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[5].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17811__A0 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[6].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17676__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[6].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17674__B (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[6].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17808__A0 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[7].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17669__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[7].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17667__B (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[7].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17805__A0 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[8].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17662__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[8].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17660__B (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[8].drv.axis_data_ff ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18681__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[9].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18546__A1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[9].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17493__B1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[9].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17475__C1 (.DIODE(\wfg_drive_pat_top.wfg_drive_pat.gen_channels[9].drv.ctrl_en_q_i ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20108__A (.DIODE(\wfg_drive_spi_top.cfg_cpol_q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19205__A1 (.DIODE(\wfg_drive_spi_top.cfg_cpol_q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10082__A0 (.DIODE(\wfg_drive_spi_top.cfg_cpol_q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20110__A (.DIODE(\wfg_drive_spi_top.cfg_dff_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19209__B2 (.DIODE(\wfg_drive_spi_top.cfg_dff_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10078__A0 (.DIODE(\wfg_drive_spi_top.cfg_dff_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20114__A (.DIODE(\wfg_drive_spi_top.cfg_lsbfirst_q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19207__B2 (.DIODE(\wfg_drive_spi_top.cfg_lsbfirst_q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10085__A0 (.DIODE(\wfg_drive_spi_top.cfg_lsbfirst_q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20116__A (.DIODE(\wfg_drive_spi_top.cfg_sspol_q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19213__B2 (.DIODE(\wfg_drive_spi_top.cfg_sspol_q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10080__A0 (.DIODE(\wfg_drive_spi_top.cfg_sspol_q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20121__A (.DIODE(\wfg_drive_spi_top.clkcfg_div_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19204__A1 (.DIODE(\wfg_drive_spi_top.clkcfg_div_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10275__A0 (.DIODE(\wfg_drive_spi_top.clkcfg_div_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20123__A (.DIODE(\wfg_drive_spi_top.clkcfg_div_q[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19207__A1 (.DIODE(\wfg_drive_spi_top.clkcfg_div_q[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10273__A0 (.DIODE(\wfg_drive_spi_top.clkcfg_div_q[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20125__A (.DIODE(\wfg_drive_spi_top.clkcfg_div_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19209__A1 (.DIODE(\wfg_drive_spi_top.clkcfg_div_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10271__A0 (.DIODE(\wfg_drive_spi_top.clkcfg_div_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20127__A (.DIODE(\wfg_drive_spi_top.clkcfg_div_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19211__A1 (.DIODE(\wfg_drive_spi_top.clkcfg_div_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10269__A0 (.DIODE(\wfg_drive_spi_top.clkcfg_div_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20131__A (.DIODE(\wfg_drive_spi_top.clkcfg_div_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19215__A1 (.DIODE(\wfg_drive_spi_top.clkcfg_div_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10265__A0 (.DIODE(\wfg_drive_spi_top.clkcfg_div_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19210__A1 (.DIODE(\wfg_drive_spi_top.wbs_dat_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17966__A1 (.DIODE(\wfg_drive_spi_top.wbs_dat_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19212__A1 (.DIODE(\wfg_drive_spi_top.wbs_dat_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17969__A1 (.DIODE(\wfg_drive_spi_top.wbs_dat_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19214__A1 (.DIODE(\wfg_drive_spi_top.wbs_dat_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17975__A1 (.DIODE(\wfg_drive_spi_top.wbs_dat_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19216__A1 (.DIODE(\wfg_drive_spi_top.wbs_dat_o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17977__A1 (.DIODE(\wfg_drive_spi_top.wbs_dat_o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19217__A (.DIODE(\wfg_drive_spi_top.wbs_dat_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17983__A1 (.DIODE(\wfg_drive_spi_top.wbs_dat_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19221__A (.DIODE(\wfg_drive_spi_top.wbs_dat_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17985__A1 (.DIODE(\wfg_drive_spi_top.wbs_dat_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13859__A1 (.DIODE(\wfg_drive_spi_top.wfg_axis_tready_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13396__A1 (.DIODE(\wfg_drive_spi_top.wfg_axis_tready_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10087__A0 (.DIODE(\wfg_drive_spi_top.wfg_axis_tready_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18160__S0 (.DIODE(\wfg_drive_spi_top.wfg_drive_spi.byte_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10251__A (.DIODE(\wfg_drive_spi_top.wfg_drive_spi.byte_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10078__A1 (.DIODE(\wfg_drive_spi_top.wfg_drive_spi.byte_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18160__S1 (.DIODE(\wfg_drive_spi_top.wfg_drive_spi.byte_cnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10250__A1 (.DIODE(\wfg_drive_spi_top.wfg_drive_spi.byte_cnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10075__A1 (.DIODE(\wfg_drive_spi_top.wfg_drive_spi.byte_cnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10242__S (.DIODE(\wfg_drive_spi_top.wfg_drive_spi.lsbfirst ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10238__S (.DIODE(\wfg_drive_spi_top.wfg_drive_spi.lsbfirst ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10234__S (.DIODE(\wfg_drive_spi_top.wfg_drive_spi.lsbfirst ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10191__A (.DIODE(\wfg_drive_spi_top.wfg_drive_spi.lsbfirst ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10142__A (.DIODE(\wfg_drive_spi_top.wfg_drive_spi.lsbfirst ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10084__A (.DIODE(\wfg_drive_spi_top.wfg_drive_spi.lsbfirst ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18161__A0 (.DIODE(\wfg_drive_spi_top.wfg_drive_spi.spi_data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10248__B2 (.DIODE(\wfg_drive_spi_top.wfg_drive_spi.spi_data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10242__A0 (.DIODE(\wfg_drive_spi_top.wfg_drive_spi.spi_data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18160__A2 (.DIODE(\wfg_drive_spi_top.wfg_drive_spi.spi_data[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10147__A1 (.DIODE(\wfg_drive_spi_top.wfg_drive_spi.spi_data[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10145__A1 (.DIODE(\wfg_drive_spi_top.wfg_drive_spi.spi_data[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10138__A0 (.DIODE(\wfg_drive_spi_top.wfg_drive_spi.spi_data[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18160__A3 (.DIODE(\wfg_drive_spi_top.wfg_drive_spi.spi_data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10112__A1 (.DIODE(\wfg_drive_spi_top.wfg_drive_spi.spi_data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10110__A1 (.DIODE(\wfg_drive_spi_top.wfg_drive_spi.spi_data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19773__B2 (.DIODE(\wfg_interconnect_top.driver0_select_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10175__B (.DIODE(\wfg_interconnect_top.driver0_select_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10105__A2 (.DIODE(\wfg_interconnect_top.driver0_select_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10065__A2 (.DIODE(\wfg_interconnect_top.driver0_select_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10058__A (.DIODE(\wfg_interconnect_top.driver0_select_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17828__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17112__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10246__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17798__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17092__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10208__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17791__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17088__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10199__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17788__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17086__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10194__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17785__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17084__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10188__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17782__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17082__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10184__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17779__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17079__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10180__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17725__A (.DIODE(\wfg_interconnect_top.stimulus_0[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17072__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10105__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17825__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17110__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10244__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17822__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17108__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10240__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17728__B2 (.DIODE(\wfg_interconnect_top.stimulus_0[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10065__A3 (.DIODE(\wfg_interconnect_top.stimulus_0[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17819__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17106__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10236__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17816__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17104__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10232__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17813__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17102__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10228__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17810__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17100__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10224__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17807__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17098__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10220__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17804__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17096__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10216__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17801__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17094__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10212__A1 (.DIODE(\wfg_interconnect_top.stimulus_0[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17728__A1 (.DIODE(\wfg_interconnect_top.stimulus_1[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10061__A2 (.DIODE(\wfg_interconnect_top.stimulus_1[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13017__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10323__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12926__B (.DIODE(\wfg_stim_mem_top.cfg_gain_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12300__B (.DIODE(\wfg_stim_mem_top.cfg_gain_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11805__B (.DIODE(\wfg_stim_mem_top.cfg_gain_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11644__B (.DIODE(\wfg_stim_mem_top.cfg_gain_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11290__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11273__B (.DIODE(\wfg_stim_mem_top.cfg_gain_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11054__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10316__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10313__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12926__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12896__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12300__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11805__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11644__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11289__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11273__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11053__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11050__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10311__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12339__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12211__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11719__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11635__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11553__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11264__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11261__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10946__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10343__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10334__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11637__B (.DIODE(\wfg_stim_mem_top.cfg_gain_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10629__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10626__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10339__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12426__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12276__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11620__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11211__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10351__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12275__B (.DIODE(\wfg_stim_mem_top.cfg_gain_q[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11619__B (.DIODE(\wfg_stim_mem_top.cfg_gain_q[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11209__B (.DIODE(\wfg_stim_mem_top.cfg_gain_q[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10357__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10354__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12416__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12359__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12265__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12184__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11770__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11691__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11609__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11526__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11199__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10365__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12266__B (.DIODE(\wfg_stim_mem_top.cfg_gain_q[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11610__B (.DIODE(\wfg_stim_mem_top.cfg_gain_q[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11190__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10371__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12263__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12262__B2 (.DIODE(\wfg_stim_mem_top.cfg_gain_q[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12182__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11524__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11173__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11095__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10430__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13017__B (.DIODE(\wfg_stim_mem_top.cfg_gain_q[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10303__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13030__B (.DIODE(\wfg_stim_mem_top.cfg_gain_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12993__B (.DIODE(\wfg_stim_mem_top.cfg_gain_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12964__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12924__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12894__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11642__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10907__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10309__A (.DIODE(\wfg_stim_mem_top.cfg_gain_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19835__A1 (.DIODE(\wfg_stim_mem_top.cfg_inc_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19418__B2 (.DIODE(\wfg_stim_mem_top.cfg_inc_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13718__A (.DIODE(\wfg_stim_mem_top.cfg_inc_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13673__A (.DIODE(\wfg_stim_mem_top.cfg_inc_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19844__A1 (.DIODE(\wfg_stim_mem_top.cfg_inc_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19435__A1 (.DIODE(\wfg_stim_mem_top.cfg_inc_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13713__A (.DIODE(\wfg_stim_mem_top.cfg_inc_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13678__A1 (.DIODE(\wfg_stim_mem_top.cfg_inc_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13677__A1 (.DIODE(\wfg_stim_mem_top.cfg_inc_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19862__A1 (.DIODE(\wfg_stim_mem_top.end_val_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19417__B2 (.DIODE(\wfg_stim_mem_top.end_val_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13720__C1 (.DIODE(\wfg_stim_mem_top.end_val_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19872__A1 (.DIODE(\wfg_stim_mem_top.end_val_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19434__B2 (.DIODE(\wfg_stim_mem_top.end_val_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13724__B2 (.DIODE(\wfg_stim_mem_top.end_val_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13723__A1 (.DIODE(\wfg_stim_mem_top.end_val_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19915__A1 (.DIODE(\wfg_stim_mem_top.start_val_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19418__A1 (.DIODE(\wfg_stim_mem_top.start_val_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13802__A (.DIODE(\wfg_stim_mem_top.start_val_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19923__A1 (.DIODE(\wfg_stim_mem_top.start_val_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19434__A1 (.DIODE(\wfg_stim_mem_top.start_val_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13790__A1 (.DIODE(\wfg_stim_mem_top.start_val_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19457__A1 (.DIODE(\wfg_stim_mem_top.wbs_dat_o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17999__B2 (.DIODE(\wfg_stim_mem_top.wbs_dat_o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19461__A1 (.DIODE(\wfg_stim_mem_top.wbs_dat_o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18002__B2 (.DIODE(\wfg_stim_mem_top.wbs_dat_o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19464__A1 (.DIODE(\wfg_stim_mem_top.wbs_dat_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18005__B2 (.DIODE(\wfg_stim_mem_top.wbs_dat_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19467__A1 (.DIODE(\wfg_stim_mem_top.wbs_dat_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18008__B2 (.DIODE(\wfg_stim_mem_top.wbs_dat_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19470__A1 (.DIODE(\wfg_stim_mem_top.wbs_dat_o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18011__B2 (.DIODE(\wfg_stim_mem_top.wbs_dat_o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19473__A1 (.DIODE(\wfg_stim_mem_top.wbs_dat_o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18014__B2 (.DIODE(\wfg_stim_mem_top.wbs_dat_o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19428__A1 (.DIODE(\wfg_stim_mem_top.wbs_dat_o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17960__B2 (.DIODE(\wfg_stim_mem_top.wbs_dat_o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19431__A1 (.DIODE(\wfg_stim_mem_top.wbs_dat_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17964__B2 (.DIODE(\wfg_stim_mem_top.wbs_dat_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19436__A1 (.DIODE(\wfg_stim_mem_top.wbs_dat_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17968__B2 (.DIODE(\wfg_stim_mem_top.wbs_dat_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19439__A1 (.DIODE(\wfg_stim_mem_top.wbs_dat_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17973__B2 (.DIODE(\wfg_stim_mem_top.wbs_dat_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19445__A1 (.DIODE(\wfg_stim_mem_top.wbs_dat_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17981__B2 (.DIODE(\wfg_stim_mem_top.wbs_dat_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19448__A1 (.DIODE(\wfg_stim_mem_top.wbs_dat_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17984__B2 (.DIODE(\wfg_stim_mem_top.wbs_dat_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19454__A1 (.DIODE(\wfg_stim_mem_top.wbs_dat_o[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17994__B2 (.DIODE(\wfg_stim_mem_top.wbs_dat_o[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17916__B1 (.DIODE(\wfg_stim_mem_top.wfg_stim_mem.cur_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13741__A2 (.DIODE(\wfg_stim_mem_top.wfg_stim_mem.cur_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13392__B (.DIODE(\wfg_stim_mem_top.wfg_stim_mem.cur_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13658__S (.DIODE(\wfg_stim_mem_top.wfg_stim_mem.cur_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13656__S (.DIODE(\wfg_stim_mem_top.wfg_stim_mem.cur_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13635__A (.DIODE(\wfg_stim_mem_top.wfg_stim_mem.cur_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13614__A (.DIODE(\wfg_stim_mem_top.wfg_stim_mem.cur_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13593__A (.DIODE(\wfg_stim_mem_top.wfg_stim_mem.cur_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13398__B1 (.DIODE(\wfg_stim_mem_top.wfg_stim_mem.cur_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20200__D (.DIODE(\wfg_stim_mem_top.wfg_stim_mem.cur_state[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13741__A1 (.DIODE(\wfg_stim_mem_top.wfg_stim_mem.cur_state[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13737__B1 (.DIODE(\wfg_stim_mem_top.wfg_stim_mem.cur_state[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13399__C_N (.DIODE(\wfg_stim_mem_top.wfg_stim_mem.cur_state[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13658__A1 (.DIODE(\wfg_stim_mem_top.wfg_stim_mem.data_calc[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13592__A1 (.DIODE(\wfg_stim_mem_top.wfg_stim_mem.data_calc[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13608__A1 (.DIODE(\wfg_stim_mem_top.wfg_stim_mem.data_calc[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13494__A1 (.DIODE(\wfg_stim_mem_top.wfg_stim_mem.data_calc[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13606__A1 (.DIODE(\wfg_stim_mem_top.wfg_stim_mem.data_calc[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13491__A1 (.DIODE(\wfg_stim_mem_top.wfg_stim_mem.data_calc[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13600__A1 (.DIODE(\wfg_stim_mem_top.wfg_stim_mem.data_calc[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13477__A1 (.DIODE(\wfg_stim_mem_top.wfg_stim_mem.data_calc[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19068__A1 (.DIODE(\wfg_stim_sine_top.ctrl_en_q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17241__A1 (.DIODE(\wfg_stim_sine_top.ctrl_en_q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17237__A (.DIODE(\wfg_stim_sine_top.ctrl_en_q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15083__A1 (.DIODE(\wfg_stim_sine_top.gain_val_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14559__A (.DIODE(\wfg_stim_sine_top.gain_val_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14557__B (.DIODE(\wfg_stim_sine_top.gain_val_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14055__A (.DIODE(\wfg_stim_sine_top.gain_val_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14052__B (.DIODE(\wfg_stim_sine_top.gain_val_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14800__B (.DIODE(\wfg_stim_sine_top.gain_val_q[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14534__A1 (.DIODE(\wfg_stim_sine_top.gain_val_q[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14524__A (.DIODE(\wfg_stim_sine_top.gain_val_q[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14513__A (.DIODE(\wfg_stim_sine_top.gain_val_q[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13966__A (.DIODE(\wfg_stim_sine_top.gain_val_q[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14508__B (.DIODE(\wfg_stim_sine_top.gain_val_q[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13954__A (.DIODE(\wfg_stim_sine_top.gain_val_q[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14755__A (.DIODE(\wfg_stim_sine_top.gain_val_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14662__A (.DIODE(\wfg_stim_sine_top.gain_val_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14597__B2 (.DIODE(\wfg_stim_sine_top.gain_val_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14596__A (.DIODE(\wfg_stim_sine_top.gain_val_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14521__A (.DIODE(\wfg_stim_sine_top.gain_val_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14520__B2 (.DIODE(\wfg_stim_sine_top.gain_val_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14509__B2 (.DIODE(\wfg_stim_sine_top.gain_val_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14508__A (.DIODE(\wfg_stim_sine_top.gain_val_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13962__A (.DIODE(\wfg_stim_sine_top.gain_val_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13960__A (.DIODE(\wfg_stim_sine_top.gain_val_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14863__A (.DIODE(\wfg_stim_sine_top.gain_val_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14748__A (.DIODE(\wfg_stim_sine_top.gain_val_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14655__A (.DIODE(\wfg_stim_sine_top.gain_val_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14590__A (.DIODE(\wfg_stim_sine_top.gain_val_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14518__A1 (.DIODE(\wfg_stim_sine_top.gain_val_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14262__C (.DIODE(\wfg_stim_sine_top.gain_val_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14190__B (.DIODE(\wfg_stim_sine_top.gain_val_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13935__A (.DIODE(\wfg_stim_sine_top.gain_val_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14862__A1 (.DIODE(\wfg_stim_sine_top.gain_val_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14861__B (.DIODE(\wfg_stim_sine_top.gain_val_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14747__A1 (.DIODE(\wfg_stim_sine_top.gain_val_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14653__B (.DIODE(\wfg_stim_sine_top.gain_val_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14589__A1 (.DIODE(\wfg_stim_sine_top.gain_val_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14267__B (.DIODE(\wfg_stim_sine_top.gain_val_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14256__B (.DIODE(\wfg_stim_sine_top.gain_val_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13975__A (.DIODE(\wfg_stim_sine_top.gain_val_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13928__A (.DIODE(\wfg_stim_sine_top.gain_val_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14862__B2 (.DIODE(\wfg_stim_sine_top.gain_val_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14861__A (.DIODE(\wfg_stim_sine_top.gain_val_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14747__B2 (.DIODE(\wfg_stim_sine_top.gain_val_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14653__A (.DIODE(\wfg_stim_sine_top.gain_val_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14267__A (.DIODE(\wfg_stim_sine_top.gain_val_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14256__A (.DIODE(\wfg_stim_sine_top.gain_val_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13974__A (.DIODE(\wfg_stim_sine_top.gain_val_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13921__A (.DIODE(\wfg_stim_sine_top.gain_val_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15083__B2 (.DIODE(\wfg_stim_sine_top.gain_val_q[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14560__A (.DIODE(\wfg_stim_sine_top.gain_val_q[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14557__A (.DIODE(\wfg_stim_sine_top.gain_val_q[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14054__A (.DIODE(\wfg_stim_sine_top.gain_val_q[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14052__A (.DIODE(\wfg_stim_sine_top.gain_val_q[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15226__A (.DIODE(\wfg_stim_sine_top.gain_val_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15187__A (.DIODE(\wfg_stim_sine_top.gain_val_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15128__A (.DIODE(\wfg_stim_sine_top.gain_val_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15120__A (.DIODE(\wfg_stim_sine_top.gain_val_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15080__A (.DIODE(\wfg_stim_sine_top.gain_val_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15026__A (.DIODE(\wfg_stim_sine_top.gain_val_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14556__A (.DIODE(\wfg_stim_sine_top.gain_val_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14120__A (.DIODE(\wfg_stim_sine_top.gain_val_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14058__A (.DIODE(\wfg_stim_sine_top.gain_val_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15191__A (.DIODE(\wfg_stim_sine_top.gain_val_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15132__A (.DIODE(\wfg_stim_sine_top.gain_val_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15112__A (.DIODE(\wfg_stim_sine_top.gain_val_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15074__A (.DIODE(\wfg_stim_sine_top.gain_val_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15020__A (.DIODE(\wfg_stim_sine_top.gain_val_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14816__A (.DIODE(\wfg_stim_sine_top.gain_val_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14730__A (.DIODE(\wfg_stim_sine_top.gain_val_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14546__A (.DIODE(\wfg_stim_sine_top.gain_val_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14060__A (.DIODE(\wfg_stim_sine_top.gain_val_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15134__B (.DIODE(\wfg_stim_sine_top.gain_val_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15133__A1 (.DIODE(\wfg_stim_sine_top.gain_val_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15076__B (.DIODE(\wfg_stim_sine_top.gain_val_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15022__B (.DIODE(\wfg_stim_sine_top.gain_val_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15021__A1 (.DIODE(\wfg_stim_sine_top.gain_val_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14818__B (.DIODE(\wfg_stim_sine_top.gain_val_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14817__A1 (.DIODE(\wfg_stim_sine_top.gain_val_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14728__B (.DIODE(\wfg_stim_sine_top.gain_val_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14446__A (.DIODE(\wfg_stim_sine_top.gain_val_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14064__A (.DIODE(\wfg_stim_sine_top.gain_val_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15134__A (.DIODE(\wfg_stim_sine_top.gain_val_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15022__A (.DIODE(\wfg_stim_sine_top.gain_val_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15021__B2 (.DIODE(\wfg_stim_sine_top.gain_val_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14818__A (.DIODE(\wfg_stim_sine_top.gain_val_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14817__B2 (.DIODE(\wfg_stim_sine_top.gain_val_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14728__A (.DIODE(\wfg_stim_sine_top.gain_val_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14445__A (.DIODE(\wfg_stim_sine_top.gain_val_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14062__A (.DIODE(\wfg_stim_sine_top.gain_val_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14532__A (.DIODE(\wfg_stim_sine_top.gain_val_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14000__A (.DIODE(\wfg_stim_sine_top.gain_val_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15060__B (.DIODE(\wfg_stim_sine_top.gain_val_q[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15005__A1 (.DIODE(\wfg_stim_sine_top.gain_val_q[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15004__B (.DIODE(\wfg_stim_sine_top.gain_val_q[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14804__A1 (.DIODE(\wfg_stim_sine_top.gain_val_q[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14803__B (.DIODE(\wfg_stim_sine_top.gain_val_q[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14607__B (.DIODE(\wfg_stim_sine_top.gain_val_q[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14531__A1 (.DIODE(\wfg_stim_sine_top.gain_val_q[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14530__B (.DIODE(\wfg_stim_sine_top.gain_val_q[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14006__A (.DIODE(\wfg_stim_sine_top.gain_val_q[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14004__A (.DIODE(\wfg_stim_sine_top.gain_val_q[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15060__A (.DIODE(\wfg_stim_sine_top.gain_val_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15005__B2 (.DIODE(\wfg_stim_sine_top.gain_val_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15004__A (.DIODE(\wfg_stim_sine_top.gain_val_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14803__A (.DIODE(\wfg_stim_sine_top.gain_val_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14531__B2 (.DIODE(\wfg_stim_sine_top.gain_val_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14530__A (.DIODE(\wfg_stim_sine_top.gain_val_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14229__A (.DIODE(\wfg_stim_sine_top.gain_val_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14003__A (.DIODE(\wfg_stim_sine_top.gain_val_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19567__A1 (.DIODE(\wfg_stim_sine_top.inc_val_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19065__A1 (.DIODE(\wfg_stim_sine_top.inc_val_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13916__A (.DIODE(\wfg_stim_sine_top.inc_val_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13824__A (.DIODE(\wfg_stim_sine_top.inc_val_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19598__A1 (.DIODE(\wfg_stim_sine_top.inc_val_q[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19107__B2 (.DIODE(\wfg_stim_sine_top.inc_val_q[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13846__A (.DIODE(\wfg_stim_sine_top.inc_val_q[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13812__A (.DIODE(\wfg_stim_sine_top.inc_val_q[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19601__A1 (.DIODE(\wfg_stim_sine_top.inc_val_q[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19111__B2 (.DIODE(\wfg_stim_sine_top.inc_val_q[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13848__A (.DIODE(\wfg_stim_sine_top.inc_val_q[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13811__A (.DIODE(\wfg_stim_sine_top.inc_val_q[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19604__A1 (.DIODE(\wfg_stim_sine_top.inc_val_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19114__B2 (.DIODE(\wfg_stim_sine_top.inc_val_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13850__A (.DIODE(\wfg_stim_sine_top.inc_val_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13810__A (.DIODE(\wfg_stim_sine_top.inc_val_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19607__A1 (.DIODE(\wfg_stim_sine_top.inc_val_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19117__B2 (.DIODE(\wfg_stim_sine_top.inc_val_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13869__A (.DIODE(\wfg_stim_sine_top.inc_val_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13853__A1 (.DIODE(\wfg_stim_sine_top.inc_val_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13852__A1 (.DIODE(\wfg_stim_sine_top.inc_val_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19610__A1 (.DIODE(\wfg_stim_sine_top.inc_val_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19120__B2 (.DIODE(\wfg_stim_sine_top.inc_val_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13808__A (.DIODE(\wfg_stim_sine_top.inc_val_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13807__A (.DIODE(\wfg_stim_sine_top.inc_val_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19613__A1 (.DIODE(\wfg_stim_sine_top.inc_val_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19123__B2 (.DIODE(\wfg_stim_sine_top.inc_val_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13806__A (.DIODE(\wfg_stim_sine_top.inc_val_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19570__A1 (.DIODE(\wfg_stim_sine_top.inc_val_q[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19078__B2 (.DIODE(\wfg_stim_sine_top.inc_val_q[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13826__A (.DIODE(\wfg_stim_sine_top.inc_val_q[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13825__A (.DIODE(\wfg_stim_sine_top.inc_val_q[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19573__A1 (.DIODE(\wfg_stim_sine_top.inc_val_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19083__B2 (.DIODE(\wfg_stim_sine_top.inc_val_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13829__A (.DIODE(\wfg_stim_sine_top.inc_val_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13823__A (.DIODE(\wfg_stim_sine_top.inc_val_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19576__A1 (.DIODE(\wfg_stim_sine_top.inc_val_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19086__B2 (.DIODE(\wfg_stim_sine_top.inc_val_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13903__A (.DIODE(\wfg_stim_sine_top.inc_val_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13831__A1 (.DIODE(\wfg_stim_sine_top.inc_val_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13822__A (.DIODE(\wfg_stim_sine_top.inc_val_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19579__A1 (.DIODE(\wfg_stim_sine_top.inc_val_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19089__B2 (.DIODE(\wfg_stim_sine_top.inc_val_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13821__A (.DIODE(\wfg_stim_sine_top.inc_val_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13820__A (.DIODE(\wfg_stim_sine_top.inc_val_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19582__A1 (.DIODE(\wfg_stim_sine_top.inc_val_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19092__B2 (.DIODE(\wfg_stim_sine_top.inc_val_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13833__A (.DIODE(\wfg_stim_sine_top.inc_val_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13819__A (.DIODE(\wfg_stim_sine_top.inc_val_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19586__A1 (.DIODE(\wfg_stim_sine_top.inc_val_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19095__B2 (.DIODE(\wfg_stim_sine_top.inc_val_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13837__A (.DIODE(\wfg_stim_sine_top.inc_val_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13818__A (.DIODE(\wfg_stim_sine_top.inc_val_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19589__A1 (.DIODE(\wfg_stim_sine_top.inc_val_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19098__B2 (.DIODE(\wfg_stim_sine_top.inc_val_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13839__A (.DIODE(\wfg_stim_sine_top.inc_val_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13817__A (.DIODE(\wfg_stim_sine_top.inc_val_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19592__A1 (.DIODE(\wfg_stim_sine_top.inc_val_q[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19101__B2 (.DIODE(\wfg_stim_sine_top.inc_val_q[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13816__A (.DIODE(\wfg_stim_sine_top.inc_val_q[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13814__A (.DIODE(\wfg_stim_sine_top.inc_val_q[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19595__A1 (.DIODE(\wfg_stim_sine_top.inc_val_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19104__B2 (.DIODE(\wfg_stim_sine_top.inc_val_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13842__A (.DIODE(\wfg_stim_sine_top.inc_val_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13813__A (.DIODE(\wfg_stim_sine_top.inc_val_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19619__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19065__B2 (.DIODE(\wfg_stim_sine_top.offset_val_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17354__A (.DIODE(\wfg_stim_sine_top.offset_val_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17254__A (.DIODE(\wfg_stim_sine_top.offset_val_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19650__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19108__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17273__A (.DIODE(\wfg_stim_sine_top.offset_val_q[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17246__A (.DIODE(\wfg_stim_sine_top.offset_val_q[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19654__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19112__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17310__A (.DIODE(\wfg_stim_sine_top.offset_val_q[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17276__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17275__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19657__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19115__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17277__A (.DIODE(\wfg_stim_sine_top.offset_val_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17245__A (.DIODE(\wfg_stim_sine_top.offset_val_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19660__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19117__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17302__A (.DIODE(\wfg_stim_sine_top.offset_val_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17280__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17279__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19663__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19120__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17281__A (.DIODE(\wfg_stim_sine_top.offset_val_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17244__A (.DIODE(\wfg_stim_sine_top.offset_val_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19666__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19124__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17294__A (.DIODE(\wfg_stim_sine_top.offset_val_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17284__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17283__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19669__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19126__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17285__A (.DIODE(\wfg_stim_sine_top.offset_val_q[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17243__A (.DIODE(\wfg_stim_sine_top.offset_val_q[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19672__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19128__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17070__A (.DIODE(\wfg_stim_sine_top.offset_val_q[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17068__A (.DIODE(\wfg_stim_sine_top.offset_val_q[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19626__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19083__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17257__A (.DIODE(\wfg_stim_sine_top.offset_val_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17252__A (.DIODE(\wfg_stim_sine_top.offset_val_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19629__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19087__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17342__A (.DIODE(\wfg_stim_sine_top.offset_val_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17260__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17259__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19632__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19089__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17261__A (.DIODE(\wfg_stim_sine_top.offset_val_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17251__A (.DIODE(\wfg_stim_sine_top.offset_val_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19635__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19092__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17263__A (.DIODE(\wfg_stim_sine_top.offset_val_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17250__A (.DIODE(\wfg_stim_sine_top.offset_val_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19638__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19096__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17265__A (.DIODE(\wfg_stim_sine_top.offset_val_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17249__A (.DIODE(\wfg_stim_sine_top.offset_val_q[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19641__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19098__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17267__A (.DIODE(\wfg_stim_sine_top.offset_val_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17248__A (.DIODE(\wfg_stim_sine_top.offset_val_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19644__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19102__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17269__A (.DIODE(\wfg_stim_sine_top.offset_val_q[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17247__A (.DIODE(\wfg_stim_sine_top.offset_val_q[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19647__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19104__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17318__A (.DIODE(\wfg_stim_sine_top.offset_val_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17272__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17271__A1 (.DIODE(\wfg_stim_sine_top.offset_val_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19088__A1 (.DIODE(\wfg_stim_sine_top.wbs_dat_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17971__A1 (.DIODE(\wfg_stim_sine_top.wbs_dat_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19094__A1 (.DIODE(\wfg_stim_sine_top.wbs_dat_o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17979__A1 (.DIODE(\wfg_stim_sine_top.wbs_dat_o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17240__B1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.cur_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17232__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.cur_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17157__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.cur_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17154__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.cur_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16599__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.cur_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16462__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.cur_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16454__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.cur_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16432__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.cur_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13918__C (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.cur_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13855__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.cur_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17240__A2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.cur_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17232__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.cur_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17157__C_N (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.cur_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17154__C_N (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.cur_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16431__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.cur_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16428__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.cur_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13918__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.cur_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13855__A_N (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.cur_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17240__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.cur_state[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17232__C_N (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.cur_state[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17157__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.cur_state[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17154__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.cur_state[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16431__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.cur_state[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16428__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.cur_state[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13918__A_N (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.cur_state[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13855__C (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.cur_state[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16895__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.iteration[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16885__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.iteration[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16682__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.iteration[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16499__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.iteration[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16488__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.iteration[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16476__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.iteration[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16446__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.iteration[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16439__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.iteration[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17228__S (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.quadrant[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17176__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.quadrant[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17170__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.quadrant[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17162__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.quadrant[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17161__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.quadrant[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17152__S (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.quadrant[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17113__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.quadrant[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16465__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.quadrant[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17205__B1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.quadrant[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17197__B1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.quadrant[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17189__B1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.quadrant[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17181__B1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.quadrant[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17170__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.quadrant[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17162__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.quadrant[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17161__B1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.quadrant[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17150__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.quadrant[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17113__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.quadrant[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16463__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.quadrant[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16012__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15917__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15916__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15060__D (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14491__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15717__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15658__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15640__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15083__A2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15082__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14685__D (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13931__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15684__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15640__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15608__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15028__A2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14823__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14729__B1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14728__D (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14685__C (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13929__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15660__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15608__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15603__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14823__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14729__A2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14728__C (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14558__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13937__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15615__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15609__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15603__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14558__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13958__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15626__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15617__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15615__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15605__B1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15604__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14447__D (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13956__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15626__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15616__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13968__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15917__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15916__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15875__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15328__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15134__D (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15060__C (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15004__D (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14489__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14486__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15841__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15811__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15316__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15280__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14803__C (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14511__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14498__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14411__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15789__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15779__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15256__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15227__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14818__D (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14530__D (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14266__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15810__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15779__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15738__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15184__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14530__C (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14254__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14252__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13942__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.sin_17[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17070__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.temp[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17068__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.temp[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15601__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.temp[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17228__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17114__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17067__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17065__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16979__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16676__C (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17190__B2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17136__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17040__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17004__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16950__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16670__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16664__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17186__B2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17138__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17037__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17009__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17007__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16670__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16662__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17182__B2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17141__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17034__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16944__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16943__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16672__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16662__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17178__B2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17143__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17032__B2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17011__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16940__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16672__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16657__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17171__A2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17146__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17030__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17014__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16937__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16657__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16653__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17148__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16856__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16653__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16646__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17152__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17024__B1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16808__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16654__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16650__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16648__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16647__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16646__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17226__B2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17115__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17064__B2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16978__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16977__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16688__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16677__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17222__B2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17117__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17062__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16981__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16974__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16688__B2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16675__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17218__B2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17119__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17059__B2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16983__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16971__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16687__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16675__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17214__B2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17121__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17057__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16986__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16968__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16687__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16678__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17210__B2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17123__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17054__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16989__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16965__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16685__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16678__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17206__B2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17126__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17051__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16992__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16962__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16685__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16679__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17202__B2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17128__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17048__B2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16995__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16959__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16679__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16665__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17198__B2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17131__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17046__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16998__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16956__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16669__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16665__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17194__B2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17133__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17043__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17001__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16953__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16669__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16664__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.x[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17190__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17136__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16873__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16867__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16828__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16794__A_N (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16740__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17186__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17138__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16873__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16864__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16825__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16797__A_N (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16737__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17182__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17141__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16875__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16864__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16821__B2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16802__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16800__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17178__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17143__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16875__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16865__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16819__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16731__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16730__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17172__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17146__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16876__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16865__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16817__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16727__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16726__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17165__B2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17148__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16876__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16857__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16815__B2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16805__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16724__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17152__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16898__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16861__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16859__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16858__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16857__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16813__B1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16808__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17214__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17121__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16889__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16879__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16844__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16777__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16758__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17210__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17123__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16892__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16879__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16841__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16779__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16755__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17206__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17126__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16892__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16880__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16838__B2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16782__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16752__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17202__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17128__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16880__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16868__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16836__B2 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16785__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16749__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17198__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17131__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16872__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16868__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16834__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16788__A_N (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16746__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17194__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17133__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16872__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16867__A0 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16831__A1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16791__A_N (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16743__B (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.y[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16975__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.z[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16972__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.z[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16969__B1 (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.z[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16767__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.z[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16764__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.z[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16544__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.z[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16541__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.z[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16467__A (.DIODE(\wfg_stim_sine_top.wfg_stim_sine.z[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19190__B1 (.DIODE(\wfg_subcore_top.active_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18404__A1 (.DIODE(\wfg_subcore_top.active_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18156__A (.DIODE(\wfg_subcore_top.active_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18146__C1 (.DIODE(\wfg_subcore_top.active_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18143__C1 (.DIODE(\wfg_subcore_top.active_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18112__A (.DIODE(\wfg_subcore_top.active_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17411__A (.DIODE(\wfg_subcore_top.active_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17408__B1 (.DIODE(\wfg_subcore_top.active_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17359__A (.DIODE(\wfg_subcore_top.active_o ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19144__A (.DIODE(\wfg_subcore_top.cfg_subcycle_q[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18434__A1 (.DIODE(\wfg_subcore_top.cfg_subcycle_q[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18122__A1 (.DIODE(\wfg_subcore_top.cfg_subcycle_q[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19148__A (.DIODE(\wfg_subcore_top.cfg_subcycle_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18438__A1 (.DIODE(\wfg_subcore_top.cfg_subcycle_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18128__A1 (.DIODE(\wfg_subcore_top.cfg_subcycle_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12515__D (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__12418__D (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__12417__B1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__12384__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__12263__D (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__11610__D (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__11523__B1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__11519__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__11197__D (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__11780__D (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__11611__A2 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__11610__C (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__11183__D (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__11177__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__11780__C (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11201__D (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11179__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11175__D (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__12263__C (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11619__D (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11201__C (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11187__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__12262__A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__12182__C (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11619__C (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11229__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11186__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__12181__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__12178__C (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11311__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11227__C (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11209__D (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11097__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__12065__C (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11209__C (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11091__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11014__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11935__C (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11637__C (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11245__D (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11210__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__10968__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11848__C (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11266__D (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11101__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__10853__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11844__C (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11768__C (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11266__C (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__10703__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__12417__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12361__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12360__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12262__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12261__D (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12182__D (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11383__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11098__C (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__10375__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11094__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__11015__C (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__10374__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__12416__B (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__12360__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__12267__B1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__12266__D (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__12181__B1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__12178__D (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__12103__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__10628__C (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__10368__A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__10362__B (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__B (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10305__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__12425__D (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__12359__B (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__12267__A2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__12266__C (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__12098__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__12065__D (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__12425__C (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__12265__B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__12186__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11934__A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__12426__B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__12355__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__12277__B1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__12275__D (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__12184__B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__12108__C (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__12107__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__11929__A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__11848__D (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__12277__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__12275__C (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11843__A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11768__D (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11939__A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__11767__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__11763__A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__11689__D (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__11772__D (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11687__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11684__D (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11607__D (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11772__C (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11602__A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11524__D (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__18223__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__17945__D (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__17921__D (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__18222__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__17946__D (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__17923__B (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__18222__D (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__17947__C (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__17923__D (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__18222__C (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__17947__B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__17922__C (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__19061__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__18492__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__18487__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__18324__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__18214__B_N (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__19061__A2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__18493__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__18487__B (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__18398__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__18325__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__18214__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__19194__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__19060__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__19028__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__18331__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__18046__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__17933__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__17920__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__17939__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__17932__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__17930__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__18648__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__17950__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__17925__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__19133__B (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__18402__B_N (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__18394__B (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__18333__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__18216__B (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__19191__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__18647__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__18327__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__18287__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__19945__A0 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__19893__A0 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__18237__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__19948__A0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__19897__A0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__18241__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__19951__A0 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__19604__A0 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__18245__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__19954__A0 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__19903__A0 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__18249__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__19957__A0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__19558__A0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__18253__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__19960__A0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__19909__A0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__18257__A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__19809__A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__19669__A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__19155__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__18961__A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__18857__A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__18757__A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__18703__A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__18261__A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__19812__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__19672__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__19157__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__18964__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__18860__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__18706__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__18264__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__19815__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__19161__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__18967__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__18863__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__18710__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__18268__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__19819__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__19163__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__18970__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__18866__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__18713__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__18271__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__19866__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__19838__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__19623__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__19570__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__19518__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__18913__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__18291__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__19822__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__19166__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__18974__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__18870__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__18717__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__18275__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__19825__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__19168__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__18977__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__18873__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__18720__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__18278__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__19829__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__19170__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__18980__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__18876__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__18723__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__18281__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__19832__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__19172__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__18984__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__18879__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__18726__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__18284__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__18987__A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__18882__A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__18729__A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__18990__A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__18887__A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__18732__A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__18993__A0 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__18890__A0 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__18735__A0 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__18996__A0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__18893__A0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__18738__A0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__18999__A0 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__18896__A0 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__18742__A0 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__19002__A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__18899__A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__18745__A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__19920__A0 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__19869__A0 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__19841__A0 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__19626__A0 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__18295__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__19005__A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__18902__A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__18748__A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__19008__A0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__18905__A0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__18751__A0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__19923__A0 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__19872__A0 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__19844__A0 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__19629__A0 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__18299__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__19926__A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__19875__A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__19847__A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__19632__A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__18303__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__19929__A0 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__19878__A0 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__19850__A0 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__19635__A0 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__18307__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__19933__A0 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__19881__A0 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__19853__A0 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__18312__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__19936__A0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__19884__A0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__19856__A0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__18316__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__19939__A0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__19783__A0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__18212__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__19942__A0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__19890__A0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__18232__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__19727__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__19346__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__18585__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__18166__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__18163__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__18217__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__19133__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__18402__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__18394__A_N (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__18216__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__13767__A0 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__13660__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__19779__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__17916__B2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_output122_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_output123_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_output124_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_output126_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_output127_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_output128_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_output135_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_output138_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_output139_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_output140_A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_output141_A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_output142_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_output143_A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_output144_A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_output145_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__17658__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_output146_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__17651__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_output147_A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__17644__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_output148_A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__17633__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_output149_A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__17626__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_output150_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__17619__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_output151_A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__17612__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_output152_A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__17605__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_output153_A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__17597__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_output154_A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__17590__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_output155_A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__17721__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_output156_A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__17583__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_output157_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__17576__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_output158_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__17569__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_output159_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__17558__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_output160_A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__17551__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_output161_A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__17544__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_output162_A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__17537__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_output163_A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__17530__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_output164_A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__17522__A1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_output165_A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__17515__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_output166_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__17714__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_output167_A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__17508__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_output168_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__17501__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_output169_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__17707__A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_output170_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__17700__A1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_output171_A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__17693__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_output172_A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__17686__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_output173_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__17679__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_output174_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__17672__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_output175_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__17665__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_output176_A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__17494__A1 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_output177_A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_output178_A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_output179_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__20462__CLK (.DIODE(clknet_leaf_12_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20512__CLK (.DIODE(clknet_leaf_12_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20511__CLK (.DIODE(clknet_leaf_12_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20458__CLK (.DIODE(clknet_leaf_12_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20457__CLK (.DIODE(clknet_leaf_12_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20510__CLK (.DIODE(clknet_leaf_12_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20509__CLK (.DIODE(clknet_leaf_12_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20444__CLK (.DIODE(clknet_leaf_12_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20498__CLK (.DIODE(clknet_leaf_12_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20497__CLK (.DIODE(clknet_leaf_12_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20442__CLK (.DIODE(clknet_leaf_12_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20443__CLK (.DIODE(clknet_leaf_12_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20375__CLK (.DIODE(clknet_leaf_41_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20383__CLK (.DIODE(clknet_leaf_41_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20407__CLK (.DIODE(clknet_leaf_41_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20327__CLK (.DIODE(clknet_leaf_41_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20408__CLK (.DIODE(clknet_leaf_41_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20310__CLK (.DIODE(clknet_leaf_41_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20571__CLK (.DIODE(clknet_leaf_41_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20588__CLK (.DIODE(clknet_leaf_41_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20306__CLK (.DIODE(clknet_leaf_41_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20360__CLK (.DIODE(clknet_leaf_41_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20376__CLK (.DIODE(clknet_leaf_41_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20367__CLK (.DIODE(clknet_leaf_41_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20225__CLK (.DIODE(clknet_leaf_61_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20224__CLK (.DIODE(clknet_leaf_61_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20222__CLK (.DIODE(clknet_leaf_61_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20943__CLK (.DIODE(clknet_leaf_61_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20944__CLK (.DIODE(clknet_leaf_61_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20234__CLK (.DIODE(clknet_leaf_61_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20227__CLK (.DIODE(clknet_leaf_61_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20235__CLK (.DIODE(clknet_leaf_61_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20236__CLK (.DIODE(clknet_leaf_61_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20284__CLK (.DIODE(clknet_leaf_61_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20508__CLK (.DIODE(clknet_leaf_88_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20505__CLK (.DIODE(clknet_leaf_88_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20271__CLK (.DIODE(clknet_leaf_88_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20265__CLK (.DIODE(clknet_leaf_88_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20504__CLK (.DIODE(clknet_leaf_88_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20501__CLK (.DIODE(clknet_leaf_88_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20502__CLK (.DIODE(clknet_leaf_88_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20446__CLK (.DIODE(clknet_leaf_88_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20503__CLK (.DIODE(clknet_leaf_88_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20448__CLK (.DIODE(clknet_leaf_88_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20552__CLK (.DIODE(clknet_leaf_88_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20298__CLK (.DIODE(clknet_leaf_90_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20261__CLK (.DIODE(clknet_leaf_90_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20251__CLK (.DIODE(clknet_leaf_90_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20495__CLK (.DIODE(clknet_leaf_90_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20496__CLK (.DIODE(clknet_leaf_90_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20500__CLK (.DIODE(clknet_leaf_90_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20445__CLK (.DIODE(clknet_leaf_90_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20499__CLK (.DIODE(clknet_leaf_90_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20268__CLK (.DIODE(clknet_leaf_90_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20266__CLK (.DIODE(clknet_leaf_90_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20262__CLK (.DIODE(clknet_leaf_90_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20263__CLK (.DIODE(clknet_leaf_90_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1_0_io_wbs_clk_A (.DIODE(clknet_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0_0_io_wbs_clk_A (.DIODE(clknet_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1_0_io_wbs_clk_A (.DIODE(clknet_1_0_1_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0_0_io_wbs_clk_A (.DIODE(clknet_1_0_1_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3_0_io_wbs_clk_A (.DIODE(clknet_1_1_1_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2_0_io_wbs_clk_A (.DIODE(clknet_1_1_1_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1_0_io_wbs_clk_A (.DIODE(clknet_2_0_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0_0_io_wbs_clk_A (.DIODE(clknet_2_0_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3_0_io_wbs_clk_A (.DIODE(clknet_2_1_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2_0_io_wbs_clk_A (.DIODE(clknet_2_1_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5_0_io_wbs_clk_A (.DIODE(clknet_2_2_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4_0_io_wbs_clk_A (.DIODE(clknet_2_2_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7_0_io_wbs_clk_A (.DIODE(clknet_2_3_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6_0_io_wbs_clk_A (.DIODE(clknet_2_3_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_109_io_wbs_clk_A (.DIODE(clknet_3_0_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_108_io_wbs_clk_A (.DIODE(clknet_3_0_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_107_io_wbs_clk_A (.DIODE(clknet_3_0_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_106_io_wbs_clk_A (.DIODE(clknet_3_0_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_105_io_wbs_clk_A (.DIODE(clknet_3_0_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_104_io_wbs_clk_A (.DIODE(clknet_3_0_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_103_io_wbs_clk_A (.DIODE(clknet_3_0_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_102_io_wbs_clk_A (.DIODE(clknet_3_0_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_io_wbs_clk_A (.DIODE(clknet_3_0_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_opt_1_0_io_wbs_clk_A (.DIODE(clknet_3_0_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_io_wbs_clk_A (.DIODE(clknet_3_0_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_io_wbs_clk_A (.DIODE(clknet_3_0_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_io_wbs_clk_A (.DIODE(clknet_3_0_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_io_wbs_clk_A (.DIODE(clknet_3_0_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_io_wbs_clk_A (.DIODE(clknet_3_0_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_101_io_wbs_clk_A (.DIODE(clknet_3_1_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_100_io_wbs_clk_A (.DIODE(clknet_3_1_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_99_io_wbs_clk_A (.DIODE(clknet_3_1_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_98_io_wbs_clk_A (.DIODE(clknet_3_1_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_97_io_wbs_clk_A (.DIODE(clknet_3_1_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_96_io_wbs_clk_A (.DIODE(clknet_3_1_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_95_io_wbs_clk_A (.DIODE(clknet_3_1_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_94_io_wbs_clk_A (.DIODE(clknet_3_1_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_93_io_wbs_clk_A (.DIODE(clknet_3_1_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_92_io_wbs_clk_A (.DIODE(clknet_3_1_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_91_io_wbs_clk_A (.DIODE(clknet_3_1_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_90_io_wbs_clk_A (.DIODE(clknet_3_1_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_89_io_wbs_clk_A (.DIODE(clknet_3_1_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_88_io_wbs_clk_A (.DIODE(clknet_3_1_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_84_io_wbs_clk_A (.DIODE(clknet_3_1_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_81_io_wbs_clk_A (.DIODE(clknet_3_1_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_79_io_wbs_clk_A (.DIODE(clknet_3_1_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_io_wbs_clk_A (.DIODE(clknet_3_1_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__20845__CLK (.DIODE(clknet_3_2_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_io_wbs_clk_A (.DIODE(clknet_3_2_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_io_wbs_clk_A (.DIODE(clknet_3_2_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_io_wbs_clk_A (.DIODE(clknet_3_2_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_io_wbs_clk_A (.DIODE(clknet_3_2_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_io_wbs_clk_A (.DIODE(clknet_3_2_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_io_wbs_clk_A (.DIODE(clknet_3_2_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_io_wbs_clk_A (.DIODE(clknet_3_2_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_io_wbs_clk_A (.DIODE(clknet_3_2_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_io_wbs_clk_A (.DIODE(clknet_3_2_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_io_wbs_clk_A (.DIODE(clknet_3_2_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_io_wbs_clk_A (.DIODE(clknet_3_2_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_io_wbs_clk_A (.DIODE(clknet_3_2_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_io_wbs_clk_A (.DIODE(clknet_3_2_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_opt_2_0_io_wbs_clk_A (.DIODE(clknet_3_2_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_87_io_wbs_clk_A (.DIODE(clknet_3_3_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_86_io_wbs_clk_A (.DIODE(clknet_3_3_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_io_wbs_clk_A (.DIODE(clknet_3_3_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_io_wbs_clk_A (.DIODE(clknet_3_3_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_io_wbs_clk_A (.DIODE(clknet_3_3_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_io_wbs_clk_A (.DIODE(clknet_3_3_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_io_wbs_clk_A (.DIODE(clknet_3_3_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_io_wbs_clk_A (.DIODE(clknet_3_3_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_io_wbs_clk_A (.DIODE(clknet_3_3_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_io_wbs_clk_A (.DIODE(clknet_3_3_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_io_wbs_clk_A (.DIODE(clknet_3_3_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_io_wbs_clk_A (.DIODE(clknet_3_3_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_io_wbs_clk_A (.DIODE(clknet_3_3_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_io_wbs_clk_A (.DIODE(clknet_3_4_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_io_wbs_clk_A (.DIODE(clknet_3_4_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_io_wbs_clk_A (.DIODE(clknet_3_4_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_io_wbs_clk_A (.DIODE(clknet_3_4_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_io_wbs_clk_A (.DIODE(clknet_3_4_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_io_wbs_clk_A (.DIODE(clknet_3_4_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_io_wbs_clk_A (.DIODE(clknet_3_4_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_io_wbs_clk_A (.DIODE(clknet_3_4_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_io_wbs_clk_A (.DIODE(clknet_3_4_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_io_wbs_clk_A (.DIODE(clknet_3_4_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_85_io_wbs_clk_A (.DIODE(clknet_3_5_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_83_io_wbs_clk_A (.DIODE(clknet_3_5_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_82_io_wbs_clk_A (.DIODE(clknet_3_5_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_80_io_wbs_clk_A (.DIODE(clknet_3_5_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_opt_3_0_io_wbs_clk_A (.DIODE(clknet_3_5_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_77_io_wbs_clk_A (.DIODE(clknet_3_5_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_76_io_wbs_clk_A (.DIODE(clknet_3_5_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_75_io_wbs_clk_A (.DIODE(clknet_3_5_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_74_io_wbs_clk_A (.DIODE(clknet_3_5_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_73_io_wbs_clk_A (.DIODE(clknet_3_5_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_72_io_wbs_clk_A (.DIODE(clknet_3_5_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_71_io_wbs_clk_A (.DIODE(clknet_3_6_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_70_io_wbs_clk_A (.DIODE(clknet_3_6_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_69_io_wbs_clk_A (.DIODE(clknet_3_6_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_52_io_wbs_clk_A (.DIODE(clknet_3_6_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_io_wbs_clk_A (.DIODE(clknet_3_6_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_io_wbs_clk_A (.DIODE(clknet_3_6_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_io_wbs_clk_A (.DIODE(clknet_3_6_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_io_wbs_clk_A (.DIODE(clknet_3_6_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_io_wbs_clk_A (.DIODE(clknet_3_6_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_io_wbs_clk_A (.DIODE(clknet_3_6_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_io_wbs_clk_A (.DIODE(clknet_3_6_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_io_wbs_clk_A (.DIODE(clknet_3_6_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_68_io_wbs_clk_A (.DIODE(clknet_3_7_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_67_io_wbs_clk_A (.DIODE(clknet_3_7_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_66_io_wbs_clk_A (.DIODE(clknet_3_7_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_65_io_wbs_clk_A (.DIODE(clknet_3_7_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_64_io_wbs_clk_A (.DIODE(clknet_3_7_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_63_io_wbs_clk_A (.DIODE(clknet_3_7_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_62_io_wbs_clk_A (.DIODE(clknet_3_7_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_61_io_wbs_clk_A (.DIODE(clknet_3_7_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_60_io_wbs_clk_A (.DIODE(clknet_3_7_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_59_io_wbs_clk_A (.DIODE(clknet_3_7_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_58_io_wbs_clk_A (.DIODE(clknet_3_7_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_opt_4_0_io_wbs_clk_A (.DIODE(clknet_3_7_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_io_wbs_clk_A (.DIODE(clknet_3_7_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_io_wbs_clk_A (.DIODE(clknet_3_7_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_io_wbs_clk_A (.DIODE(clknet_3_7_0_io_wbs_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_53_io_wbs_clk_A (.DIODE(clknet_3_7_0_io_wbs_clk));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1534 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1094 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1210 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1247 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1253 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1286 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1295 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1302 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1311 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1317 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1325 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1351 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1363 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1413 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1433 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1441 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1446 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1471 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1495 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1511 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1531 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1543 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1555 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_891 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1194 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1227 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1283 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1294 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1305 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1327 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1338 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1344 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1350 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1361 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1382 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1392 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1405 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1424 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1483 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1490 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1496 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1508 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1520 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1528 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1535 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1162 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1260 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1282 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1299 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1305 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1323 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1326 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1332 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1341 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1359 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1375 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1380 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1386 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1419 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1426 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1432 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1271 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1313 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1323 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1326 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1384 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1396 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1405 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1416 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1429 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1447 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1461 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1473 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1103 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1159 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1207 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1248 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1264 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1320 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1411 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1418 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1430 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1436 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1442 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1493 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1505 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1522 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1534 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1546 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1558 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1566 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1282 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1449 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1460 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1472 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1497 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1509 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1524 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1534 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1304 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1314 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1323 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1378 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1425 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1437 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1452 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1466 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1470 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1478 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1488 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1494 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1506 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1523 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1530 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1536 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1548 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1560 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_898 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1299 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1308 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1336 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1389 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1400 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1408 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1420 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1444 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1456 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1462 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1466 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1478 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1491 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1505 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1515 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1526 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1538 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1211 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1263 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1303 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1311 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1322 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1330 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1338 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1366 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1372 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1375 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1387 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1406 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1418 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1437 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1448 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1482 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1489 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1501 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1509 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1518 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1530 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1542 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1554 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1566 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1163 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1251 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1286 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1292 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1298 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1322 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1334 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1348 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1440 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1446 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1458 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1470 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1482 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1485 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1497 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1503 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1507 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1515 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1526 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1532 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1263 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1322 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1330 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1379 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1425 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1437 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1511 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1524 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1532 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1544 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1556 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1066 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1176 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1251 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1278 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1296 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1308 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1325 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1373 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1395 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1407 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1427 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1441 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1450 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1458 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1467 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1474 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1494 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1506 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1514 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1517 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1524 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1530 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1538 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1597 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1148 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1263 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1376 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1415 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1421 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1428 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1457 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1478 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1490 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1502 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1510 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1513 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1531 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1547 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1559 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1601 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1247 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1371 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1383 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1394 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1402 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1405 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1411 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1422 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1440 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1452 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1464 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1468 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1480 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1496 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1508 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1520 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1532 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1538 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1550 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1562 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1574 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1586 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1594 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1304 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1316 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1327 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1376 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1399 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1410 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1438 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1450 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1468 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1479 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1487 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1496 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1503 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1513 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1534 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1546 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1558 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1566 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1271 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1283 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1291 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1337 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1355 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1370 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1391 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1403 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1407 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1410 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1419 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1481 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1505 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1517 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1532 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1541 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1553 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1559 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1563 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1575 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1587 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1114 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1223 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1263 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1358 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1389 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1413 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1425 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1433 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1437 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1443 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1479 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1487 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1490 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1496 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1502 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1510 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1513 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1521 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1535 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1547 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1555 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1564 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1574 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1586 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1598 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1602 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1168 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1238 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1277 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1283 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1295 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1391 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1405 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1417 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1423 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1438 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1451 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1463 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1468 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1474 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1478 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1494 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1498 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1512 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1522 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1541 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1553 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1572 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1583 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1298 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1318 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1369 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1389 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1413 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1425 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1433 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1439 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1455 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1457 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1465 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1470 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1477 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1486 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1496 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1511 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1517 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1529 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1601 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1291 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1311 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1322 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1338 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1350 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1358 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1394 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1404 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1448 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1460 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1468 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1472 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1478 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1493 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1499 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1505 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1517 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1529 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1537 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1557 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1593 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1085 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1263 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1296 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1302 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1314 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1326 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1333 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1338 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1365 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1378 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1421 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1424 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1434 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1457 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1474 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1491 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1503 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1513 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1525 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1558 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1566 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1601 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1153 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1191 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1275 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1281 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1294 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1303 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1405 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1416 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1422 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1450 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1462 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1470 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1500 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1506 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1525 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1535 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1539 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1550 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1562 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1572 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1584 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1153 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1247 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1270 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1298 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1307 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1319 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1387 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1394 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1413 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1421 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1432 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1472 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1489 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1495 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1502 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1513 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1525 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1531 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1543 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1555 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1566 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1575 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1589 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1601 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1182 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1271 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1290 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1298 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1365 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1383 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1395 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1407 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1427 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1437 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1452 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1464 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1472 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1476 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1489 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1495 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1501 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1511 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1523 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1531 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1538 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1550 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1561 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1572 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1085 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1199 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1220 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1226 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1266 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1278 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1293 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1357 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1385 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1394 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1425 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1431 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1438 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1448 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1481 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1501 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1567 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1578 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1588 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1600 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1046 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1185 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1218 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1246 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1335 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1342 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1358 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1361 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1398 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1410 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1444 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1456 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1460 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1466 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1475 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1479 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1494 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1506 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1514 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1528 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_975 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1271 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1285 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1295 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1312 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1324 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1332 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1372 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1389 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1413 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1430 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1442 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1454 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1461 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1467 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1474 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1478 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1486 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1496 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1504 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1522 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1534 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1546 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1558 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1566 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1575 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1582 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1594 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1602 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1183 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1227 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1271 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1326 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1352 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1364 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1390 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1402 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1410 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1434 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1462 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1468 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1472 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1516 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1528 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1538 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1550 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1561 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1569 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1585 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1593 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1087 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1151 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1223 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1275 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1355 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1367 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1379 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1399 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1417 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1453 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1463 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1466 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1474 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1486 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1498 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1510 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1525 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1537 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1545 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1553 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1564 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1599 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1195 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1235 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1291 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1350 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1389 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1411 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1420 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1435 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1483 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1496 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1508 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1516 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1521 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1532 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1559 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1571 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1594 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1154 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1250 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1272 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1305 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1342 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1377 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1383 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1391 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1399 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1407 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1414 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1433 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1450 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1472 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1480 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1491 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1504 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1567 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1573 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1577 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1587 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1599 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1179 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1221 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1227 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1315 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1324 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1334 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1346 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1350 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1380 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1388 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1391 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1402 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1414 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1426 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1446 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1455 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1461 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1465 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1480 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1494 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1506 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1516 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1528 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1534 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1264 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1279 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1313 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1319 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1333 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1340 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1363 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1386 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1394 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1407 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1411 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1417 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1429 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1433 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1439 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1447 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1487 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1493 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1505 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1510 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1523 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1529 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1540 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1555 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1585 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_842 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1134 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1221 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1306 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1312 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1330 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1348 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1360 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1364 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1378 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1393 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1407 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1427 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1437 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1440 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1464 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1476 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1485 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1497 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1502 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1508 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1519 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1528 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1534 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1558 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1566 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1570 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1580 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1590 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_982 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1254 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1260 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1266 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1293 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1304 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1334 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1369 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1381 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1408 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1420 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1432 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1442 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1493 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1505 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1510 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1513 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1519 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1527 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1533 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1551 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1563 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1567 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1579 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1590 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1602 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1059 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1079 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1222 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1254 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1270 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1286 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1295 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1327 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1379 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1382 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1394 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1406 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1412 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1441 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1451 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1461 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1473 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1481 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1485 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1502 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1516 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1526 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1553 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1561 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1583 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1597 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1206 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1248 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1254 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1264 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1315 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1331 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1361 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1368 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1374 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1388 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1405 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1411 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1420 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1432 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1438 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1441 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1454 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1461 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1481 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1493 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1502 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1510 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1513 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1525 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1531 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1567 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1578 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1587 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1599 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1215 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1226 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1270 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1307 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1327 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1339 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1361 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1377 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1389 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1397 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1437 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1447 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1459 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1471 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1505 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1517 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1529 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1538 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1546 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1558 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1566 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1573 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1585 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1593 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1223 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1252 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1296 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1304 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1314 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1320 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1326 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1332 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1357 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1365 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1413 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1428 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1444 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1455 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1457 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1465 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1471 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1483 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1490 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1499 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1503 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1513 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1525 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1531 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1538 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1546 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1558 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1566 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1601 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1269 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1281 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1303 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1330 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1338 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1348 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1360 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1393 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1405 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1413 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1424 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1449 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1464 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1482 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1489 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1521 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1533 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1538 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1545 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1552 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1563 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1575 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1587 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1243 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1355 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1367 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1374 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1413 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1425 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1438 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1468 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1481 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1495 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1511 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1522 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1534 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1542 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1548 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1552 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1557 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1565 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1575 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1582 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1594 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1602 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1296 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1302 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1310 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1368 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1389 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1411 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1427 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1450 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1462 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1470 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1473 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1479 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1483 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1489 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1501 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1504 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1510 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1517 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1523 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1535 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1539 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1545 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1549 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1564 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1572 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1582 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1594 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_927 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1206 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1242 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1255 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1318 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1322 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1326 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1333 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1351 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1363 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1413 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1425 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1432 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1453 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1470 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1474 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1493 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1508 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1528 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1540 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1546 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1552 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1564 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1601 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1188 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1198 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1270 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1280 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1288 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1294 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1307 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1310 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1323 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1332 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1347 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1358 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1368 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1389 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1395 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1406 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1426 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1433 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1450 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1464 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1479 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1497 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1501 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1504 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1530 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1538 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1556 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1568 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1576 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1585 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1594 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1039 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1051 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1108 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1148 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1199 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1256 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1264 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1282 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1308 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1324 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1336 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1342 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1360 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1372 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1384 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1410 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1416 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1428 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1436 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1444 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1448 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1462 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1468 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1478 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1491 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1503 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1525 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1546 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1558 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1566 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1601 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1209 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1215 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1223 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1271 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1283 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1311 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1336 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1344 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1360 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1385 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1400 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1406 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1416 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1429 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1437 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1446 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1454 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1462 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1468 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1476 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1503 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1515 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1519 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1526 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1537 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1547 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1551 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1558 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1577 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1584 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1592 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1255 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1286 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1305 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1319 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1343 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1362 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1382 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1388 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1398 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1455 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1466 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1472 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1480 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1492 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1496 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1551 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1563 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1588 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1600 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1104 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1181 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1209 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1281 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1307 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1333 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1385 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1397 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1403 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1411 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1417 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1465 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1489 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1501 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1509 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1512 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1538 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1549 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1561 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1573 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1586 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1594 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1597 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_926 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1082 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1194 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1206 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1298 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1308 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1314 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1318 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1324 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1354 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1378 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1423 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1432 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1444 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1462 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1470 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1476 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1488 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1500 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1519 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1525 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1536 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1546 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1558 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1566 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1569 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1577 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1585 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_954 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1169 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1198 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1239 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1299 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1333 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1347 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1397 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1422 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1433 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1444 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1456 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1459 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1466 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1478 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1497 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1509 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1519 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1531 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1538 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1565 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1577 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1581 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1585 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1591 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1154 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1260 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1287 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1309 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1321 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1341 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1355 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1367 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1379 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1387 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1396 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1405 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1413 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1432 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1445 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1455 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1465 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1474 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1486 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1498 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1513 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1529 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1565 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1583 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1592 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1600 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1221 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1247 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1281 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1298 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1306 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1312 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1340 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1350 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1354 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1370 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1373 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1387 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1404 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1411 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1417 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1425 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1434 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1440 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1464 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1476 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1494 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1506 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1516 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1522 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1525 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1535 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1561 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1567 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1576 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1585 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1592 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1597 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_926 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1088 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1204 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1311 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1323 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1335 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1361 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1370 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1376 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1384 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1392 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1406 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1418 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1430 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1442 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1450 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1454 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1464 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1471 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1488 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1499 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1511 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1522 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1529 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1537 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1543 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1567 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1584 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1592 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1600 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1294 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1298 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1303 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1344 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1356 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1382 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1400 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1412 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1441 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1452 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1460 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1475 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1483 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1492 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1500 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1511 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1539 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1552 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1564 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1572 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1579 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1586 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1594 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1168 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1286 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1302 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1352 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1399 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1415 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1439 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1455 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1463 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1476 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1488 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1496 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1503 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1511 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1521 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1527 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1533 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1543 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1557 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1566 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1577 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1584 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1596 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1602 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1224 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1247 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1335 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1395 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1406 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1410 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1418 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1441 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1445 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1452 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1458 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1470 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1482 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1485 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1497 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1503 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1507 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1519 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1531 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1539 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1547 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1551 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1563 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1571 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1593 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1307 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1323 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1351 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1369 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1375 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1393 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1407 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1414 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1423 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1430 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1442 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1455 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1462 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1473 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1493 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1501 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1509 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1526 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1534 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1547 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1558 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1564 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1569 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1576 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1582 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1587 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1222 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1234 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1247 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1275 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1281 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1304 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1326 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1338 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1341 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1347 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1362 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1368 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1391 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1403 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1412 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1429 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1433 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1448 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1458 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1471 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1482 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1497 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1509 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1515 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1525 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1531 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1539 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1547 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1560 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1576 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1587 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1593 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1218 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1260 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1266 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1278 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1284 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1309 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1328 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1342 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1367 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1383 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1389 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1395 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1398 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1410 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1417 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1423 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1443 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1450 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1461 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1469 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1473 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1479 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1497 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1504 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1549 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1561 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1564 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1575 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1580 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1588 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1600 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1220 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1247 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1306 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1327 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1331 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1334 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1340 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1346 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1363 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1397 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1407 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1420 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1433 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1445 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1521 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1536 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1548 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1560 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1572 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1580 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1592 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1206 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1228 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1244 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1282 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1303 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1309 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1332 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1338 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1361 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1375 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1387 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1392 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1398 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1414 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1455 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1465 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1477 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1486 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1494 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1506 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1522 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1528 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1540 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1552 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1564 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1575 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1582 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1592 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1600 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1010 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1284 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1314 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1360 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1378 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1386 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1390 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1400 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1408 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1411 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1441 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1447 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1453 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1463 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1474 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1492 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1499 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1505 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1517 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1526 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1536 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1548 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1560 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1564 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1572 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1578 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1585 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1593 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1183 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1279 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1323 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1327 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1378 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1382 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1394 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1412 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1424 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1432 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1439 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1447 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1454 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1461 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1473 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1489 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1496 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1504 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1513 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1525 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1529 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1536 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1548 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1556 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1566 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1580 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1590 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1602 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1209 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1278 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1291 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1314 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1325 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1334 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1346 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1370 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1387 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1399 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1407 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1417 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1425 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1448 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1460 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1472 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1490 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1503 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1515 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1532 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1538 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1546 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1553 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1557 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1575 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1583 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1590 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1215 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1266 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1299 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1323 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1367 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1378 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1388 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1394 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1425 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1438 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1447 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1481 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1490 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1509 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1513 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1522 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1535 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1542 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1552 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1558 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1564 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1573 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1195 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1347 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1390 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1396 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1408 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1420 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1438 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1448 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1455 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1471 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1483 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1489 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1492 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1500 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1506 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1529 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1547 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1550 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1556 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1562 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1568 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1574 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1593 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1260 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1307 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1324 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1332 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1354 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1366 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1374 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1390 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1396 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1416 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1428 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1434 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1439 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1453 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1467 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1477 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1487 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1497 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1503 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1532 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1538 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1544 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1550 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1559 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1565 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1573 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1579 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1585 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1270 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1280 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1304 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1327 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1333 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1344 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1361 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1367 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1389 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1399 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1402 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1408 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1414 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1420 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1426 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1435 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1443 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1455 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1463 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1473 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1485 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1497 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1503 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1506 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1516 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1522 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1528 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1534 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1554 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1566 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1573 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1579 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1585 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1591 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1038 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1134 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1206 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1223 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1263 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1312 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1323 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1335 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1349 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1352 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1360 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1366 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1372 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1386 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1392 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1398 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1405 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1412 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1422 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1428 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1443 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1455 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1461 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1476 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1488 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1492 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1495 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1501 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1511 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1526 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1532 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1538 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1544 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1555 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1559 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1565 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1582 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1594 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1602 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1135 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1224 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1238 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1250 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1281 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1287 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1307 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1326 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1336 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1342 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1348 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1382 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1420 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1433 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1439 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1447 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1453 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1459 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1483 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1489 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1495 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1505 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1511 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1519 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1525 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1538 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1550 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1554 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1561 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1568 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1574 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1580 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1592 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1597 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_972 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1194 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1220 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1255 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1263 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1275 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1299 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1311 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1319 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1331 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1363 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1391 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1405 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1411 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1417 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1428 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1434 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1440 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1454 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1467 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1486 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1493 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1501 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1513 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1517 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1531 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1539 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1547 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1560 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1566 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1569 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1578 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1584 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1588 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1600 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_886 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1113 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1179 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1268 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1284 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1292 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1298 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1304 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1327 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1330 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1352 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1358 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1364 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1387 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1393 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1413 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1420 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1426 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1429 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1443 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1449 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1452 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1466 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1472 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1490 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1508 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1514 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1520 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1526 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1532 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1538 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1557 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1563 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1569 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1581 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1185 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1220 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1247 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1271 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1298 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1308 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1314 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1320 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1326 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1359 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1365 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1383 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1398 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1405 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1408 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1412 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1420 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1426 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1432 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1438 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1446 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1455 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1463 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1470 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1482 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1490 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1496 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1500 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1503 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1518 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1524 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1538 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1544 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1556 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1562 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1113 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1305 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1334 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1338 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1342 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1361 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1379 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1383 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1392 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1400 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1406 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1419 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1425 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1433 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1437 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1441 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1447 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1454 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1465 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1474 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1478 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1489 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1495 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1501 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1511 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1517 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1523 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1529 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1535 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1539 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1552 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1561 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1568 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1580 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1584 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1588 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1215 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1260 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1286 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1306 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1312 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1318 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1326 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1354 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1360 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1366 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1372 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1378 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1392 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1419 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1430 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1436 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1442 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1448 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1454 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1466 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1472 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1476 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1479 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1491 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1497 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1505 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1520 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1529 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1535 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1549 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1558 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1566 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1573 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1591 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1281 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1284 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1290 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1296 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1303 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1315 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1331 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1340 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1344 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1360 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1378 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1390 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1396 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1408 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1416 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1433 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1439 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1451 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1460 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1466 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1479 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1483 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1485 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1489 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1497 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1510 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1522 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1539 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1545 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1551 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1563 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1575 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1579 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1584 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1168 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1220 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1294 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1305 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1312 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1318 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1324 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1332 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1335 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1366 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1383 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1389 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1415 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1433 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1465 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1468 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1474 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1483 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1494 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1500 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1506 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1522 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1548 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1559 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1567 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1577 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1585 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1282 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1294 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1311 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1337 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1347 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1397 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1415 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1433 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1447 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1460 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1472 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1497 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1503 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1513 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1519 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1525 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1531 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1539 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1549 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1552 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1564 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1576 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1584 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1591 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1094 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1332 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1354 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1362 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1380 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1386 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1415 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1422 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1426 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1431 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1438 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1444 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1455 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1461 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1470 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1489 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1501 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1509 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1522 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1534 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1546 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1558 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1562 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1566 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1573 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1577 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1587 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1023 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1270 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1282 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1290 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1295 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1317 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1350 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1378 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1396 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1400 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1404 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1416 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1438 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1446 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1451 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1463 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1475 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1509 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1521 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1529 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1554 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1562 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1571 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1583 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1312 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1324 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1410 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1417 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1439 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1455 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1463 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1467 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1479 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1489 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1501 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1509 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1522 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1531 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1543 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1555 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1561 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1566 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1577 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1589 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1601 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1083 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1299 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1314 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1331 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1366 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1382 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1394 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1406 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1418 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1444 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1456 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1468 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1480 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1489 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1496 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1503 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1515 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1537 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1549 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1561 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1573 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1584 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1143 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1242 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1271 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1287 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1295 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1313 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1325 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1357 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1365 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1374 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1384 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1392 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1417 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1455 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1461 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1473 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1478 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1486 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1494 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1501 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1509 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1513 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1528 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1540 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1550 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1562 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1566 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1573 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1591 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1187 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1246 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1284 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1296 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1302 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1346 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1358 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1383 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1395 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1407 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1436 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1442 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1454 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1462 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1468 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1472 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1479 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1497 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1515 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1527 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1539 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1549 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1553 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1573 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1585 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1593 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1197 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1253 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1284 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1311 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1326 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1369 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1389 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1419 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1439 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1454 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1466 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1472 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1484 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1496 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1504 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1521 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1528 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1534 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1546 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1558 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1566 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1573 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1601 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1003 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1068 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1128 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1268 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1292 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1337 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1350 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1417 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1441 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1456 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1472 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1492 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1504 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1508 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1511 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1522 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1531 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1549 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1562 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1573 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1580 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1592 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_751 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1095 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1253 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1310 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1399 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1406 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1410 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1418 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1436 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1448 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1463 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1480 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1491 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1503 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1523 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1532 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1544 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1556 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1582 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1594 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1602 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_891 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1257 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1284 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1296 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1302 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1373 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1390 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1400 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1412 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1419 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1425 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1436 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1442 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1450 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1459 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1468 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1480 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1491 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1511 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1517 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1523 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1553 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1565 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1571 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1579 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1590 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1597 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_914 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1314 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1326 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1330 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1358 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1362 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1365 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1374 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1380 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1384 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1388 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1408 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1414 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1431 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1438 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1453 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1465 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1488 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1496 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1508 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1525 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1529 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1533 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1540 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1549 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1556 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1575 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1580 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1587 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1599 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1003 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1127 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1180 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1258 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1294 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1326 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1338 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1361 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1379 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1389 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1399 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1411 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1419 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1426 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1440 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1483 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1491 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1498 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1504 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1516 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1519 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1528 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1535 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1539 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1548 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1555 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1561 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1573 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1585 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1593 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1263 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1313 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1319 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1326 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1335 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1352 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1364 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1376 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1425 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1431 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1435 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1483 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1492 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1501 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1513 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1525 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1530 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1536 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1540 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1546 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1552 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1562 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1578 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1590 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1602 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1290 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1317 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1347 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1378 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1402 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1411 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1427 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1435 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1448 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1460 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1472 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1490 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1499 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1505 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1517 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1526 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1539 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1547 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1553 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1559 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1573 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1584 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1016 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1167 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1253 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1268 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1279 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1305 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1312 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1323 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1327 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1350 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1362 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1374 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1386 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1398 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1412 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1436 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1448 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1467 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1479 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1487 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1491 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1500 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1508 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1513 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1525 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1531 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1543 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1555 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1560 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1589 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1601 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_952 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1179 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1284 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1296 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1324 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1393 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1397 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1408 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1417 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1449 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1497 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1501 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1504 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1516 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1530 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1537 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1548 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1554 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1566 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1578 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1590 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1597 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1160 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1207 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1219 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1287 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1340 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1397 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1413 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1423 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1433 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1444 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1465 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1474 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1486 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1501 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1513 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1525 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1536 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1545 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1553 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1560 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1589 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1192 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1236 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1271 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1279 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1284 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1306 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1312 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1325 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1349 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1405 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1414 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1422 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1440 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1449 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1456 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1465 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1474 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1482 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1493 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1501 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1505 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1523 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1535 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1538 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1552 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1561 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1571 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1586 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1594 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1163 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1199 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1286 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1294 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1302 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1308 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1312 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1318 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1343 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1378 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1390 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1396 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1408 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1416 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1422 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1436 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1447 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1455 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1461 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1466 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1499 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1510 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1523 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1531 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1543 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1546 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1554 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1562 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1576 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1583 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1082 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1156 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1247 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1280 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1292 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1305 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1314 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1330 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1336 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1350 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1363 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1385 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1407 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1427 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1439 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1447 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1459 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1471 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1541 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1553 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1559 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1566 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1572 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1582 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1336 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1362 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1374 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1385 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1394 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1401 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1418 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1436 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1448 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1461 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1466 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1478 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1486 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1489 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1500 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1519 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1531 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1543 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1548 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1559 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1567 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1569 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1576 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1586 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1598 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1602 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1292 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1348 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1360 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1397 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1409 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1422 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1438 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1446 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1450 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1462 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1468 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1476 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1497 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1505 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1508 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1519 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1531 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1539 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1541 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1549 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1556 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1092 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1104 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1112 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1252 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1307 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1310 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1399 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1418 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1428 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1442 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1481 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1497 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1567 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1575 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1587 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1599 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1200 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1292 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1314 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1330 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1336 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1348 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1354 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1405 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1418 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1425 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1433 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1444 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1456 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1468 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1495 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1519 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1526 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1534 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1553 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1561 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1568 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1579 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1585 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1593 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1226 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1264 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1299 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1320 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1332 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1396 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1407 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1421 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1427 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1436 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1442 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1457 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1465 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1497 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1505 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1520 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1524 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1531 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1543 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1555 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1566 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1577 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1589 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1601 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1128 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1179 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1236 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1277 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1291 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1348 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1397 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1405 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1408 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1414 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1418 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1441 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1451 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1467 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1473 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1480 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1497 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1509 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1517 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1526 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1538 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1553 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1557 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1563 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1574 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1220 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1264 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1282 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1296 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1316 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1336 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1358 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1368 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1374 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1380 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1392 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1405 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1417 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1422 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1434 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1442 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1447 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1454 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1464 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1509 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1518 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1531 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1543 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1555 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1567 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1578 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1589 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1188 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1333 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1349 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1369 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1393 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1406 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1426 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1439 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1446 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1455 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1464 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1473 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1497 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1501 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1505 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1511 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1517 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1523 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1535 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_960 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1135 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1206 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1246 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1260 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1279 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1311 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1323 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1361 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1368 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1376 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1379 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1431 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1443 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1454 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1466 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1475 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1483 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1495 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1498 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1525 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1529 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1533 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1545 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1557 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1565 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1584 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1596 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1602 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_972 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1028 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1067 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1254 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1278 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1321 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1327 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1339 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1342 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1348 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1351 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1360 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1392 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1441 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1453 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1461 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1479 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1485 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1497 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1506 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1516 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1530 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1538 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1548 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1560 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1570 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1582 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1594 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1597 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1167 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1250 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1262 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1276 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1287 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1320 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1331 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1343 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1354 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1360 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1378 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1390 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1396 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1413 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1423 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1435 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1447 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1478 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1490 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1494 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1504 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1513 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1521 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1531 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1542 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1546 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1553 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1559 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1566 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1577 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1589 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1268 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1291 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1327 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1333 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1344 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1368 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1383 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1395 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1400 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1406 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1419 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1436 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1442 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1454 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1462 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1470 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1480 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1497 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1500 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1511 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1523 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1531 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1535 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1553 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1557 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1572 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1584 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1237 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1254 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1263 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1322 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1334 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1338 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1363 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1376 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1383 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1395 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1423 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1436 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1442 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1477 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1487 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1495 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1500 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1506 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1533 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1545 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1557 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1601 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_843 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1120 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1176 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1280 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1292 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1298 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1301 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1337 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1342 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1357 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1366 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1391 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1403 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1433 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1445 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1322 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1361 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1393 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1408 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1417 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1430 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1442 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1008 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1171 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1243 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1291 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1307 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1322 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1335 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1347 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1355 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1378 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1384 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1396 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1408 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1434 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1446 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1458 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1470 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1482 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1163 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1242 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1262 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1305 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1308 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1319 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1330 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1342 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1362 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1384 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1398 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1401 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1428 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1440 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1601 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1142 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1176 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1242 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1280 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1291 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1298 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1327 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1335 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1370 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1393 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1411 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1156 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1199 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1255 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1307 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1310 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1326 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1338 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1365 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1383 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1601 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_898 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_930 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1283 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1356 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1378 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1384 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1396 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1408 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1420 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1082 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1262 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1266 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1282 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1322 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1367 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1380 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1386 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1392 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1439 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1186 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1292 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1307 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1314 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1323 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1327 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1339 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1363 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1395 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1402 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1434 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1446 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1458 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1470 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1482 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1597 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1083 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1144 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1264 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1305 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1311 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1340 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1412 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1438 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1450 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1194 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1258 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1274 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1296 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1308 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1317 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1331 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1337 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1354 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1361 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1408 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1420 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1597 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_975 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1031 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1151 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1279 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1294 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1306 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1318 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1365 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1377 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1389 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1417 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1433 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1187 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1251 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1296 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1314 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1326 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1333 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1378 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1390 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1401 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1597 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1082 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1163 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1263 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1306 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1310 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1313 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1338 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1350 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1358 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1381 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1389 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1394 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1059 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1211 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1308 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1331 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1356 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1362 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1366 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1392 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1412 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1420 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1424 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1434 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1446 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1458 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1470 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1482 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1597 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_982 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1054 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1096 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1256 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1262 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1312 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1324 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1327 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1333 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1337 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1356 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1362 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1396 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1407 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1431 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1443 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1008 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1254 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1266 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1284 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1290 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1300 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1333 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1340 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1352 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1366 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1395 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1408 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1412 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1419 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1155 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1228 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1254 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1303 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1327 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1368 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1380 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1431 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1443 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1601 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1003 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1059 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1221 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1279 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1282 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1288 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1307 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1322 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1352 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1387 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1411 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1597 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1267 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1286 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1323 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1365 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1375 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1399 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1411 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1423 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1435 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1447 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1601 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1067 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1222 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1247 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1278 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1293 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1332 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1338 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1351 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1368 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1382 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1390 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1394 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1400 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1404 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1434 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1440 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1464 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1476 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1110 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1188 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1206 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1250 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1253 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1266 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1278 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1311 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1320 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1374 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1387 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1408 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1434 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1440 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1601 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1108 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1240 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1270 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1282 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1288 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1298 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1314 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1323 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1344 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1350 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1370 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1393 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1414 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1425 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1434 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1440 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1464 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1476 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1597 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1302 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1312 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1327 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1335 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1376 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1388 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1394 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1408 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1414 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1435 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1447 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1601 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1154 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1290 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1301 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1322 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1336 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1348 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1360 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1387 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1398 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1411 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1422 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1434 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1440 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1464 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1476 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1152 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1167 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1194 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1298 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1322 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1342 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1359 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1376 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1388 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1405 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1411 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1423 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1435 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1447 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_787 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1153 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1279 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1301 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1321 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1327 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1335 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1352 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1371 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1397 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1400 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1413 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1424 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1434 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1440 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1464 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1476 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1188 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1264 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1274 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1301 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1313 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1323 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1342 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1384 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1408 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1412 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1433 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1142 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1211 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1224 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1258 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1284 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1294 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1303 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1326 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1332 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1356 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1393 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1406 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1417 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1434 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1440 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1464 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1476 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1182 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1367 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1391 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1405 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1431 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1443 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1079 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1098 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1292 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1304 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1324 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1330 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1342 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1354 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1360 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1397 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1405 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1597 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_815 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1206 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1221 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1268 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1286 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1298 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1302 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1306 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1601 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1008 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1286 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1347 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1367 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1378 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1404 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1416 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1597 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1212 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1306 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1314 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1319 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1327 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1350 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1358 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1379 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1388 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_955 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1266 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1293 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1322 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1350 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1358 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1380 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1393 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1411 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1199 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1211 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1266 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1294 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1306 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1318 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1330 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1364 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1376 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1382 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1394 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1601 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1286 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1377 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1387 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1395 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1407 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1194 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1319 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1331 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1338 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1350 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1362 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1391 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1406 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1412 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1436 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1448 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1601 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_787 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1285 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1302 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1322 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1330 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1358 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1364 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1399 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1406 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1412 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1038 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1314 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1338 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1367 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_1375 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1406 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1418 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1430 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1442 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1601 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1160 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1180 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1268 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1275 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1291 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1304 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1324 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1331 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1344 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1365 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1387 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1411 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1038 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1244 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1275 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1299 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1361 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1379 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1396 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1601 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1183 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1239 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1247 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1283 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1295 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1597 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1263 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1354 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1360 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1597 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1343 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1361 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1601 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1097 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1597 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1260 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1106 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1168 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1296 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1326 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1350 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1183 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1254 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1269 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_1281 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1299 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1322 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1334 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1338 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1358 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1364 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1377 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1406 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1418 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1430 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1442 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1446 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1601 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_730 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1270 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1290 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1326 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1334 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1340 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1358 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1366 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1383 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1398 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1406 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1412 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1427 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1429 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1437 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1447 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1481 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1500 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1512 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1524 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1536 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1597 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1253 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1265 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1296 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1305 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1323 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1352 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1358 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1365 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1378 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1386 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1410 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1433 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1453 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1466 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1478 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1489 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1500 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1510 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1601 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1067 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1155 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1281 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1332 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1344 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1359 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1366 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1390 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1396 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1402 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1413 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1427 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1437 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1440 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1460 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1472 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1498 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_924 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1298 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1309 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1318 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1362 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1374 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1386 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1405 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1411 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1423 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1435 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1455 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1473 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1496 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1500 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1506 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1601 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1176 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1188 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1281 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1290 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1303 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1403 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1427 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1434 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1445 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1461 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1473 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1481 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1485 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1493 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1505 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1597 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1071 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1098 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1110 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1246 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1264 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1278 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1303 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1353 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1358 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1366 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1379 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1399 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1416 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1423 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1431 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1436 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1443 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1452 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1464 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1471 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1495 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1510 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1601 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1026 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1270 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1283 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1295 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1307 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1310 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1321 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1341 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1380 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1387 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1395 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1403 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1414 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1434 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1440 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1450 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1458 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1464 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1476 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1497 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1501 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1516 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1528 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_982 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1270 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1293 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1306 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1328 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1363 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1378 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1396 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1407 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1413 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1427 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1439 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1447 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1453 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1465 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1477 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1489 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1501 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1533 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1545 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1557 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1130 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1243 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1252 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1275 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1299 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1307 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1324 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1338 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1350 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1393 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1402 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1441 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1470 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1500 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1518 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1530 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1538 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_973 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1248 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1260 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1304 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1312 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1326 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1455 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1464 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1474 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1509 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1518 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1530 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1542 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1554 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1566 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1268 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1280 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1292 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1300 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1405 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1414 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1441 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1462 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1474 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1482 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1508 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1520 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1532 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1039 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1114 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1326 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1338 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1354 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1382 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1394 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1409 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1415 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1428 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1440 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1477 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1485 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1497 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1503 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1528 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1540 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1552 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1564 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1097 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1258 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1274 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1325 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1352 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1378 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1391 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1398 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1406 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1414 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1427 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1439 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1447 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1454 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1460 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1466 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1479 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1527 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1597 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1251 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1271 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1294 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1306 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1312 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1320 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1378 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1398 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1425 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1443 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1455 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1457 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1465 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1477 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1484 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1491 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1503 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1511 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1518 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1530 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1542 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1554 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1566 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1123 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1209 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1280 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1296 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1324 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1331 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1429 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1441 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1447 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1456 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1463 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1479 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1483 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1499 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1505 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_887 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_980 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1260 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1276 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1280 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1298 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1322 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1342 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1351 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1355 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1391 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1394 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1477 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1484 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1488 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1496 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1508 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1067 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1075 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1295 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1303 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1358 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1390 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1410 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1416 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1464 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1476 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1501 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1187 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1254 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1302 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1311 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1318 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1324 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1332 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1335 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1370 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1377 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1389 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1411 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1418 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1424 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1439 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1484 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1496 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1508 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1601 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1288 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1322 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1344 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1356 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1383 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_1395 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1404 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1411 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1465 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_1477 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1491 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1503 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1515 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1527 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1322 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1342 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1353 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1358 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1396 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1425 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1437 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1444 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1482 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1491 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1502 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1179 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1307 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1385 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1410 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1422 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1433 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1441 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1453 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1459 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1470 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1490 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1500 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1507 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1519 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1531 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1084 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1226 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1332 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1358 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1379 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1410 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1420 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1426 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1433 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1442 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1446 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1450 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1457 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1474 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1489 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1501 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1601 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1290 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1314 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1364 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1381 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1408 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1412 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1416 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1438 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1447 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1456 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1468 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1480 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1500 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1512 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1524 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1536 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1286 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1306 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1318 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1330 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1378 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1398 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1411 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1425 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1428 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1440 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1447 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_842 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1122 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1235 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1288 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1389 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1392 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1402 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1426 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1439 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1445 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1210 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1282 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1312 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1324 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1350 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1365 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1379 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1387 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1398 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1412 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1424 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1430 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1438 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1450 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1601 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1225 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1247 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1298 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1310 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1317 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1325 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1332 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1355 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1391 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1403 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1151 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1267 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1294 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1298 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1320 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1326 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1367 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1379 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1601 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1068 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1220 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1275 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1292 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1298 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1323 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1333 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1344 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1355 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1359 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1597 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1087 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1206 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1298 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1304 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1316 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1342 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1351 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1375 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1601 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1256 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1293 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1305 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1350 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1370 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1396 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1401 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1413 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1441 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1449 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1490 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1502 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1510 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1524 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1536 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1541 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1553 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1559 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1569 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1581 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1589 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1594 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1597 ();
 assign io_oeb[0] = net180;
 assign io_oeb[10] = net190;
 assign io_oeb[1] = net181;
 assign io_oeb[2] = net182;
 assign io_oeb[3] = net183;
 assign io_oeb[4] = net184;
 assign io_oeb[5] = net185;
 assign io_oeb[6] = net186;
 assign io_oeb[7] = net187;
 assign io_oeb[8] = net188;
 assign io_oeb[9] = net189;
endmodule

