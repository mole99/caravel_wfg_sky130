// This is the unpowered netlist.
module wb_mux (io_wbs_ack,
    io_wbs_ack_0,
    io_wbs_ack_1,
    io_wbs_cyc,
    io_wbs_cyc_0,
    io_wbs_cyc_1,
    io_wbs_stb,
    io_wbs_stb_0,
    io_wbs_stb_1,
    io_wbs_we,
    io_wbs_we_0,
    io_wbs_we_1,
    io_wbs_adr,
    io_wbs_adr_0,
    io_wbs_adr_1,
    io_wbs_datrd,
    io_wbs_datrd_0,
    io_wbs_datrd_1,
    io_wbs_datwr,
    io_wbs_datwr_0,
    io_wbs_datwr_1,
    io_wbs_sel,
    io_wbs_sel_0,
    io_wbs_sel_1);
 output io_wbs_ack;
 input io_wbs_ack_0;
 input io_wbs_ack_1;
 input io_wbs_cyc;
 output io_wbs_cyc_0;
 output io_wbs_cyc_1;
 input io_wbs_stb;
 output io_wbs_stb_0;
 output io_wbs_stb_1;
 input io_wbs_we;
 output io_wbs_we_0;
 output io_wbs_we_1;
 input [31:0] io_wbs_adr;
 output [31:0] io_wbs_adr_0;
 output [31:0] io_wbs_adr_1;
 output [31:0] io_wbs_datrd;
 input [31:0] io_wbs_datrd_0;
 input [31:0] io_wbs_datrd_1;
 input [31:0] io_wbs_datwr;
 output [31:0] io_wbs_datwr_0;
 output [31:0] io_wbs_datwr_1;
 input [3:0] io_wbs_sel;
 output [3:0] io_wbs_sel_0;
 output [3:0] io_wbs_sel_1;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;

 sky130_fd_sc_hd__or4_1 _021_ (.A(net16),
    .B(net15),
    .C(net18),
    .D(net17),
    .X(_000_));
 sky130_fd_sc_hd__or4bb_1 _022_ (.A(net27),
    .B(net26),
    .C_N(net24),
    .D_N(net23),
    .X(_001_));
 sky130_fd_sc_hd__nor2_1 _023_ (.A(_000_),
    .B(_001_),
    .Y(_002_));
 sky130_fd_sc_hd__or3_1 _024_ (.A(net9),
    .B(net8),
    .C(net7),
    .X(_003_));
 sky130_fd_sc_hd__or4_1 _025_ (.A(net11),
    .B(net10),
    .C(net13),
    .D(net12),
    .X(_004_));
 sky130_fd_sc_hd__or4_1 _026_ (.A(net20),
    .B(net19),
    .C(net22),
    .D(net21),
    .X(_005_));
 sky130_fd_sc_hd__nor3_1 _027_ (.A(_003_),
    .B(_004_),
    .C(_005_),
    .Y(_006_));
 sky130_fd_sc_hd__and3b_1 _028_ (.A_N(net6),
    .B(_002_),
    .C(_006_),
    .X(_007_));
 sky130_fd_sc_hd__buf_2 _029_ (.A(_007_),
    .X(_008_));
 sky130_fd_sc_hd__buf_2 _030_ (.A(_008_),
    .X(_009_));
 sky130_fd_sc_hd__and3_1 _031_ (.A(net6),
    .B(_002_),
    .C(_006_),
    .X(_010_));
 sky130_fd_sc_hd__buf_2 _032_ (.A(_010_),
    .X(_011_));
 sky130_fd_sc_hd__buf_2 _033_ (.A(_011_),
    .X(_012_));
 sky130_fd_sc_hd__a22o_2 _034_ (.A1(net1),
    .A2(_009_),
    .B1(_012_),
    .B2(net2),
    .X(net138));
 sky130_fd_sc_hd__a22o_2 _035_ (.A1(net36),
    .A2(_009_),
    .B1(_012_),
    .B2(net68),
    .X(net205));
 sky130_fd_sc_hd__a22o_2 _036_ (.A1(net47),
    .A2(_009_),
    .B1(_012_),
    .B2(net79),
    .X(net216));
 sky130_fd_sc_hd__a22o_2 _037_ (.A1(net58),
    .A2(_009_),
    .B1(_012_),
    .B2(net90),
    .X(net227));
 sky130_fd_sc_hd__a22o_2 _038_ (.A1(net61),
    .A2(_009_),
    .B1(_012_),
    .B2(net93),
    .X(net230));
 sky130_fd_sc_hd__a22o_2 _039_ (.A1(net62),
    .A2(_009_),
    .B1(_012_),
    .B2(net94),
    .X(net231));
 sky130_fd_sc_hd__a22o_2 _040_ (.A1(net63),
    .A2(_009_),
    .B1(_012_),
    .B2(net95),
    .X(net232));
 sky130_fd_sc_hd__a22o_2 _041_ (.A1(net64),
    .A2(_009_),
    .B1(_012_),
    .B2(net96),
    .X(net233));
 sky130_fd_sc_hd__a22o_2 _042_ (.A1(net65),
    .A2(_009_),
    .B1(_012_),
    .B2(net97),
    .X(net234));
 sky130_fd_sc_hd__a22o_2 _043_ (.A1(net66),
    .A2(_009_),
    .B1(_012_),
    .B2(net98),
    .X(net235));
 sky130_fd_sc_hd__buf_2 _044_ (.A(_008_),
    .X(_013_));
 sky130_fd_sc_hd__buf_2 _045_ (.A(_011_),
    .X(_014_));
 sky130_fd_sc_hd__a22o_2 _046_ (.A1(net67),
    .A2(_013_),
    .B1(_014_),
    .B2(net99),
    .X(net236));
 sky130_fd_sc_hd__a22o_2 _047_ (.A1(net37),
    .A2(_013_),
    .B1(_014_),
    .B2(net69),
    .X(net206));
 sky130_fd_sc_hd__a22o_2 _048_ (.A1(net38),
    .A2(_013_),
    .B1(_014_),
    .B2(net70),
    .X(net207));
 sky130_fd_sc_hd__a22o_2 _049_ (.A1(net39),
    .A2(_013_),
    .B1(_014_),
    .B2(net71),
    .X(net208));
 sky130_fd_sc_hd__a22o_2 _050_ (.A1(net40),
    .A2(_013_),
    .B1(_014_),
    .B2(net72),
    .X(net209));
 sky130_fd_sc_hd__a22o_2 _051_ (.A1(net41),
    .A2(_013_),
    .B1(_014_),
    .B2(net73),
    .X(net210));
 sky130_fd_sc_hd__a22o_2 _052_ (.A1(net42),
    .A2(_013_),
    .B1(_014_),
    .B2(net74),
    .X(net211));
 sky130_fd_sc_hd__a22o_2 _053_ (.A1(net43),
    .A2(_013_),
    .B1(_014_),
    .B2(net75),
    .X(net212));
 sky130_fd_sc_hd__a22o_2 _054_ (.A1(net44),
    .A2(_013_),
    .B1(_014_),
    .B2(net76),
    .X(net213));
 sky130_fd_sc_hd__a22o_2 _055_ (.A1(net45),
    .A2(_013_),
    .B1(_014_),
    .B2(net77),
    .X(net214));
 sky130_fd_sc_hd__buf_2 _056_ (.A(_008_),
    .X(_015_));
 sky130_fd_sc_hd__buf_2 _057_ (.A(_011_),
    .X(_016_));
 sky130_fd_sc_hd__a22o_2 _058_ (.A1(net46),
    .A2(_015_),
    .B1(_016_),
    .B2(net78),
    .X(net215));
 sky130_fd_sc_hd__a22o_2 _059_ (.A1(net48),
    .A2(_015_),
    .B1(_016_),
    .B2(net80),
    .X(net217));
 sky130_fd_sc_hd__a22o_2 _060_ (.A1(net49),
    .A2(_015_),
    .B1(_016_),
    .B2(net81),
    .X(net218));
 sky130_fd_sc_hd__a22o_2 _061_ (.A1(net50),
    .A2(_015_),
    .B1(_016_),
    .B2(net82),
    .X(net219));
 sky130_fd_sc_hd__a22o_2 _062_ (.A1(net51),
    .A2(_015_),
    .B1(_016_),
    .B2(net83),
    .X(net220));
 sky130_fd_sc_hd__a22o_2 _063_ (.A1(net52),
    .A2(_015_),
    .B1(_016_),
    .B2(net84),
    .X(net221));
 sky130_fd_sc_hd__a22o_2 _064_ (.A1(net53),
    .A2(_015_),
    .B1(_016_),
    .B2(net85),
    .X(net222));
 sky130_fd_sc_hd__a22o_2 _065_ (.A1(net54),
    .A2(_015_),
    .B1(_016_),
    .B2(net86),
    .X(net223));
 sky130_fd_sc_hd__a22o_2 _066_ (.A1(net55),
    .A2(_015_),
    .B1(_016_),
    .B2(net87),
    .X(net224));
 sky130_fd_sc_hd__a22o_2 _067_ (.A1(net56),
    .A2(_015_),
    .B1(_016_),
    .B2(net88),
    .X(net225));
 sky130_fd_sc_hd__a22o_2 _068_ (.A1(net57),
    .A2(_008_),
    .B1(_011_),
    .B2(net89),
    .X(net226));
 sky130_fd_sc_hd__a22o_2 _069_ (.A1(net59),
    .A2(_008_),
    .B1(_011_),
    .B2(net91),
    .X(net228));
 sky130_fd_sc_hd__a22o_2 _070_ (.A1(net60),
    .A2(_008_),
    .B1(_011_),
    .B2(net92),
    .X(net229));
 sky130_fd_sc_hd__and2_1 _071_ (.A(net136),
    .B(_008_),
    .X(_017_));
 sky130_fd_sc_hd__clkbuf_1 _072_ (.A(_017_),
    .X(net309));
 sky130_fd_sc_hd__and2_1 _073_ (.A(net35),
    .B(_008_),
    .X(_018_));
 sky130_fd_sc_hd__clkbuf_1 _074_ (.A(_018_),
    .X(net203));
 sky130_fd_sc_hd__and2_1 _075_ (.A(net136),
    .B(_011_),
    .X(_019_));
 sky130_fd_sc_hd__buf_2 _076_ (.A(_019_),
    .X(net310));
 sky130_fd_sc_hd__and2_1 _077_ (.A(net35),
    .B(_011_),
    .X(_020_));
 sky130_fd_sc_hd__buf_2 _078_ (.A(_020_),
    .X(net204));
 sky130_fd_sc_hd__buf_2 _079_ (.A(net3),
    .X(net139));
 sky130_fd_sc_hd__buf_2 _080_ (.A(net14),
    .X(net150));
 sky130_fd_sc_hd__buf_2 _081_ (.A(net25),
    .X(net161));
 sky130_fd_sc_hd__buf_2 _082_ (.A(net28),
    .X(net164));
 sky130_fd_sc_hd__buf_2 _083_ (.A(net29),
    .X(net165));
 sky130_fd_sc_hd__buf_2 _084_ (.A(net30),
    .X(net166));
 sky130_fd_sc_hd__buf_2 _085_ (.A(net31),
    .X(net167));
 sky130_fd_sc_hd__buf_2 _086_ (.A(net32),
    .X(net168));
 sky130_fd_sc_hd__buf_2 _087_ (.A(net33),
    .X(net169));
 sky130_fd_sc_hd__buf_2 _088_ (.A(net34),
    .X(net170));
 sky130_fd_sc_hd__buf_2 _089_ (.A(net4),
    .X(net140));
 sky130_fd_sc_hd__buf_2 _090_ (.A(net5),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_2 _091_ (.A(net6),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_2 _092_ (.A(net7),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_2 _093_ (.A(net8),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_2 _094_ (.A(net9),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_2 _095_ (.A(net10),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 _096_ (.A(net11),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_2 _097_ (.A(net12),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_2 _098_ (.A(net13),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_2 _099_ (.A(net15),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_2 _100_ (.A(net16),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_2 _101_ (.A(net17),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_2 _102_ (.A(net18),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_2 _103_ (.A(net19),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_2 _104_ (.A(net20),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_2 _105_ (.A(net21),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_2 _106_ (.A(net22),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_2 _107_ (.A(net23),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_2 _108_ (.A(net24),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_2 _109_ (.A(net26),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_2 _110_ (.A(net27),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 _111_ (.A(net3),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_1 _112_ (.A(net14),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 _113_ (.A(net25),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 _114_ (.A(net28),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_1 _115_ (.A(net29),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_1 _116_ (.A(net30),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_1 _117_ (.A(net31),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_1 _118_ (.A(net32),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_1 _119_ (.A(net33),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_1 _120_ (.A(net34),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 _121_ (.A(net4),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 _122_ (.A(net5),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_1 _123_ (.A(net6),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 _124_ (.A(net7),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 _125_ (.A(net8),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 _126_ (.A(net9),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 _127_ (.A(net10),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 _128_ (.A(net11),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_1 _129_ (.A(net12),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_1 _130_ (.A(net13),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 _131_ (.A(net15),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 _132_ (.A(net16),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 _133_ (.A(net17),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 _134_ (.A(net18),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_1 _135_ (.A(net19),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 _136_ (.A(net20),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_1 _137_ (.A(net21),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_1 _138_ (.A(net22),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_1 _139_ (.A(net23),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_2 _140_ (.A(net24),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_1 _141_ (.A(net26),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_2 _142_ (.A(net27),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_2 _143_ (.A(net100),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_2 _144_ (.A(net111),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_2 _145_ (.A(net122),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_2 _146_ (.A(net125),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_2 _147_ (.A(net126),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_2 _148_ (.A(net127),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_2 _149_ (.A(net128),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_2 _150_ (.A(net129),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_2 _151_ (.A(net130),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_2 _152_ (.A(net131),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_2 _153_ (.A(net101),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_2 _154_ (.A(net102),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_2 _155_ (.A(net103),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_2 _156_ (.A(net104),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_2 _157_ (.A(net105),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_2 _158_ (.A(net106),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_2 _159_ (.A(net107),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_2 _160_ (.A(net108),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_2 _161_ (.A(net109),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_2 _162_ (.A(net110),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_2 _163_ (.A(net112),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_2 _164_ (.A(net113),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_2 _165_ (.A(net114),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_2 _166_ (.A(net115),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_2 _167_ (.A(net116),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_2 _168_ (.A(net117),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_2 _169_ (.A(net118),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_2 _170_ (.A(net119),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_2 _171_ (.A(net120),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_2 _172_ (.A(net121),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_2 _173_ (.A(net123),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_2 _174_ (.A(net124),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_2 _175_ (.A(net100),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_2 _176_ (.A(net111),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_2 _177_ (.A(net122),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_2 _178_ (.A(net125),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_2 _179_ (.A(net126),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_2 _180_ (.A(net127),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_2 _181_ (.A(net128),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_2 _182_ (.A(net129),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_2 _183_ (.A(net130),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_2 _184_ (.A(net131),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_2 _185_ (.A(net101),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_2 _186_ (.A(net102),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_2 _187_ (.A(net103),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_2 _188_ (.A(net104),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_2 _189_ (.A(net105),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_2 _190_ (.A(net106),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_2 _191_ (.A(net107),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_2 _192_ (.A(net108),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_2 _193_ (.A(net109),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_2 _194_ (.A(net110),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_2 _195_ (.A(net112),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_2 _196_ (.A(net113),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_2 _197_ (.A(net114),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_2 _198_ (.A(net115),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_2 _199_ (.A(net116),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_2 _200_ (.A(net117),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_2 _201_ (.A(net118),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_2 _202_ (.A(net119),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_2 _203_ (.A(net120),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_2 _204_ (.A(net121),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_2 _205_ (.A(net123),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_2 _206_ (.A(net124),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_1 _207_ (.A(net132),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_1 _208_ (.A(net133),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_1 _209_ (.A(net134),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_1 _210_ (.A(net135),
    .X(net304));
 sky130_fd_sc_hd__buf_2 _211_ (.A(net132),
    .X(net305));
 sky130_fd_sc_hd__buf_2 _212_ (.A(net133),
    .X(net306));
 sky130_fd_sc_hd__buf_2 _213_ (.A(net134),
    .X(net307));
 sky130_fd_sc_hd__buf_2 _214_ (.A(net135),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_1 _215_ (.A(net137),
    .X(net311));
 sky130_fd_sc_hd__buf_2 _216_ (.A(net137),
    .X(net312));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(io_wbs_ack_0),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input2 (.A(io_wbs_ack_1),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(io_wbs_adr[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(io_wbs_adr[10]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(io_wbs_adr[11]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input6 (.A(io_wbs_adr[12]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(io_wbs_adr[13]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(io_wbs_adr[14]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(io_wbs_adr[15]),
    .X(net9));
 sky130_fd_sc_hd__dlymetal6s2s_1 input10 (.A(io_wbs_adr[16]),
    .X(net10));
 sky130_fd_sc_hd__dlymetal6s2s_1 input11 (.A(io_wbs_adr[17]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(io_wbs_adr[18]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(io_wbs_adr[19]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(io_wbs_adr[1]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(io_wbs_adr[20]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(io_wbs_adr[21]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(io_wbs_adr[22]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(io_wbs_adr[23]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(io_wbs_adr[24]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(io_wbs_adr[25]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(io_wbs_adr[26]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(io_wbs_adr[27]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(io_wbs_adr[28]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(io_wbs_adr[29]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(io_wbs_adr[2]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(io_wbs_adr[30]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(io_wbs_adr[31]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(io_wbs_adr[3]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(io_wbs_adr[4]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(io_wbs_adr[5]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(io_wbs_adr[6]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(io_wbs_adr[7]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(io_wbs_adr[8]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(io_wbs_adr[9]),
    .X(net34));
 sky130_fd_sc_hd__buf_2 input35 (.A(io_wbs_cyc),
    .X(net35));
 sky130_fd_sc_hd__dlymetal6s2s_1 input36 (.A(io_wbs_datrd_0[0]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(io_wbs_datrd_0[10]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(io_wbs_datrd_0[11]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(io_wbs_datrd_0[12]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(io_wbs_datrd_0[13]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(io_wbs_datrd_0[14]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(io_wbs_datrd_0[15]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(io_wbs_datrd_0[16]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(io_wbs_datrd_0[17]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(io_wbs_datrd_0[18]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(io_wbs_datrd_0[19]),
    .X(net46));
 sky130_fd_sc_hd__dlymetal6s2s_1 input47 (.A(io_wbs_datrd_0[1]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(io_wbs_datrd_0[20]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(io_wbs_datrd_0[21]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(io_wbs_datrd_0[22]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(io_wbs_datrd_0[23]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(io_wbs_datrd_0[24]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(io_wbs_datrd_0[25]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(io_wbs_datrd_0[26]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(io_wbs_datrd_0[27]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(io_wbs_datrd_0[28]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(io_wbs_datrd_0[29]),
    .X(net57));
 sky130_fd_sc_hd__dlymetal6s2s_1 input58 (.A(io_wbs_datrd_0[2]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(io_wbs_datrd_0[30]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(io_wbs_datrd_0[31]),
    .X(net60));
 sky130_fd_sc_hd__dlymetal6s2s_1 input61 (.A(io_wbs_datrd_0[3]),
    .X(net61));
 sky130_fd_sc_hd__dlymetal6s2s_1 input62 (.A(io_wbs_datrd_0[4]),
    .X(net62));
 sky130_fd_sc_hd__dlymetal6s2s_1 input63 (.A(io_wbs_datrd_0[5]),
    .X(net63));
 sky130_fd_sc_hd__dlymetal6s2s_1 input64 (.A(io_wbs_datrd_0[6]),
    .X(net64));
 sky130_fd_sc_hd__dlymetal6s2s_1 input65 (.A(io_wbs_datrd_0[7]),
    .X(net65));
 sky130_fd_sc_hd__dlymetal6s2s_1 input66 (.A(io_wbs_datrd_0[8]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(io_wbs_datrd_0[9]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 input68 (.A(io_wbs_datrd_1[0]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 input69 (.A(io_wbs_datrd_1[10]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 input70 (.A(io_wbs_datrd_1[11]),
    .X(net70));
 sky130_fd_sc_hd__buf_2 input71 (.A(io_wbs_datrd_1[12]),
    .X(net71));
 sky130_fd_sc_hd__buf_2 input72 (.A(io_wbs_datrd_1[13]),
    .X(net72));
 sky130_fd_sc_hd__buf_2 input73 (.A(io_wbs_datrd_1[14]),
    .X(net73));
 sky130_fd_sc_hd__buf_2 input74 (.A(io_wbs_datrd_1[15]),
    .X(net74));
 sky130_fd_sc_hd__buf_2 input75 (.A(io_wbs_datrd_1[16]),
    .X(net75));
 sky130_fd_sc_hd__buf_2 input76 (.A(io_wbs_datrd_1[17]),
    .X(net76));
 sky130_fd_sc_hd__buf_2 input77 (.A(io_wbs_datrd_1[18]),
    .X(net77));
 sky130_fd_sc_hd__buf_2 input78 (.A(io_wbs_datrd_1[19]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 input79 (.A(io_wbs_datrd_1[1]),
    .X(net79));
 sky130_fd_sc_hd__buf_2 input80 (.A(io_wbs_datrd_1[20]),
    .X(net80));
 sky130_fd_sc_hd__buf_2 input81 (.A(io_wbs_datrd_1[21]),
    .X(net81));
 sky130_fd_sc_hd__buf_2 input82 (.A(io_wbs_datrd_1[22]),
    .X(net82));
 sky130_fd_sc_hd__buf_2 input83 (.A(io_wbs_datrd_1[23]),
    .X(net83));
 sky130_fd_sc_hd__buf_2 input84 (.A(io_wbs_datrd_1[24]),
    .X(net84));
 sky130_fd_sc_hd__buf_2 input85 (.A(io_wbs_datrd_1[25]),
    .X(net85));
 sky130_fd_sc_hd__buf_2 input86 (.A(io_wbs_datrd_1[26]),
    .X(net86));
 sky130_fd_sc_hd__buf_2 input87 (.A(io_wbs_datrd_1[27]),
    .X(net87));
 sky130_fd_sc_hd__buf_2 input88 (.A(io_wbs_datrd_1[28]),
    .X(net88));
 sky130_fd_sc_hd__buf_2 input89 (.A(io_wbs_datrd_1[29]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 input90 (.A(io_wbs_datrd_1[2]),
    .X(net90));
 sky130_fd_sc_hd__buf_2 input91 (.A(io_wbs_datrd_1[30]),
    .X(net91));
 sky130_fd_sc_hd__buf_2 input92 (.A(io_wbs_datrd_1[31]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_2 input93 (.A(io_wbs_datrd_1[3]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 input94 (.A(io_wbs_datrd_1[4]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 input95 (.A(io_wbs_datrd_1[5]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 input96 (.A(io_wbs_datrd_1[6]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 input97 (.A(io_wbs_datrd_1[7]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 input98 (.A(io_wbs_datrd_1[8]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 input99 (.A(io_wbs_datrd_1[9]),
    .X(net99));
 sky130_fd_sc_hd__dlymetal6s2s_1 input100 (.A(io_wbs_datwr[0]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_2 input101 (.A(io_wbs_datwr[10]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 input102 (.A(io_wbs_datwr[11]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 input103 (.A(io_wbs_datwr[12]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_2 input104 (.A(io_wbs_datwr[13]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 input105 (.A(io_wbs_datwr[14]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 input106 (.A(io_wbs_datwr[15]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 input107 (.A(io_wbs_datwr[16]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_2 input108 (.A(io_wbs_datwr[17]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 input109 (.A(io_wbs_datwr[18]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 input110 (.A(io_wbs_datwr[19]),
    .X(net110));
 sky130_fd_sc_hd__dlymetal6s2s_1 input111 (.A(io_wbs_datwr[1]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_2 input112 (.A(io_wbs_datwr[20]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_2 input113 (.A(io_wbs_datwr[21]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 input114 (.A(io_wbs_datwr[22]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_2 input115 (.A(io_wbs_datwr[23]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_2 input116 (.A(io_wbs_datwr[24]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_2 input117 (.A(io_wbs_datwr[25]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 input118 (.A(io_wbs_datwr[26]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_2 input119 (.A(io_wbs_datwr[27]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_2 input120 (.A(io_wbs_datwr[28]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 input121 (.A(io_wbs_datwr[29]),
    .X(net121));
 sky130_fd_sc_hd__dlymetal6s2s_1 input122 (.A(io_wbs_datwr[2]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 input123 (.A(io_wbs_datwr[30]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 input124 (.A(io_wbs_datwr[31]),
    .X(net124));
 sky130_fd_sc_hd__dlymetal6s2s_1 input125 (.A(io_wbs_datwr[3]),
    .X(net125));
 sky130_fd_sc_hd__dlymetal6s2s_1 input126 (.A(io_wbs_datwr[4]),
    .X(net126));
 sky130_fd_sc_hd__dlymetal6s2s_1 input127 (.A(io_wbs_datwr[5]),
    .X(net127));
 sky130_fd_sc_hd__dlymetal6s2s_1 input128 (.A(io_wbs_datwr[6]),
    .X(net128));
 sky130_fd_sc_hd__dlymetal6s2s_1 input129 (.A(io_wbs_datwr[7]),
    .X(net129));
 sky130_fd_sc_hd__dlymetal6s2s_1 input130 (.A(io_wbs_datwr[8]),
    .X(net130));
 sky130_fd_sc_hd__dlymetal6s2s_1 input131 (.A(io_wbs_datwr[9]),
    .X(net131));
 sky130_fd_sc_hd__buf_2 input132 (.A(io_wbs_sel[0]),
    .X(net132));
 sky130_fd_sc_hd__buf_2 input133 (.A(io_wbs_sel[1]),
    .X(net133));
 sky130_fd_sc_hd__buf_2 input134 (.A(io_wbs_sel[2]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_4 input135 (.A(io_wbs_sel[3]),
    .X(net135));
 sky130_fd_sc_hd__buf_2 input136 (.A(io_wbs_stb),
    .X(net136));
 sky130_fd_sc_hd__buf_2 input137 (.A(io_wbs_we),
    .X(net137));
 sky130_fd_sc_hd__buf_2 output138 (.A(net138),
    .X(io_wbs_ack));
 sky130_fd_sc_hd__buf_2 output139 (.A(net139),
    .X(io_wbs_adr_0[0]));
 sky130_fd_sc_hd__buf_2 output140 (.A(net140),
    .X(io_wbs_adr_0[10]));
 sky130_fd_sc_hd__buf_2 output141 (.A(net141),
    .X(io_wbs_adr_0[11]));
 sky130_fd_sc_hd__buf_2 output142 (.A(net142),
    .X(io_wbs_adr_0[12]));
 sky130_fd_sc_hd__buf_2 output143 (.A(net143),
    .X(io_wbs_adr_0[13]));
 sky130_fd_sc_hd__buf_2 output144 (.A(net144),
    .X(io_wbs_adr_0[14]));
 sky130_fd_sc_hd__buf_2 output145 (.A(net145),
    .X(io_wbs_adr_0[15]));
 sky130_fd_sc_hd__buf_2 output146 (.A(net146),
    .X(io_wbs_adr_0[16]));
 sky130_fd_sc_hd__buf_2 output147 (.A(net147),
    .X(io_wbs_adr_0[17]));
 sky130_fd_sc_hd__buf_2 output148 (.A(net148),
    .X(io_wbs_adr_0[18]));
 sky130_fd_sc_hd__buf_2 output149 (.A(net149),
    .X(io_wbs_adr_0[19]));
 sky130_fd_sc_hd__buf_2 output150 (.A(net150),
    .X(io_wbs_adr_0[1]));
 sky130_fd_sc_hd__buf_2 output151 (.A(net151),
    .X(io_wbs_adr_0[20]));
 sky130_fd_sc_hd__buf_2 output152 (.A(net152),
    .X(io_wbs_adr_0[21]));
 sky130_fd_sc_hd__buf_2 output153 (.A(net153),
    .X(io_wbs_adr_0[22]));
 sky130_fd_sc_hd__buf_2 output154 (.A(net154),
    .X(io_wbs_adr_0[23]));
 sky130_fd_sc_hd__buf_2 output155 (.A(net155),
    .X(io_wbs_adr_0[24]));
 sky130_fd_sc_hd__buf_2 output156 (.A(net156),
    .X(io_wbs_adr_0[25]));
 sky130_fd_sc_hd__buf_2 output157 (.A(net157),
    .X(io_wbs_adr_0[26]));
 sky130_fd_sc_hd__buf_2 output158 (.A(net158),
    .X(io_wbs_adr_0[27]));
 sky130_fd_sc_hd__buf_2 output159 (.A(net159),
    .X(io_wbs_adr_0[28]));
 sky130_fd_sc_hd__buf_2 output160 (.A(net160),
    .X(io_wbs_adr_0[29]));
 sky130_fd_sc_hd__buf_2 output161 (.A(net161),
    .X(io_wbs_adr_0[2]));
 sky130_fd_sc_hd__buf_2 output162 (.A(net162),
    .X(io_wbs_adr_0[30]));
 sky130_fd_sc_hd__buf_2 output163 (.A(net163),
    .X(io_wbs_adr_0[31]));
 sky130_fd_sc_hd__buf_2 output164 (.A(net164),
    .X(io_wbs_adr_0[3]));
 sky130_fd_sc_hd__buf_2 output165 (.A(net165),
    .X(io_wbs_adr_0[4]));
 sky130_fd_sc_hd__buf_2 output166 (.A(net166),
    .X(io_wbs_adr_0[5]));
 sky130_fd_sc_hd__buf_2 output167 (.A(net167),
    .X(io_wbs_adr_0[6]));
 sky130_fd_sc_hd__buf_2 output168 (.A(net168),
    .X(io_wbs_adr_0[7]));
 sky130_fd_sc_hd__buf_2 output169 (.A(net169),
    .X(io_wbs_adr_0[8]));
 sky130_fd_sc_hd__buf_2 output170 (.A(net170),
    .X(io_wbs_adr_0[9]));
 sky130_fd_sc_hd__buf_2 output171 (.A(net171),
    .X(io_wbs_adr_1[0]));
 sky130_fd_sc_hd__buf_2 output172 (.A(net172),
    .X(io_wbs_adr_1[10]));
 sky130_fd_sc_hd__buf_2 output173 (.A(net173),
    .X(io_wbs_adr_1[11]));
 sky130_fd_sc_hd__buf_2 output174 (.A(net174),
    .X(io_wbs_adr_1[12]));
 sky130_fd_sc_hd__buf_2 output175 (.A(net175),
    .X(io_wbs_adr_1[13]));
 sky130_fd_sc_hd__buf_2 output176 (.A(net176),
    .X(io_wbs_adr_1[14]));
 sky130_fd_sc_hd__buf_2 output177 (.A(net177),
    .X(io_wbs_adr_1[15]));
 sky130_fd_sc_hd__buf_2 output178 (.A(net178),
    .X(io_wbs_adr_1[16]));
 sky130_fd_sc_hd__buf_2 output179 (.A(net179),
    .X(io_wbs_adr_1[17]));
 sky130_fd_sc_hd__buf_2 output180 (.A(net180),
    .X(io_wbs_adr_1[18]));
 sky130_fd_sc_hd__buf_2 output181 (.A(net181),
    .X(io_wbs_adr_1[19]));
 sky130_fd_sc_hd__buf_2 output182 (.A(net182),
    .X(io_wbs_adr_1[1]));
 sky130_fd_sc_hd__buf_2 output183 (.A(net183),
    .X(io_wbs_adr_1[20]));
 sky130_fd_sc_hd__buf_2 output184 (.A(net184),
    .X(io_wbs_adr_1[21]));
 sky130_fd_sc_hd__buf_2 output185 (.A(net185),
    .X(io_wbs_adr_1[22]));
 sky130_fd_sc_hd__buf_2 output186 (.A(net186),
    .X(io_wbs_adr_1[23]));
 sky130_fd_sc_hd__buf_2 output187 (.A(net187),
    .X(io_wbs_adr_1[24]));
 sky130_fd_sc_hd__buf_2 output188 (.A(net188),
    .X(io_wbs_adr_1[25]));
 sky130_fd_sc_hd__buf_2 output189 (.A(net189),
    .X(io_wbs_adr_1[26]));
 sky130_fd_sc_hd__buf_2 output190 (.A(net190),
    .X(io_wbs_adr_1[27]));
 sky130_fd_sc_hd__buf_2 output191 (.A(net191),
    .X(io_wbs_adr_1[28]));
 sky130_fd_sc_hd__buf_2 output192 (.A(net192),
    .X(io_wbs_adr_1[29]));
 sky130_fd_sc_hd__buf_2 output193 (.A(net193),
    .X(io_wbs_adr_1[2]));
 sky130_fd_sc_hd__buf_2 output194 (.A(net194),
    .X(io_wbs_adr_1[30]));
 sky130_fd_sc_hd__buf_2 output195 (.A(net195),
    .X(io_wbs_adr_1[31]));
 sky130_fd_sc_hd__buf_2 output196 (.A(net196),
    .X(io_wbs_adr_1[3]));
 sky130_fd_sc_hd__buf_2 output197 (.A(net197),
    .X(io_wbs_adr_1[4]));
 sky130_fd_sc_hd__buf_2 output198 (.A(net198),
    .X(io_wbs_adr_1[5]));
 sky130_fd_sc_hd__buf_2 output199 (.A(net199),
    .X(io_wbs_adr_1[6]));
 sky130_fd_sc_hd__buf_2 output200 (.A(net200),
    .X(io_wbs_adr_1[7]));
 sky130_fd_sc_hd__buf_2 output201 (.A(net201),
    .X(io_wbs_adr_1[8]));
 sky130_fd_sc_hd__buf_2 output202 (.A(net202),
    .X(io_wbs_adr_1[9]));
 sky130_fd_sc_hd__buf_2 output203 (.A(net203),
    .X(io_wbs_cyc_0));
 sky130_fd_sc_hd__buf_2 output204 (.A(net204),
    .X(io_wbs_cyc_1));
 sky130_fd_sc_hd__buf_2 output205 (.A(net205),
    .X(io_wbs_datrd[0]));
 sky130_fd_sc_hd__buf_2 output206 (.A(net206),
    .X(io_wbs_datrd[10]));
 sky130_fd_sc_hd__buf_2 output207 (.A(net207),
    .X(io_wbs_datrd[11]));
 sky130_fd_sc_hd__buf_2 output208 (.A(net208),
    .X(io_wbs_datrd[12]));
 sky130_fd_sc_hd__buf_2 output209 (.A(net209),
    .X(io_wbs_datrd[13]));
 sky130_fd_sc_hd__buf_2 output210 (.A(net210),
    .X(io_wbs_datrd[14]));
 sky130_fd_sc_hd__buf_2 output211 (.A(net211),
    .X(io_wbs_datrd[15]));
 sky130_fd_sc_hd__buf_2 output212 (.A(net212),
    .X(io_wbs_datrd[16]));
 sky130_fd_sc_hd__buf_2 output213 (.A(net213),
    .X(io_wbs_datrd[17]));
 sky130_fd_sc_hd__buf_2 output214 (.A(net214),
    .X(io_wbs_datrd[18]));
 sky130_fd_sc_hd__buf_2 output215 (.A(net215),
    .X(io_wbs_datrd[19]));
 sky130_fd_sc_hd__buf_2 output216 (.A(net216),
    .X(io_wbs_datrd[1]));
 sky130_fd_sc_hd__buf_2 output217 (.A(net217),
    .X(io_wbs_datrd[20]));
 sky130_fd_sc_hd__buf_2 output218 (.A(net218),
    .X(io_wbs_datrd[21]));
 sky130_fd_sc_hd__buf_2 output219 (.A(net219),
    .X(io_wbs_datrd[22]));
 sky130_fd_sc_hd__buf_2 output220 (.A(net220),
    .X(io_wbs_datrd[23]));
 sky130_fd_sc_hd__buf_2 output221 (.A(net221),
    .X(io_wbs_datrd[24]));
 sky130_fd_sc_hd__buf_2 output222 (.A(net222),
    .X(io_wbs_datrd[25]));
 sky130_fd_sc_hd__buf_2 output223 (.A(net223),
    .X(io_wbs_datrd[26]));
 sky130_fd_sc_hd__buf_2 output224 (.A(net224),
    .X(io_wbs_datrd[27]));
 sky130_fd_sc_hd__buf_2 output225 (.A(net225),
    .X(io_wbs_datrd[28]));
 sky130_fd_sc_hd__buf_2 output226 (.A(net226),
    .X(io_wbs_datrd[29]));
 sky130_fd_sc_hd__buf_2 output227 (.A(net227),
    .X(io_wbs_datrd[2]));
 sky130_fd_sc_hd__buf_2 output228 (.A(net228),
    .X(io_wbs_datrd[30]));
 sky130_fd_sc_hd__buf_2 output229 (.A(net229),
    .X(io_wbs_datrd[31]));
 sky130_fd_sc_hd__buf_2 output230 (.A(net230),
    .X(io_wbs_datrd[3]));
 sky130_fd_sc_hd__buf_2 output231 (.A(net231),
    .X(io_wbs_datrd[4]));
 sky130_fd_sc_hd__buf_2 output232 (.A(net232),
    .X(io_wbs_datrd[5]));
 sky130_fd_sc_hd__buf_2 output233 (.A(net233),
    .X(io_wbs_datrd[6]));
 sky130_fd_sc_hd__buf_2 output234 (.A(net234),
    .X(io_wbs_datrd[7]));
 sky130_fd_sc_hd__buf_2 output235 (.A(net235),
    .X(io_wbs_datrd[8]));
 sky130_fd_sc_hd__buf_2 output236 (.A(net236),
    .X(io_wbs_datrd[9]));
 sky130_fd_sc_hd__buf_2 output237 (.A(net237),
    .X(io_wbs_datwr_0[0]));
 sky130_fd_sc_hd__buf_2 output238 (.A(net238),
    .X(io_wbs_datwr_0[10]));
 sky130_fd_sc_hd__buf_2 output239 (.A(net239),
    .X(io_wbs_datwr_0[11]));
 sky130_fd_sc_hd__buf_2 output240 (.A(net240),
    .X(io_wbs_datwr_0[12]));
 sky130_fd_sc_hd__buf_2 output241 (.A(net241),
    .X(io_wbs_datwr_0[13]));
 sky130_fd_sc_hd__buf_2 output242 (.A(net242),
    .X(io_wbs_datwr_0[14]));
 sky130_fd_sc_hd__buf_2 output243 (.A(net243),
    .X(io_wbs_datwr_0[15]));
 sky130_fd_sc_hd__buf_2 output244 (.A(net244),
    .X(io_wbs_datwr_0[16]));
 sky130_fd_sc_hd__buf_2 output245 (.A(net245),
    .X(io_wbs_datwr_0[17]));
 sky130_fd_sc_hd__buf_2 output246 (.A(net246),
    .X(io_wbs_datwr_0[18]));
 sky130_fd_sc_hd__buf_2 output247 (.A(net247),
    .X(io_wbs_datwr_0[19]));
 sky130_fd_sc_hd__buf_2 output248 (.A(net248),
    .X(io_wbs_datwr_0[1]));
 sky130_fd_sc_hd__buf_2 output249 (.A(net249),
    .X(io_wbs_datwr_0[20]));
 sky130_fd_sc_hd__buf_2 output250 (.A(net250),
    .X(io_wbs_datwr_0[21]));
 sky130_fd_sc_hd__buf_2 output251 (.A(net251),
    .X(io_wbs_datwr_0[22]));
 sky130_fd_sc_hd__buf_2 output252 (.A(net252),
    .X(io_wbs_datwr_0[23]));
 sky130_fd_sc_hd__buf_2 output253 (.A(net253),
    .X(io_wbs_datwr_0[24]));
 sky130_fd_sc_hd__buf_2 output254 (.A(net254),
    .X(io_wbs_datwr_0[25]));
 sky130_fd_sc_hd__buf_2 output255 (.A(net255),
    .X(io_wbs_datwr_0[26]));
 sky130_fd_sc_hd__buf_2 output256 (.A(net256),
    .X(io_wbs_datwr_0[27]));
 sky130_fd_sc_hd__buf_2 output257 (.A(net257),
    .X(io_wbs_datwr_0[28]));
 sky130_fd_sc_hd__buf_2 output258 (.A(net258),
    .X(io_wbs_datwr_0[29]));
 sky130_fd_sc_hd__buf_2 output259 (.A(net259),
    .X(io_wbs_datwr_0[2]));
 sky130_fd_sc_hd__buf_2 output260 (.A(net260),
    .X(io_wbs_datwr_0[30]));
 sky130_fd_sc_hd__buf_2 output261 (.A(net261),
    .X(io_wbs_datwr_0[31]));
 sky130_fd_sc_hd__buf_2 output262 (.A(net262),
    .X(io_wbs_datwr_0[3]));
 sky130_fd_sc_hd__buf_2 output263 (.A(net263),
    .X(io_wbs_datwr_0[4]));
 sky130_fd_sc_hd__buf_2 output264 (.A(net264),
    .X(io_wbs_datwr_0[5]));
 sky130_fd_sc_hd__buf_2 output265 (.A(net265),
    .X(io_wbs_datwr_0[6]));
 sky130_fd_sc_hd__buf_2 output266 (.A(net266),
    .X(io_wbs_datwr_0[7]));
 sky130_fd_sc_hd__buf_2 output267 (.A(net267),
    .X(io_wbs_datwr_0[8]));
 sky130_fd_sc_hd__buf_2 output268 (.A(net268),
    .X(io_wbs_datwr_0[9]));
 sky130_fd_sc_hd__buf_2 output269 (.A(net269),
    .X(io_wbs_datwr_1[0]));
 sky130_fd_sc_hd__buf_2 output270 (.A(net270),
    .X(io_wbs_datwr_1[10]));
 sky130_fd_sc_hd__buf_2 output271 (.A(net271),
    .X(io_wbs_datwr_1[11]));
 sky130_fd_sc_hd__buf_2 output272 (.A(net272),
    .X(io_wbs_datwr_1[12]));
 sky130_fd_sc_hd__buf_2 output273 (.A(net273),
    .X(io_wbs_datwr_1[13]));
 sky130_fd_sc_hd__buf_2 output274 (.A(net274),
    .X(io_wbs_datwr_1[14]));
 sky130_fd_sc_hd__buf_2 output275 (.A(net275),
    .X(io_wbs_datwr_1[15]));
 sky130_fd_sc_hd__buf_2 output276 (.A(net276),
    .X(io_wbs_datwr_1[16]));
 sky130_fd_sc_hd__buf_2 output277 (.A(net277),
    .X(io_wbs_datwr_1[17]));
 sky130_fd_sc_hd__buf_2 output278 (.A(net278),
    .X(io_wbs_datwr_1[18]));
 sky130_fd_sc_hd__buf_2 output279 (.A(net279),
    .X(io_wbs_datwr_1[19]));
 sky130_fd_sc_hd__buf_2 output280 (.A(net280),
    .X(io_wbs_datwr_1[1]));
 sky130_fd_sc_hd__buf_2 output281 (.A(net281),
    .X(io_wbs_datwr_1[20]));
 sky130_fd_sc_hd__buf_2 output282 (.A(net282),
    .X(io_wbs_datwr_1[21]));
 sky130_fd_sc_hd__buf_2 output283 (.A(net283),
    .X(io_wbs_datwr_1[22]));
 sky130_fd_sc_hd__buf_2 output284 (.A(net284),
    .X(io_wbs_datwr_1[23]));
 sky130_fd_sc_hd__buf_2 output285 (.A(net285),
    .X(io_wbs_datwr_1[24]));
 sky130_fd_sc_hd__buf_2 output286 (.A(net286),
    .X(io_wbs_datwr_1[25]));
 sky130_fd_sc_hd__buf_2 output287 (.A(net287),
    .X(io_wbs_datwr_1[26]));
 sky130_fd_sc_hd__buf_2 output288 (.A(net288),
    .X(io_wbs_datwr_1[27]));
 sky130_fd_sc_hd__buf_2 output289 (.A(net289),
    .X(io_wbs_datwr_1[28]));
 sky130_fd_sc_hd__buf_2 output290 (.A(net290),
    .X(io_wbs_datwr_1[29]));
 sky130_fd_sc_hd__buf_2 output291 (.A(net291),
    .X(io_wbs_datwr_1[2]));
 sky130_fd_sc_hd__buf_2 output292 (.A(net292),
    .X(io_wbs_datwr_1[30]));
 sky130_fd_sc_hd__buf_2 output293 (.A(net293),
    .X(io_wbs_datwr_1[31]));
 sky130_fd_sc_hd__buf_2 output294 (.A(net294),
    .X(io_wbs_datwr_1[3]));
 sky130_fd_sc_hd__buf_2 output295 (.A(net295),
    .X(io_wbs_datwr_1[4]));
 sky130_fd_sc_hd__buf_2 output296 (.A(net296),
    .X(io_wbs_datwr_1[5]));
 sky130_fd_sc_hd__buf_2 output297 (.A(net297),
    .X(io_wbs_datwr_1[6]));
 sky130_fd_sc_hd__buf_2 output298 (.A(net298),
    .X(io_wbs_datwr_1[7]));
 sky130_fd_sc_hd__buf_2 output299 (.A(net299),
    .X(io_wbs_datwr_1[8]));
 sky130_fd_sc_hd__buf_2 output300 (.A(net300),
    .X(io_wbs_datwr_1[9]));
 sky130_fd_sc_hd__buf_2 output301 (.A(net301),
    .X(io_wbs_sel_0[0]));
 sky130_fd_sc_hd__buf_2 output302 (.A(net302),
    .X(io_wbs_sel_0[1]));
 sky130_fd_sc_hd__buf_2 output303 (.A(net303),
    .X(io_wbs_sel_0[2]));
 sky130_fd_sc_hd__buf_2 output304 (.A(net304),
    .X(io_wbs_sel_0[3]));
 sky130_fd_sc_hd__buf_2 output305 (.A(net305),
    .X(io_wbs_sel_1[0]));
 sky130_fd_sc_hd__buf_2 output306 (.A(net306),
    .X(io_wbs_sel_1[1]));
 sky130_fd_sc_hd__buf_2 output307 (.A(net307),
    .X(io_wbs_sel_1[2]));
 sky130_fd_sc_hd__buf_2 output308 (.A(net308),
    .X(io_wbs_sel_1[3]));
 sky130_fd_sc_hd__buf_2 output309 (.A(net309),
    .X(io_wbs_stb_0));
 sky130_fd_sc_hd__buf_2 output310 (.A(net310),
    .X(io_wbs_stb_1));
 sky130_fd_sc_hd__buf_2 output311 (.A(net311),
    .X(io_wbs_we_0));
 sky130_fd_sc_hd__buf_2 output312 (.A(net312),
    .X(io_wbs_we_1));
 sky130_fd_sc_hd__diode_2 ANTENNA__029__A (.DIODE(_007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__073__B (.DIODE(_008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__071__B (.DIODE(_008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__070__A2 (.DIODE(_008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__069__A2 (.DIODE(_008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__068__A2 (.DIODE(_008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__056__A (.DIODE(_008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__044__A (.DIODE(_008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__030__A (.DIODE(_008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__032__A (.DIODE(_010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__077__B (.DIODE(_011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__075__B (.DIODE(_011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__070__B1 (.DIODE(_011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__069__B1 (.DIODE(_011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__068__B1 (.DIODE(_011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__057__A (.DIODE(_011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__045__A (.DIODE(_011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__033__A (.DIODE(_011_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_wbs_ack_0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(io_wbs_ack_1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(io_wbs_adr[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(io_wbs_adr[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(io_wbs_adr[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(io_wbs_adr[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(io_wbs_adr[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(io_wbs_adr[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(io_wbs_adr[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(io_wbs_adr[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(io_wbs_adr[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(io_wbs_adr[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(io_wbs_adr[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(io_wbs_adr[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(io_wbs_adr[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(io_wbs_adr[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(io_wbs_adr[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(io_wbs_adr[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(io_wbs_adr[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(io_wbs_adr[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(io_wbs_adr[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(io_wbs_adr[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(io_wbs_adr[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(io_wbs_adr[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(io_wbs_adr[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(io_wbs_adr[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(io_wbs_adr[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(io_wbs_adr[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(io_wbs_adr[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(io_wbs_adr[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(io_wbs_adr[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(io_wbs_adr[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(io_wbs_adr[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(io_wbs_adr[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(io_wbs_cyc));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(io_wbs_datrd_0[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(io_wbs_datrd_0[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(io_wbs_datrd_0[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(io_wbs_datrd_0[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(io_wbs_datrd_0[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(io_wbs_datrd_0[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(io_wbs_datrd_0[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(io_wbs_datrd_0[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(io_wbs_datrd_0[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(io_wbs_datrd_0[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(io_wbs_datrd_0[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(io_wbs_datrd_0[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(io_wbs_datrd_0[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(io_wbs_datrd_0[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(io_wbs_datrd_0[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(io_wbs_datrd_0[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(io_wbs_datrd_0[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(io_wbs_datrd_0[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(io_wbs_datrd_0[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(io_wbs_datrd_0[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(io_wbs_datrd_0[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(io_wbs_datrd_0[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(io_wbs_datrd_0[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(io_wbs_datrd_0[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(io_wbs_datrd_0[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(io_wbs_datrd_0[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(io_wbs_datrd_0[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(io_wbs_datrd_0[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(io_wbs_datrd_0[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(io_wbs_datrd_0[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(io_wbs_datrd_0[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(io_wbs_datrd_0[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(io_wbs_datrd_1[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(io_wbs_datrd_1[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(io_wbs_datrd_1[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(io_wbs_datrd_1[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(io_wbs_datrd_1[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(io_wbs_datrd_1[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(io_wbs_datrd_1[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(io_wbs_datrd_1[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(io_wbs_datrd_1[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(io_wbs_datrd_1[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(io_wbs_datrd_1[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(io_wbs_datrd_1[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(io_wbs_datrd_1[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(io_wbs_datrd_1[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(io_wbs_datrd_1[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(io_wbs_datrd_1[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(io_wbs_datrd_1[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(io_wbs_datrd_1[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(io_wbs_datrd_1[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(io_wbs_datrd_1[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(io_wbs_datrd_1[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(io_wbs_datrd_1[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(io_wbs_datrd_1[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(io_wbs_datrd_1[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(io_wbs_datrd_1[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(io_wbs_datrd_1[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(io_wbs_datrd_1[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(io_wbs_datrd_1[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(io_wbs_datrd_1[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(io_wbs_datrd_1[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_A (.DIODE(io_wbs_datrd_1[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_A (.DIODE(io_wbs_datrd_1[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input100_A (.DIODE(io_wbs_datwr[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input101_A (.DIODE(io_wbs_datwr[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input102_A (.DIODE(io_wbs_datwr[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input103_A (.DIODE(io_wbs_datwr[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input104_A (.DIODE(io_wbs_datwr[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input105_A (.DIODE(io_wbs_datwr[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input106_A (.DIODE(io_wbs_datwr[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input107_A (.DIODE(io_wbs_datwr[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input108_A (.DIODE(io_wbs_datwr[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input109_A (.DIODE(io_wbs_datwr[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input110_A (.DIODE(io_wbs_datwr[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input111_A (.DIODE(io_wbs_datwr[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input112_A (.DIODE(io_wbs_datwr[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input113_A (.DIODE(io_wbs_datwr[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input114_A (.DIODE(io_wbs_datwr[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input115_A (.DIODE(io_wbs_datwr[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input116_A (.DIODE(io_wbs_datwr[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input117_A (.DIODE(io_wbs_datwr[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input118_A (.DIODE(io_wbs_datwr[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input119_A (.DIODE(io_wbs_datwr[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input120_A (.DIODE(io_wbs_datwr[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input121_A (.DIODE(io_wbs_datwr[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input122_A (.DIODE(io_wbs_datwr[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input123_A (.DIODE(io_wbs_datwr[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input124_A (.DIODE(io_wbs_datwr[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input125_A (.DIODE(io_wbs_datwr[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input126_A (.DIODE(io_wbs_datwr[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input127_A (.DIODE(io_wbs_datwr[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input128_A (.DIODE(io_wbs_datwr[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input129_A (.DIODE(io_wbs_datwr[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input130_A (.DIODE(io_wbs_datwr[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input131_A (.DIODE(io_wbs_datwr[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input132_A (.DIODE(io_wbs_sel[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input133_A (.DIODE(io_wbs_sel[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input134_A (.DIODE(io_wbs_sel[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input135_A (.DIODE(io_wbs_sel[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input136_A (.DIODE(io_wbs_stb));
 sky130_fd_sc_hd__diode_2 ANTENNA_input137_A (.DIODE(io_wbs_we));
 sky130_fd_sc_hd__diode_2 ANTENNA__034__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__034__B2 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__123__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__091__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__031__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__028__A_N (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__124__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__092__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__024__C (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__125__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__093__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__024__B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__126__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__094__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__024__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__127__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__095__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__025__B (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__128__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__096__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__025__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__129__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__097__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__025__D (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__130__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__098__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__025__C (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__131__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__099__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__021__B (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__132__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__100__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__021__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__133__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__101__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__021__D (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__134__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__102__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__021__C (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__135__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__103__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__026__B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__136__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__104__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__026__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__137__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__105__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__026__D (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__138__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__106__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__026__C (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__139__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__107__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__022__D_N (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__140__A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__108__A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__022__C_N (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__141__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__109__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__022__B (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__142__A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__110__A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__022__A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__077__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__073__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__035__A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__047__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__048__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__049__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__050__A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__051__A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__052__A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__053__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__054__A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__055__A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__036__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__067__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__068__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__037__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__069__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__070__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__038__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__039__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__040__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__041__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__042__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__043__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__046__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__035__B2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__047__B2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__048__B2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__049__B2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__050__B2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__051__B2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__052__B2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__053__B2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__054__B2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__055__B2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__058__B2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__036__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__059__B2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__060__B2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__061__B2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__062__B2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__063__B2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__064__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__065__B2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__066__B2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__067__B2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__068__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__037__B2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__069__B2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__070__B2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__038__B2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__039__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__040__B2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__041__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__042__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__043__B2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__046__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__175__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__143__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__185__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__153__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__186__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__154__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__187__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__155__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__188__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__156__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__189__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__157__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__190__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__158__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__191__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__159__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__192__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__160__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__193__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__161__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__194__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__162__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__176__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__144__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__195__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__163__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__196__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__164__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__197__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__165__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__198__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__166__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__199__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__167__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__200__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__168__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__201__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__169__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__202__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__170__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__203__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__171__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__204__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__172__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__177__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__145__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__205__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__173__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__206__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__174__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__178__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__146__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__179__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__147__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__180__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__148__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__181__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__149__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__182__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__150__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__183__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__151__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__184__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__152__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__211__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__207__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__212__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__208__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__213__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__209__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__214__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__210__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__075__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__071__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__216__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__215__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_output138_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_output139_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_output140_A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_output141_A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_output142_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_output143_A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_output144_A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_output145_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_output146_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_output147_A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_output148_A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_output149_A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_output150_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_output151_A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_output152_A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_output153_A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_output154_A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_output155_A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_output156_A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_output157_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_output158_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_output159_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_output160_A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_output161_A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_output162_A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_output163_A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_output164_A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_output165_A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_output166_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_output167_A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_output168_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_output169_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_output170_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_output189_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_output190_A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_output191_A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_output192_A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_output194_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_output195_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_output203_A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_output204_A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_output205_A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_output206_A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_output207_A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_output208_A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_output209_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_output210_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_output211_A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_output212_A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_output213_A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_output214_A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_output215_A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_output216_A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_output217_A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_output218_A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_output219_A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_output220_A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_output221_A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_output222_A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_output223_A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_output224_A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_output225_A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_output226_A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_output227_A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_output228_A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_output229_A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_output230_A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_output231_A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_output232_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_output233_A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_output234_A (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_output235_A (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_output236_A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_output237_A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_output238_A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_output239_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_output240_A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_output241_A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_output242_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_output243_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_output244_A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_output245_A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_output246_A (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_output247_A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_output248_A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_output249_A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_output250_A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_output251_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_output252_A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_output253_A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_output254_A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_output255_A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_output256_A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_output257_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_output258_A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_output259_A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_output260_A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_output261_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_output262_A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_output263_A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_output264_A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_output265_A (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_output266_A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_output267_A (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_output268_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_output269_A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_output270_A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_output271_A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_output272_A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_output273_A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_output274_A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_output275_A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_output276_A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_output277_A (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_output278_A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_output279_A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_output280_A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_output281_A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_output282_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_output283_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_output284_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_output285_A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_output286_A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_output287_A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_output288_A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_output289_A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_output290_A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_output291_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_output292_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_output293_A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_output294_A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_output295_A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_output296_A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_output297_A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_output298_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_output299_A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_output300_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_output305_A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_output306_A (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_output307_A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_output308_A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_output309_A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_output310_A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_output312_A (.DIODE(net312));
 sky130_fd_sc_hd__decap_6 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_841 ();
endmodule

