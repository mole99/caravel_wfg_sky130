VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_memory
  CLASS BLOCK ;
  FOREIGN wb_memory ;
  ORIGIN 0.000 0.000 ;
  SIZE 750.000 BY 200.000 ;
  PIN addr_mem0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 196.000 22.910 200.000 ;
    END
  END addr_mem0[0]
  PIN addr_mem0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 196.000 41.310 200.000 ;
    END
  END addr_mem0[1]
  PIN addr_mem0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 196.000 59.710 200.000 ;
    END
  END addr_mem0[2]
  PIN addr_mem0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 196.000 78.110 200.000 ;
    END
  END addr_mem0[3]
  PIN addr_mem0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 196.000 96.510 200.000 ;
    END
  END addr_mem0[4]
  PIN addr_mem0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 196.000 110.310 200.000 ;
    END
  END addr_mem0[5]
  PIN addr_mem0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 196.000 124.110 200.000 ;
    END
  END addr_mem0[6]
  PIN addr_mem0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 196.000 137.910 200.000 ;
    END
  END addr_mem0[7]
  PIN addr_mem0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 196.000 151.710 200.000 ;
    END
  END addr_mem0[8]
  PIN addr_mem1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 196.000 386.310 200.000 ;
    END
  END addr_mem1[0]
  PIN addr_mem1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.430 196.000 404.710 200.000 ;
    END
  END addr_mem1[1]
  PIN addr_mem1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 196.000 423.110 200.000 ;
    END
  END addr_mem1[2]
  PIN addr_mem1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 196.000 441.510 200.000 ;
    END
  END addr_mem1[3]
  PIN addr_mem1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.630 196.000 459.910 200.000 ;
    END
  END addr_mem1[4]
  PIN addr_mem1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 196.000 473.710 200.000 ;
    END
  END addr_mem1[5]
  PIN addr_mem1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 196.000 487.510 200.000 ;
    END
  END addr_mem1[6]
  PIN addr_mem1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.030 196.000 501.310 200.000 ;
    END
  END addr_mem1[7]
  PIN addr_mem1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 196.000 515.110 200.000 ;
    END
  END addr_mem1[8]
  PIN csb_mem0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 196.000 13.710 200.000 ;
    END
  END csb_mem0
  PIN csb_mem1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 196.000 377.110 200.000 ;
    END
  END csb_mem1
  PIN din_mem0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 196.000 27.510 200.000 ;
    END
  END din_mem0[0]
  PIN din_mem0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 196.000 174.710 200.000 ;
    END
  END din_mem0[10]
  PIN din_mem0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 196.000 183.910 200.000 ;
    END
  END din_mem0[11]
  PIN din_mem0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 196.000 193.110 200.000 ;
    END
  END din_mem0[12]
  PIN din_mem0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 196.000 202.310 200.000 ;
    END
  END din_mem0[13]
  PIN din_mem0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 196.000 211.510 200.000 ;
    END
  END din_mem0[14]
  PIN din_mem0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 196.000 220.710 200.000 ;
    END
  END din_mem0[15]
  PIN din_mem0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 196.000 229.910 200.000 ;
    END
  END din_mem0[16]
  PIN din_mem0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 196.000 239.110 200.000 ;
    END
  END din_mem0[17]
  PIN din_mem0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 196.000 248.310 200.000 ;
    END
  END din_mem0[18]
  PIN din_mem0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 196.000 257.510 200.000 ;
    END
  END din_mem0[19]
  PIN din_mem0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 196.000 45.910 200.000 ;
    END
  END din_mem0[1]
  PIN din_mem0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 196.000 266.710 200.000 ;
    END
  END din_mem0[20]
  PIN din_mem0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 196.000 275.910 200.000 ;
    END
  END din_mem0[21]
  PIN din_mem0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 196.000 285.110 200.000 ;
    END
  END din_mem0[22]
  PIN din_mem0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 196.000 294.310 200.000 ;
    END
  END din_mem0[23]
  PIN din_mem0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 196.000 303.510 200.000 ;
    END
  END din_mem0[24]
  PIN din_mem0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 196.000 312.710 200.000 ;
    END
  END din_mem0[25]
  PIN din_mem0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 196.000 321.910 200.000 ;
    END
  END din_mem0[26]
  PIN din_mem0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 196.000 331.110 200.000 ;
    END
  END din_mem0[27]
  PIN din_mem0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 196.000 340.310 200.000 ;
    END
  END din_mem0[28]
  PIN din_mem0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 196.000 349.510 200.000 ;
    END
  END din_mem0[29]
  PIN din_mem0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 196.000 64.310 200.000 ;
    END
  END din_mem0[2]
  PIN din_mem0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 196.000 358.710 200.000 ;
    END
  END din_mem0[30]
  PIN din_mem0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 196.000 367.910 200.000 ;
    END
  END din_mem0[31]
  PIN din_mem0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 196.000 82.710 200.000 ;
    END
  END din_mem0[3]
  PIN din_mem0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 196.000 101.110 200.000 ;
    END
  END din_mem0[4]
  PIN din_mem0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 196.000 114.910 200.000 ;
    END
  END din_mem0[5]
  PIN din_mem0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 196.000 128.710 200.000 ;
    END
  END din_mem0[6]
  PIN din_mem0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 196.000 142.510 200.000 ;
    END
  END din_mem0[7]
  PIN din_mem0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 196.000 156.310 200.000 ;
    END
  END din_mem0[8]
  PIN din_mem0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 196.000 165.510 200.000 ;
    END
  END din_mem0[9]
  PIN din_mem1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 196.000 390.910 200.000 ;
    END
  END din_mem1[0]
  PIN din_mem1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 196.000 538.110 200.000 ;
    END
  END din_mem1[10]
  PIN din_mem1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.030 196.000 547.310 200.000 ;
    END
  END din_mem1[11]
  PIN din_mem1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 196.000 556.510 200.000 ;
    END
  END din_mem1[12]
  PIN din_mem1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.430 196.000 565.710 200.000 ;
    END
  END din_mem1[13]
  PIN din_mem1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.630 196.000 574.910 200.000 ;
    END
  END din_mem1[14]
  PIN din_mem1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.830 196.000 584.110 200.000 ;
    END
  END din_mem1[15]
  PIN din_mem1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.030 196.000 593.310 200.000 ;
    END
  END din_mem1[16]
  PIN din_mem1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 196.000 602.510 200.000 ;
    END
  END din_mem1[17]
  PIN din_mem1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.430 196.000 611.710 200.000 ;
    END
  END din_mem1[18]
  PIN din_mem1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.630 196.000 620.910 200.000 ;
    END
  END din_mem1[19]
  PIN din_mem1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 196.000 409.310 200.000 ;
    END
  END din_mem1[1]
  PIN din_mem1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.830 196.000 630.110 200.000 ;
    END
  END din_mem1[20]
  PIN din_mem1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.030 196.000 639.310 200.000 ;
    END
  END din_mem1[21]
  PIN din_mem1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.230 196.000 648.510 200.000 ;
    END
  END din_mem1[22]
  PIN din_mem1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.430 196.000 657.710 200.000 ;
    END
  END din_mem1[23]
  PIN din_mem1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 196.000 666.910 200.000 ;
    END
  END din_mem1[24]
  PIN din_mem1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.830 196.000 676.110 200.000 ;
    END
  END din_mem1[25]
  PIN din_mem1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 196.000 685.310 200.000 ;
    END
  END din_mem1[26]
  PIN din_mem1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 196.000 694.510 200.000 ;
    END
  END din_mem1[27]
  PIN din_mem1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.430 196.000 703.710 200.000 ;
    END
  END din_mem1[28]
  PIN din_mem1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.630 196.000 712.910 200.000 ;
    END
  END din_mem1[29]
  PIN din_mem1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 196.000 427.710 200.000 ;
    END
  END din_mem1[2]
  PIN din_mem1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.830 196.000 722.110 200.000 ;
    END
  END din_mem1[30]
  PIN din_mem1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 196.000 731.310 200.000 ;
    END
  END din_mem1[31]
  PIN din_mem1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 196.000 446.110 200.000 ;
    END
  END din_mem1[3]
  PIN din_mem1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.230 196.000 464.510 200.000 ;
    END
  END din_mem1[4]
  PIN din_mem1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.030 196.000 478.310 200.000 ;
    END
  END din_mem1[5]
  PIN din_mem1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.830 196.000 492.110 200.000 ;
    END
  END din_mem1[6]
  PIN din_mem1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 196.000 505.910 200.000 ;
    END
  END din_mem1[7]
  PIN din_mem1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 196.000 519.710 200.000 ;
    END
  END din_mem1[8]
  PIN din_mem1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.630 196.000 528.910 200.000 ;
    END
  END din_mem1[9]
  PIN dout_mem0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 196.000 32.110 200.000 ;
    END
  END dout_mem0[0]
  PIN dout_mem0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 196.000 179.310 200.000 ;
    END
  END dout_mem0[10]
  PIN dout_mem0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 196.000 188.510 200.000 ;
    END
  END dout_mem0[11]
  PIN dout_mem0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 196.000 197.710 200.000 ;
    END
  END dout_mem0[12]
  PIN dout_mem0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 196.000 206.910 200.000 ;
    END
  END dout_mem0[13]
  PIN dout_mem0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 196.000 216.110 200.000 ;
    END
  END dout_mem0[14]
  PIN dout_mem0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 196.000 225.310 200.000 ;
    END
  END dout_mem0[15]
  PIN dout_mem0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 196.000 234.510 200.000 ;
    END
  END dout_mem0[16]
  PIN dout_mem0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 196.000 243.710 200.000 ;
    END
  END dout_mem0[17]
  PIN dout_mem0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 196.000 252.910 200.000 ;
    END
  END dout_mem0[18]
  PIN dout_mem0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 196.000 262.110 200.000 ;
    END
  END dout_mem0[19]
  PIN dout_mem0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 196.000 50.510 200.000 ;
    END
  END dout_mem0[1]
  PIN dout_mem0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 196.000 271.310 200.000 ;
    END
  END dout_mem0[20]
  PIN dout_mem0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 196.000 280.510 200.000 ;
    END
  END dout_mem0[21]
  PIN dout_mem0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 196.000 289.710 200.000 ;
    END
  END dout_mem0[22]
  PIN dout_mem0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 196.000 298.910 200.000 ;
    END
  END dout_mem0[23]
  PIN dout_mem0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 196.000 308.110 200.000 ;
    END
  END dout_mem0[24]
  PIN dout_mem0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 196.000 317.310 200.000 ;
    END
  END dout_mem0[25]
  PIN dout_mem0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 196.000 326.510 200.000 ;
    END
  END dout_mem0[26]
  PIN dout_mem0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 196.000 335.710 200.000 ;
    END
  END dout_mem0[27]
  PIN dout_mem0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 196.000 344.910 200.000 ;
    END
  END dout_mem0[28]
  PIN dout_mem0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 196.000 354.110 200.000 ;
    END
  END dout_mem0[29]
  PIN dout_mem0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 196.000 68.910 200.000 ;
    END
  END dout_mem0[2]
  PIN dout_mem0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 196.000 363.310 200.000 ;
    END
  END dout_mem0[30]
  PIN dout_mem0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 196.000 372.510 200.000 ;
    END
  END dout_mem0[31]
  PIN dout_mem0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 196.000 87.310 200.000 ;
    END
  END dout_mem0[3]
  PIN dout_mem0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 196.000 105.710 200.000 ;
    END
  END dout_mem0[4]
  PIN dout_mem0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 196.000 119.510 200.000 ;
    END
  END dout_mem0[5]
  PIN dout_mem0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 196.000 133.310 200.000 ;
    END
  END dout_mem0[6]
  PIN dout_mem0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 196.000 147.110 200.000 ;
    END
  END dout_mem0[7]
  PIN dout_mem0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 196.000 160.910 200.000 ;
    END
  END dout_mem0[8]
  PIN dout_mem0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 196.000 170.110 200.000 ;
    END
  END dout_mem0[9]
  PIN dout_mem1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 196.000 395.510 200.000 ;
    END
  END dout_mem1[0]
  PIN dout_mem1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 196.000 542.710 200.000 ;
    END
  END dout_mem1[10]
  PIN dout_mem1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 196.000 551.910 200.000 ;
    END
  END dout_mem1[11]
  PIN dout_mem1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 196.000 561.110 200.000 ;
    END
  END dout_mem1[12]
  PIN dout_mem1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 196.000 570.310 200.000 ;
    END
  END dout_mem1[13]
  PIN dout_mem1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 196.000 579.510 200.000 ;
    END
  END dout_mem1[14]
  PIN dout_mem1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.430 196.000 588.710 200.000 ;
    END
  END dout_mem1[15]
  PIN dout_mem1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 196.000 597.910 200.000 ;
    END
  END dout_mem1[16]
  PIN dout_mem1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.830 196.000 607.110 200.000 ;
    END
  END dout_mem1[17]
  PIN dout_mem1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.030 196.000 616.310 200.000 ;
    END
  END dout_mem1[18]
  PIN dout_mem1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.230 196.000 625.510 200.000 ;
    END
  END dout_mem1[19]
  PIN dout_mem1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 196.000 413.910 200.000 ;
    END
  END dout_mem1[1]
  PIN dout_mem1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 196.000 634.710 200.000 ;
    END
  END dout_mem1[20]
  PIN dout_mem1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.630 196.000 643.910 200.000 ;
    END
  END dout_mem1[21]
  PIN dout_mem1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.830 196.000 653.110 200.000 ;
    END
  END dout_mem1[22]
  PIN dout_mem1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.030 196.000 662.310 200.000 ;
    END
  END dout_mem1[23]
  PIN dout_mem1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.230 196.000 671.510 200.000 ;
    END
  END dout_mem1[24]
  PIN dout_mem1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 196.000 680.710 200.000 ;
    END
  END dout_mem1[25]
  PIN dout_mem1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.630 196.000 689.910 200.000 ;
    END
  END dout_mem1[26]
  PIN dout_mem1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 196.000 699.110 200.000 ;
    END
  END dout_mem1[27]
  PIN dout_mem1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.030 196.000 708.310 200.000 ;
    END
  END dout_mem1[28]
  PIN dout_mem1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.230 196.000 717.510 200.000 ;
    END
  END dout_mem1[29]
  PIN dout_mem1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 196.000 432.310 200.000 ;
    END
  END dout_mem1[2]
  PIN dout_mem1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.430 196.000 726.710 200.000 ;
    END
  END dout_mem1[30]
  PIN dout_mem1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.630 196.000 735.910 200.000 ;
    END
  END dout_mem1[31]
  PIN dout_mem1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.430 196.000 450.710 200.000 ;
    END
  END dout_mem1[3]
  PIN dout_mem1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.830 196.000 469.110 200.000 ;
    END
  END dout_mem1[4]
  PIN dout_mem1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.630 196.000 482.910 200.000 ;
    END
  END dout_mem1[5]
  PIN dout_mem1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 196.000 496.710 200.000 ;
    END
  END dout_mem1[6]
  PIN dout_mem1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.230 196.000 510.510 200.000 ;
    END
  END dout_mem1[7]
  PIN dout_mem1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 196.000 524.310 200.000 ;
    END
  END dout_mem1[8]
  PIN dout_mem1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.230 196.000 533.510 200.000 ;
    END
  END dout_mem1[9]
  PIN io_wbs_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 4.000 ;
    END
  END io_wbs_ack
  PIN io_wbs_adr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END io_wbs_adr[0]
  PIN io_wbs_adr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END io_wbs_adr[10]
  PIN io_wbs_adr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END io_wbs_adr[11]
  PIN io_wbs_adr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 0.000 330.190 4.000 ;
    END
  END io_wbs_adr[12]
  PIN io_wbs_adr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END io_wbs_adr[13]
  PIN io_wbs_adr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 0.000 371.590 4.000 ;
    END
  END io_wbs_adr[14]
  PIN io_wbs_adr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END io_wbs_adr[15]
  PIN io_wbs_adr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 0.000 412.990 4.000 ;
    END
  END io_wbs_adr[16]
  PIN io_wbs_adr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 0.000 433.690 4.000 ;
    END
  END io_wbs_adr[17]
  PIN io_wbs_adr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END io_wbs_adr[18]
  PIN io_wbs_adr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.810 0.000 475.090 4.000 ;
    END
  END io_wbs_adr[19]
  PIN io_wbs_adr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 4.000 ;
    END
  END io_wbs_adr[1]
  PIN io_wbs_adr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 0.000 495.790 4.000 ;
    END
  END io_wbs_adr[20]
  PIN io_wbs_adr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 0.000 516.490 4.000 ;
    END
  END io_wbs_adr[21]
  PIN io_wbs_adr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 0.000 537.190 4.000 ;
    END
  END io_wbs_adr[22]
  PIN io_wbs_adr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.610 0.000 557.890 4.000 ;
    END
  END io_wbs_adr[23]
  PIN io_wbs_adr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 0.000 578.590 4.000 ;
    END
  END io_wbs_adr[24]
  PIN io_wbs_adr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END io_wbs_adr[25]
  PIN io_wbs_adr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 0.000 619.990 4.000 ;
    END
  END io_wbs_adr[26]
  PIN io_wbs_adr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.410 0.000 640.690 4.000 ;
    END
  END io_wbs_adr[27]
  PIN io_wbs_adr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.110 0.000 661.390 4.000 ;
    END
  END io_wbs_adr[28]
  PIN io_wbs_adr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.810 0.000 682.090 4.000 ;
    END
  END io_wbs_adr[29]
  PIN io_wbs_adr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END io_wbs_adr[2]
  PIN io_wbs_adr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 0.000 702.790 4.000 ;
    END
  END io_wbs_adr[30]
  PIN io_wbs_adr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.210 0.000 723.490 4.000 ;
    END
  END io_wbs_adr[31]
  PIN io_wbs_adr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END io_wbs_adr[3]
  PIN io_wbs_adr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END io_wbs_adr[4]
  PIN io_wbs_adr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END io_wbs_adr[5]
  PIN io_wbs_adr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END io_wbs_adr[6]
  PIN io_wbs_adr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END io_wbs_adr[7]
  PIN io_wbs_adr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 4.000 ;
    END
  END io_wbs_adr[8]
  PIN io_wbs_adr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 4.000 ;
    END
  END io_wbs_adr[9]
  PIN io_wbs_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END io_wbs_clk
  PIN io_wbs_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END io_wbs_cyc
  PIN io_wbs_datrd[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END io_wbs_datrd[0]
  PIN io_wbs_datrd[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END io_wbs_datrd[10]
  PIN io_wbs_datrd[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 4.000 ;
    END
  END io_wbs_datrd[11]
  PIN io_wbs_datrd[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 0.000 337.090 4.000 ;
    END
  END io_wbs_datrd[12]
  PIN io_wbs_datrd[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END io_wbs_datrd[13]
  PIN io_wbs_datrd[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END io_wbs_datrd[14]
  PIN io_wbs_datrd[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 0.000 399.190 4.000 ;
    END
  END io_wbs_datrd[15]
  PIN io_wbs_datrd[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.610 0.000 419.890 4.000 ;
    END
  END io_wbs_datrd[16]
  PIN io_wbs_datrd[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 0.000 440.590 4.000 ;
    END
  END io_wbs_datrd[17]
  PIN io_wbs_datrd[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 4.000 ;
    END
  END io_wbs_datrd[18]
  PIN io_wbs_datrd[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 0.000 481.990 4.000 ;
    END
  END io_wbs_datrd[19]
  PIN io_wbs_datrd[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END io_wbs_datrd[1]
  PIN io_wbs_datrd[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END io_wbs_datrd[20]
  PIN io_wbs_datrd[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.110 0.000 523.390 4.000 ;
    END
  END io_wbs_datrd[21]
  PIN io_wbs_datrd[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 0.000 544.090 4.000 ;
    END
  END io_wbs_datrd[22]
  PIN io_wbs_datrd[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 0.000 564.790 4.000 ;
    END
  END io_wbs_datrd[23]
  PIN io_wbs_datrd[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 4.000 ;
    END
  END io_wbs_datrd[24]
  PIN io_wbs_datrd[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 0.000 606.190 4.000 ;
    END
  END io_wbs_datrd[25]
  PIN io_wbs_datrd[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.610 0.000 626.890 4.000 ;
    END
  END io_wbs_datrd[26]
  PIN io_wbs_datrd[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 0.000 647.590 4.000 ;
    END
  END io_wbs_datrd[27]
  PIN io_wbs_datrd[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.010 0.000 668.290 4.000 ;
    END
  END io_wbs_datrd[28]
  PIN io_wbs_datrd[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.710 0.000 688.990 4.000 ;
    END
  END io_wbs_datrd[29]
  PIN io_wbs_datrd[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END io_wbs_datrd[2]
  PIN io_wbs_datrd[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.410 0.000 709.690 4.000 ;
    END
  END io_wbs_datrd[30]
  PIN io_wbs_datrd[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 0.000 730.390 4.000 ;
    END
  END io_wbs_datrd[31]
  PIN io_wbs_datrd[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END io_wbs_datrd[3]
  PIN io_wbs_datrd[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END io_wbs_datrd[4]
  PIN io_wbs_datrd[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END io_wbs_datrd[5]
  PIN io_wbs_datrd[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END io_wbs_datrd[6]
  PIN io_wbs_datrd[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 0.000 233.590 4.000 ;
    END
  END io_wbs_datrd[7]
  PIN io_wbs_datrd[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END io_wbs_datrd[8]
  PIN io_wbs_datrd[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
    END
  END io_wbs_datrd[9]
  PIN io_wbs_datwr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END io_wbs_datwr[0]
  PIN io_wbs_datwr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 4.000 ;
    END
  END io_wbs_datwr[10]
  PIN io_wbs_datwr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 4.000 ;
    END
  END io_wbs_datwr[11]
  PIN io_wbs_datwr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 4.000 ;
    END
  END io_wbs_datwr[12]
  PIN io_wbs_datwr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END io_wbs_datwr[13]
  PIN io_wbs_datwr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 0.000 385.390 4.000 ;
    END
  END io_wbs_datwr[14]
  PIN io_wbs_datwr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END io_wbs_datwr[15]
  PIN io_wbs_datwr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 0.000 426.790 4.000 ;
    END
  END io_wbs_datwr[16]
  PIN io_wbs_datwr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 0.000 447.490 4.000 ;
    END
  END io_wbs_datwr[17]
  PIN io_wbs_datwr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 0.000 468.190 4.000 ;
    END
  END io_wbs_datwr[18]
  PIN io_wbs_datwr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 0.000 488.890 4.000 ;
    END
  END io_wbs_datwr[19]
  PIN io_wbs_datwr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 4.000 ;
    END
  END io_wbs_datwr[1]
  PIN io_wbs_datwr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 0.000 509.590 4.000 ;
    END
  END io_wbs_datwr[20]
  PIN io_wbs_datwr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 0.000 530.290 4.000 ;
    END
  END io_wbs_datwr[21]
  PIN io_wbs_datwr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 0.000 550.990 4.000 ;
    END
  END io_wbs_datwr[22]
  PIN io_wbs_datwr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 0.000 571.690 4.000 ;
    END
  END io_wbs_datwr[23]
  PIN io_wbs_datwr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 0.000 592.390 4.000 ;
    END
  END io_wbs_datwr[24]
  PIN io_wbs_datwr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 0.000 613.090 4.000 ;
    END
  END io_wbs_datwr[25]
  PIN io_wbs_datwr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.510 0.000 633.790 4.000 ;
    END
  END io_wbs_datwr[26]
  PIN io_wbs_datwr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.210 0.000 654.490 4.000 ;
    END
  END io_wbs_datwr[27]
  PIN io_wbs_datwr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 0.000 675.190 4.000 ;
    END
  END io_wbs_datwr[28]
  PIN io_wbs_datwr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END io_wbs_datwr[29]
  PIN io_wbs_datwr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END io_wbs_datwr[2]
  PIN io_wbs_datwr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.310 0.000 716.590 4.000 ;
    END
  END io_wbs_datwr[30]
  PIN io_wbs_datwr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 0.000 737.290 4.000 ;
    END
  END io_wbs_datwr[31]
  PIN io_wbs_datwr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END io_wbs_datwr[3]
  PIN io_wbs_datwr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 4.000 ;
    END
  END io_wbs_datwr[4]
  PIN io_wbs_datwr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END io_wbs_datwr[5]
  PIN io_wbs_datwr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 0.000 219.790 4.000 ;
    END
  END io_wbs_datwr[6]
  PIN io_wbs_datwr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 4.000 ;
    END
  END io_wbs_datwr[7]
  PIN io_wbs_datwr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END io_wbs_datwr[8]
  PIN io_wbs_datwr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 4.000 ;
    END
  END io_wbs_datwr[9]
  PIN io_wbs_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END io_wbs_rst
  PIN io_wbs_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END io_wbs_sel[0]
  PIN io_wbs_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END io_wbs_sel[1]
  PIN io_wbs_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END io_wbs_sel[2]
  PIN io_wbs_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END io_wbs_sel[3]
  PIN io_wbs_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END io_wbs_stb
  PIN io_wbs_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END io_wbs_we
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 187.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 187.920 ;
    END
  END vssd1
  PIN web_mem0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 196.000 18.310 200.000 ;
    END
  END web_mem0
  PIN web_mem1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 196.000 381.710 200.000 ;
    END
  END web_mem1
  PIN wmask_mem0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 196.000 36.710 200.000 ;
    END
  END wmask_mem0[0]
  PIN wmask_mem0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 196.000 55.110 200.000 ;
    END
  END wmask_mem0[1]
  PIN wmask_mem0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 196.000 73.510 200.000 ;
    END
  END wmask_mem0[2]
  PIN wmask_mem0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 196.000 91.910 200.000 ;
    END
  END wmask_mem0[3]
  PIN wmask_mem1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.830 196.000 400.110 200.000 ;
    END
  END wmask_mem1[0]
  PIN wmask_mem1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 196.000 418.510 200.000 ;
    END
  END wmask_mem1[1]
  PIN wmask_mem1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.630 196.000 436.910 200.000 ;
    END
  END wmask_mem1[2]
  PIN wmask_mem1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 196.000 455.310 200.000 ;
    END
  END wmask_mem1[3]
  OBS
      LAYER nwell ;
        RECT 5.330 186.265 744.470 187.870 ;
        RECT 5.330 180.825 744.470 183.655 ;
        RECT 5.330 175.385 744.470 178.215 ;
        RECT 5.330 169.945 744.470 172.775 ;
        RECT 5.330 164.505 744.470 167.335 ;
        RECT 5.330 159.065 744.470 161.895 ;
        RECT 5.330 153.625 744.470 156.455 ;
        RECT 5.330 148.185 744.470 151.015 ;
        RECT 5.330 142.745 744.470 145.575 ;
        RECT 5.330 137.305 744.470 140.135 ;
        RECT 5.330 131.865 744.470 134.695 ;
        RECT 5.330 126.425 744.470 129.255 ;
        RECT 5.330 120.985 744.470 123.815 ;
        RECT 5.330 115.545 744.470 118.375 ;
        RECT 5.330 110.105 744.470 112.935 ;
        RECT 5.330 104.665 744.470 107.495 ;
        RECT 5.330 99.225 744.470 102.055 ;
        RECT 5.330 93.785 744.470 96.615 ;
        RECT 5.330 88.345 744.470 91.175 ;
        RECT 5.330 82.905 744.470 85.735 ;
        RECT 5.330 77.465 744.470 80.295 ;
        RECT 5.330 72.025 744.470 74.855 ;
        RECT 5.330 66.585 744.470 69.415 ;
        RECT 5.330 61.145 744.470 63.975 ;
        RECT 5.330 55.705 744.470 58.535 ;
        RECT 5.330 50.265 744.470 53.095 ;
        RECT 5.330 44.825 744.470 47.655 ;
        RECT 5.330 39.385 744.470 42.215 ;
        RECT 5.330 33.945 744.470 36.775 ;
        RECT 5.330 28.505 744.470 31.335 ;
        RECT 5.330 23.065 744.470 25.895 ;
        RECT 5.330 17.625 744.470 20.455 ;
        RECT 5.330 12.185 744.470 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 744.280 187.765 ;
      LAYER met1 ;
        RECT 5.520 7.180 744.280 196.820 ;
      LAYER met2 ;
        RECT 12.520 195.720 13.150 196.850 ;
        RECT 13.990 195.720 17.750 196.850 ;
        RECT 18.590 195.720 22.350 196.850 ;
        RECT 23.190 195.720 26.950 196.850 ;
        RECT 27.790 195.720 31.550 196.850 ;
        RECT 32.390 195.720 36.150 196.850 ;
        RECT 36.990 195.720 40.750 196.850 ;
        RECT 41.590 195.720 45.350 196.850 ;
        RECT 46.190 195.720 49.950 196.850 ;
        RECT 50.790 195.720 54.550 196.850 ;
        RECT 55.390 195.720 59.150 196.850 ;
        RECT 59.990 195.720 63.750 196.850 ;
        RECT 64.590 195.720 68.350 196.850 ;
        RECT 69.190 195.720 72.950 196.850 ;
        RECT 73.790 195.720 77.550 196.850 ;
        RECT 78.390 195.720 82.150 196.850 ;
        RECT 82.990 195.720 86.750 196.850 ;
        RECT 87.590 195.720 91.350 196.850 ;
        RECT 92.190 195.720 95.950 196.850 ;
        RECT 96.790 195.720 100.550 196.850 ;
        RECT 101.390 195.720 105.150 196.850 ;
        RECT 105.990 195.720 109.750 196.850 ;
        RECT 110.590 195.720 114.350 196.850 ;
        RECT 115.190 195.720 118.950 196.850 ;
        RECT 119.790 195.720 123.550 196.850 ;
        RECT 124.390 195.720 128.150 196.850 ;
        RECT 128.990 195.720 132.750 196.850 ;
        RECT 133.590 195.720 137.350 196.850 ;
        RECT 138.190 195.720 141.950 196.850 ;
        RECT 142.790 195.720 146.550 196.850 ;
        RECT 147.390 195.720 151.150 196.850 ;
        RECT 151.990 195.720 155.750 196.850 ;
        RECT 156.590 195.720 160.350 196.850 ;
        RECT 161.190 195.720 164.950 196.850 ;
        RECT 165.790 195.720 169.550 196.850 ;
        RECT 170.390 195.720 174.150 196.850 ;
        RECT 174.990 195.720 178.750 196.850 ;
        RECT 179.590 195.720 183.350 196.850 ;
        RECT 184.190 195.720 187.950 196.850 ;
        RECT 188.790 195.720 192.550 196.850 ;
        RECT 193.390 195.720 197.150 196.850 ;
        RECT 197.990 195.720 201.750 196.850 ;
        RECT 202.590 195.720 206.350 196.850 ;
        RECT 207.190 195.720 210.950 196.850 ;
        RECT 211.790 195.720 215.550 196.850 ;
        RECT 216.390 195.720 220.150 196.850 ;
        RECT 220.990 195.720 224.750 196.850 ;
        RECT 225.590 195.720 229.350 196.850 ;
        RECT 230.190 195.720 233.950 196.850 ;
        RECT 234.790 195.720 238.550 196.850 ;
        RECT 239.390 195.720 243.150 196.850 ;
        RECT 243.990 195.720 247.750 196.850 ;
        RECT 248.590 195.720 252.350 196.850 ;
        RECT 253.190 195.720 256.950 196.850 ;
        RECT 257.790 195.720 261.550 196.850 ;
        RECT 262.390 195.720 266.150 196.850 ;
        RECT 266.990 195.720 270.750 196.850 ;
        RECT 271.590 195.720 275.350 196.850 ;
        RECT 276.190 195.720 279.950 196.850 ;
        RECT 280.790 195.720 284.550 196.850 ;
        RECT 285.390 195.720 289.150 196.850 ;
        RECT 289.990 195.720 293.750 196.850 ;
        RECT 294.590 195.720 298.350 196.850 ;
        RECT 299.190 195.720 302.950 196.850 ;
        RECT 303.790 195.720 307.550 196.850 ;
        RECT 308.390 195.720 312.150 196.850 ;
        RECT 312.990 195.720 316.750 196.850 ;
        RECT 317.590 195.720 321.350 196.850 ;
        RECT 322.190 195.720 325.950 196.850 ;
        RECT 326.790 195.720 330.550 196.850 ;
        RECT 331.390 195.720 335.150 196.850 ;
        RECT 335.990 195.720 339.750 196.850 ;
        RECT 340.590 195.720 344.350 196.850 ;
        RECT 345.190 195.720 348.950 196.850 ;
        RECT 349.790 195.720 353.550 196.850 ;
        RECT 354.390 195.720 358.150 196.850 ;
        RECT 358.990 195.720 362.750 196.850 ;
        RECT 363.590 195.720 367.350 196.850 ;
        RECT 368.190 195.720 371.950 196.850 ;
        RECT 372.790 195.720 376.550 196.850 ;
        RECT 377.390 195.720 381.150 196.850 ;
        RECT 381.990 195.720 385.750 196.850 ;
        RECT 386.590 195.720 390.350 196.850 ;
        RECT 391.190 195.720 394.950 196.850 ;
        RECT 395.790 195.720 399.550 196.850 ;
        RECT 400.390 195.720 404.150 196.850 ;
        RECT 404.990 195.720 408.750 196.850 ;
        RECT 409.590 195.720 413.350 196.850 ;
        RECT 414.190 195.720 417.950 196.850 ;
        RECT 418.790 195.720 422.550 196.850 ;
        RECT 423.390 195.720 427.150 196.850 ;
        RECT 427.990 195.720 431.750 196.850 ;
        RECT 432.590 195.720 436.350 196.850 ;
        RECT 437.190 195.720 440.950 196.850 ;
        RECT 441.790 195.720 445.550 196.850 ;
        RECT 446.390 195.720 450.150 196.850 ;
        RECT 450.990 195.720 454.750 196.850 ;
        RECT 455.590 195.720 459.350 196.850 ;
        RECT 460.190 195.720 463.950 196.850 ;
        RECT 464.790 195.720 468.550 196.850 ;
        RECT 469.390 195.720 473.150 196.850 ;
        RECT 473.990 195.720 477.750 196.850 ;
        RECT 478.590 195.720 482.350 196.850 ;
        RECT 483.190 195.720 486.950 196.850 ;
        RECT 487.790 195.720 491.550 196.850 ;
        RECT 492.390 195.720 496.150 196.850 ;
        RECT 496.990 195.720 500.750 196.850 ;
        RECT 501.590 195.720 505.350 196.850 ;
        RECT 506.190 195.720 509.950 196.850 ;
        RECT 510.790 195.720 514.550 196.850 ;
        RECT 515.390 195.720 519.150 196.850 ;
        RECT 519.990 195.720 523.750 196.850 ;
        RECT 524.590 195.720 528.350 196.850 ;
        RECT 529.190 195.720 532.950 196.850 ;
        RECT 533.790 195.720 537.550 196.850 ;
        RECT 538.390 195.720 542.150 196.850 ;
        RECT 542.990 195.720 546.750 196.850 ;
        RECT 547.590 195.720 551.350 196.850 ;
        RECT 552.190 195.720 555.950 196.850 ;
        RECT 556.790 195.720 560.550 196.850 ;
        RECT 561.390 195.720 565.150 196.850 ;
        RECT 565.990 195.720 569.750 196.850 ;
        RECT 570.590 195.720 574.350 196.850 ;
        RECT 575.190 195.720 578.950 196.850 ;
        RECT 579.790 195.720 583.550 196.850 ;
        RECT 584.390 195.720 588.150 196.850 ;
        RECT 588.990 195.720 592.750 196.850 ;
        RECT 593.590 195.720 597.350 196.850 ;
        RECT 598.190 195.720 601.950 196.850 ;
        RECT 602.790 195.720 606.550 196.850 ;
        RECT 607.390 195.720 611.150 196.850 ;
        RECT 611.990 195.720 615.750 196.850 ;
        RECT 616.590 195.720 620.350 196.850 ;
        RECT 621.190 195.720 624.950 196.850 ;
        RECT 625.790 195.720 629.550 196.850 ;
        RECT 630.390 195.720 634.150 196.850 ;
        RECT 634.990 195.720 638.750 196.850 ;
        RECT 639.590 195.720 643.350 196.850 ;
        RECT 644.190 195.720 647.950 196.850 ;
        RECT 648.790 195.720 652.550 196.850 ;
        RECT 653.390 195.720 657.150 196.850 ;
        RECT 657.990 195.720 661.750 196.850 ;
        RECT 662.590 195.720 666.350 196.850 ;
        RECT 667.190 195.720 670.950 196.850 ;
        RECT 671.790 195.720 675.550 196.850 ;
        RECT 676.390 195.720 680.150 196.850 ;
        RECT 680.990 195.720 684.750 196.850 ;
        RECT 685.590 195.720 689.350 196.850 ;
        RECT 690.190 195.720 693.950 196.850 ;
        RECT 694.790 195.720 698.550 196.850 ;
        RECT 699.390 195.720 703.150 196.850 ;
        RECT 703.990 195.720 707.750 196.850 ;
        RECT 708.590 195.720 712.350 196.850 ;
        RECT 713.190 195.720 716.950 196.850 ;
        RECT 717.790 195.720 721.550 196.850 ;
        RECT 722.390 195.720 726.150 196.850 ;
        RECT 726.990 195.720 730.750 196.850 ;
        RECT 731.590 195.720 735.350 196.850 ;
        RECT 736.190 195.720 737.280 196.850 ;
        RECT 12.520 4.280 737.280 195.720 ;
        RECT 13.070 4.000 19.130 4.280 ;
        RECT 19.970 4.000 26.030 4.280 ;
        RECT 26.870 4.000 32.930 4.280 ;
        RECT 33.770 4.000 39.830 4.280 ;
        RECT 40.670 4.000 46.730 4.280 ;
        RECT 47.570 4.000 53.630 4.280 ;
        RECT 54.470 4.000 60.530 4.280 ;
        RECT 61.370 4.000 67.430 4.280 ;
        RECT 68.270 4.000 74.330 4.280 ;
        RECT 75.170 4.000 81.230 4.280 ;
        RECT 82.070 4.000 88.130 4.280 ;
        RECT 88.970 4.000 95.030 4.280 ;
        RECT 95.870 4.000 101.930 4.280 ;
        RECT 102.770 4.000 108.830 4.280 ;
        RECT 109.670 4.000 115.730 4.280 ;
        RECT 116.570 4.000 122.630 4.280 ;
        RECT 123.470 4.000 129.530 4.280 ;
        RECT 130.370 4.000 136.430 4.280 ;
        RECT 137.270 4.000 143.330 4.280 ;
        RECT 144.170 4.000 150.230 4.280 ;
        RECT 151.070 4.000 157.130 4.280 ;
        RECT 157.970 4.000 164.030 4.280 ;
        RECT 164.870 4.000 170.930 4.280 ;
        RECT 171.770 4.000 177.830 4.280 ;
        RECT 178.670 4.000 184.730 4.280 ;
        RECT 185.570 4.000 191.630 4.280 ;
        RECT 192.470 4.000 198.530 4.280 ;
        RECT 199.370 4.000 205.430 4.280 ;
        RECT 206.270 4.000 212.330 4.280 ;
        RECT 213.170 4.000 219.230 4.280 ;
        RECT 220.070 4.000 226.130 4.280 ;
        RECT 226.970 4.000 233.030 4.280 ;
        RECT 233.870 4.000 239.930 4.280 ;
        RECT 240.770 4.000 246.830 4.280 ;
        RECT 247.670 4.000 253.730 4.280 ;
        RECT 254.570 4.000 260.630 4.280 ;
        RECT 261.470 4.000 267.530 4.280 ;
        RECT 268.370 4.000 274.430 4.280 ;
        RECT 275.270 4.000 281.330 4.280 ;
        RECT 282.170 4.000 288.230 4.280 ;
        RECT 289.070 4.000 295.130 4.280 ;
        RECT 295.970 4.000 302.030 4.280 ;
        RECT 302.870 4.000 308.930 4.280 ;
        RECT 309.770 4.000 315.830 4.280 ;
        RECT 316.670 4.000 322.730 4.280 ;
        RECT 323.570 4.000 329.630 4.280 ;
        RECT 330.470 4.000 336.530 4.280 ;
        RECT 337.370 4.000 343.430 4.280 ;
        RECT 344.270 4.000 350.330 4.280 ;
        RECT 351.170 4.000 357.230 4.280 ;
        RECT 358.070 4.000 364.130 4.280 ;
        RECT 364.970 4.000 371.030 4.280 ;
        RECT 371.870 4.000 377.930 4.280 ;
        RECT 378.770 4.000 384.830 4.280 ;
        RECT 385.670 4.000 391.730 4.280 ;
        RECT 392.570 4.000 398.630 4.280 ;
        RECT 399.470 4.000 405.530 4.280 ;
        RECT 406.370 4.000 412.430 4.280 ;
        RECT 413.270 4.000 419.330 4.280 ;
        RECT 420.170 4.000 426.230 4.280 ;
        RECT 427.070 4.000 433.130 4.280 ;
        RECT 433.970 4.000 440.030 4.280 ;
        RECT 440.870 4.000 446.930 4.280 ;
        RECT 447.770 4.000 453.830 4.280 ;
        RECT 454.670 4.000 460.730 4.280 ;
        RECT 461.570 4.000 467.630 4.280 ;
        RECT 468.470 4.000 474.530 4.280 ;
        RECT 475.370 4.000 481.430 4.280 ;
        RECT 482.270 4.000 488.330 4.280 ;
        RECT 489.170 4.000 495.230 4.280 ;
        RECT 496.070 4.000 502.130 4.280 ;
        RECT 502.970 4.000 509.030 4.280 ;
        RECT 509.870 4.000 515.930 4.280 ;
        RECT 516.770 4.000 522.830 4.280 ;
        RECT 523.670 4.000 529.730 4.280 ;
        RECT 530.570 4.000 536.630 4.280 ;
        RECT 537.470 4.000 543.530 4.280 ;
        RECT 544.370 4.000 550.430 4.280 ;
        RECT 551.270 4.000 557.330 4.280 ;
        RECT 558.170 4.000 564.230 4.280 ;
        RECT 565.070 4.000 571.130 4.280 ;
        RECT 571.970 4.000 578.030 4.280 ;
        RECT 578.870 4.000 584.930 4.280 ;
        RECT 585.770 4.000 591.830 4.280 ;
        RECT 592.670 4.000 598.730 4.280 ;
        RECT 599.570 4.000 605.630 4.280 ;
        RECT 606.470 4.000 612.530 4.280 ;
        RECT 613.370 4.000 619.430 4.280 ;
        RECT 620.270 4.000 626.330 4.280 ;
        RECT 627.170 4.000 633.230 4.280 ;
        RECT 634.070 4.000 640.130 4.280 ;
        RECT 640.970 4.000 647.030 4.280 ;
        RECT 647.870 4.000 653.930 4.280 ;
        RECT 654.770 4.000 660.830 4.280 ;
        RECT 661.670 4.000 667.730 4.280 ;
        RECT 668.570 4.000 674.630 4.280 ;
        RECT 675.470 4.000 681.530 4.280 ;
        RECT 682.370 4.000 688.430 4.280 ;
        RECT 689.270 4.000 695.330 4.280 ;
        RECT 696.170 4.000 702.230 4.280 ;
        RECT 703.070 4.000 709.130 4.280 ;
        RECT 709.970 4.000 716.030 4.280 ;
        RECT 716.870 4.000 722.930 4.280 ;
        RECT 723.770 4.000 729.830 4.280 ;
        RECT 730.670 4.000 736.730 4.280 ;
      LAYER met3 ;
        RECT 21.050 10.715 713.830 188.185 ;
  END
END wb_memory
END LIBRARY

