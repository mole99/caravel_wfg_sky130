magic
tech sky130A
magscale 1 2
timestamp 1669220310
<< obsli1 >>
rect 1104 2159 118864 117521
<< obsm1 >>
rect 14 1504 118864 117552
<< metal2 >>
rect 1950 119200 2006 120000
rect 4526 119200 4582 120000
rect 7102 119200 7158 120000
rect 9678 119200 9734 120000
rect 12254 119200 12310 120000
rect 14830 119200 14886 120000
rect 17406 119200 17462 120000
rect 19982 119200 20038 120000
rect 22558 119200 22614 120000
rect 25134 119200 25190 120000
rect 27710 119200 27766 120000
rect 30286 119200 30342 120000
rect 32862 119200 32918 120000
rect 35438 119200 35494 120000
rect 38014 119200 38070 120000
rect 40590 119200 40646 120000
rect 43166 119200 43222 120000
rect 45742 119200 45798 120000
rect 48318 119200 48374 120000
rect 50894 119200 50950 120000
rect 53470 119200 53526 120000
rect 56046 119200 56102 120000
rect 58622 119200 58678 120000
rect 61198 119200 61254 120000
rect 63774 119200 63830 120000
rect 66350 119200 66406 120000
rect 68926 119200 68982 120000
rect 71502 119200 71558 120000
rect 74078 119200 74134 120000
rect 76654 119200 76710 120000
rect 79230 119200 79286 120000
rect 81806 119200 81862 120000
rect 84382 119200 84438 120000
rect 86958 119200 87014 120000
rect 89534 119200 89590 120000
rect 92110 119200 92166 120000
rect 94686 119200 94742 120000
rect 97262 119200 97318 120000
rect 99838 119200 99894 120000
rect 102414 119200 102470 120000
rect 104990 119200 105046 120000
rect 107566 119200 107622 120000
rect 110142 119200 110198 120000
rect 112718 119200 112774 120000
rect 115294 119200 115350 120000
rect 117870 119200 117926 120000
rect 4158 0 4214 800
rect 5262 0 5318 800
rect 6366 0 6422 800
rect 7470 0 7526 800
rect 8574 0 8630 800
rect 9678 0 9734 800
rect 10782 0 10838 800
rect 11886 0 11942 800
rect 12990 0 13046 800
rect 14094 0 14150 800
rect 15198 0 15254 800
rect 16302 0 16358 800
rect 17406 0 17462 800
rect 18510 0 18566 800
rect 19614 0 19670 800
rect 20718 0 20774 800
rect 21822 0 21878 800
rect 22926 0 22982 800
rect 24030 0 24086 800
rect 25134 0 25190 800
rect 26238 0 26294 800
rect 27342 0 27398 800
rect 28446 0 28502 800
rect 29550 0 29606 800
rect 30654 0 30710 800
rect 31758 0 31814 800
rect 32862 0 32918 800
rect 33966 0 34022 800
rect 35070 0 35126 800
rect 36174 0 36230 800
rect 37278 0 37334 800
rect 38382 0 38438 800
rect 39486 0 39542 800
rect 40590 0 40646 800
rect 41694 0 41750 800
rect 42798 0 42854 800
rect 43902 0 43958 800
rect 45006 0 45062 800
rect 46110 0 46166 800
rect 47214 0 47270 800
rect 48318 0 48374 800
rect 49422 0 49478 800
rect 50526 0 50582 800
rect 51630 0 51686 800
rect 52734 0 52790 800
rect 53838 0 53894 800
rect 54942 0 54998 800
rect 56046 0 56102 800
rect 57150 0 57206 800
rect 58254 0 58310 800
rect 59358 0 59414 800
rect 60462 0 60518 800
rect 61566 0 61622 800
rect 62670 0 62726 800
rect 63774 0 63830 800
rect 64878 0 64934 800
rect 65982 0 66038 800
rect 67086 0 67142 800
rect 68190 0 68246 800
rect 69294 0 69350 800
rect 70398 0 70454 800
rect 71502 0 71558 800
rect 72606 0 72662 800
rect 73710 0 73766 800
rect 74814 0 74870 800
rect 75918 0 75974 800
rect 77022 0 77078 800
rect 78126 0 78182 800
rect 79230 0 79286 800
rect 80334 0 80390 800
rect 81438 0 81494 800
rect 82542 0 82598 800
rect 83646 0 83702 800
rect 84750 0 84806 800
rect 85854 0 85910 800
rect 86958 0 87014 800
rect 88062 0 88118 800
rect 89166 0 89222 800
rect 90270 0 90326 800
rect 91374 0 91430 800
rect 92478 0 92534 800
rect 93582 0 93638 800
rect 94686 0 94742 800
rect 95790 0 95846 800
rect 96894 0 96950 800
rect 97998 0 98054 800
rect 99102 0 99158 800
rect 100206 0 100262 800
rect 101310 0 101366 800
rect 102414 0 102470 800
rect 103518 0 103574 800
rect 104622 0 104678 800
rect 105726 0 105782 800
rect 106830 0 106886 800
rect 107934 0 107990 800
rect 109038 0 109094 800
rect 110142 0 110198 800
rect 111246 0 111302 800
rect 112350 0 112406 800
rect 113454 0 113510 800
rect 114558 0 114614 800
rect 115662 0 115718 800
<< obsm2 >>
rect 18 119144 1894 119354
rect 2062 119144 4470 119354
rect 4638 119144 7046 119354
rect 7214 119144 9622 119354
rect 9790 119144 12198 119354
rect 12366 119144 14774 119354
rect 14942 119144 17350 119354
rect 17518 119144 19926 119354
rect 20094 119144 22502 119354
rect 22670 119144 25078 119354
rect 25246 119144 27654 119354
rect 27822 119144 30230 119354
rect 30398 119144 32806 119354
rect 32974 119144 35382 119354
rect 35550 119144 37958 119354
rect 38126 119144 40534 119354
rect 40702 119144 43110 119354
rect 43278 119144 45686 119354
rect 45854 119144 48262 119354
rect 48430 119144 50838 119354
rect 51006 119144 53414 119354
rect 53582 119144 55990 119354
rect 56158 119144 58566 119354
rect 58734 119144 61142 119354
rect 61310 119144 63718 119354
rect 63886 119144 66294 119354
rect 66462 119144 68870 119354
rect 69038 119144 71446 119354
rect 71614 119144 74022 119354
rect 74190 119144 76598 119354
rect 76766 119144 79174 119354
rect 79342 119144 81750 119354
rect 81918 119144 84326 119354
rect 84494 119144 86902 119354
rect 87070 119144 89478 119354
rect 89646 119144 92054 119354
rect 92222 119144 94630 119354
rect 94798 119144 97206 119354
rect 97374 119144 99782 119354
rect 99950 119144 102358 119354
rect 102526 119144 104934 119354
rect 105102 119144 107510 119354
rect 107678 119144 110086 119354
rect 110254 119144 112662 119354
rect 112830 119144 115238 119354
rect 115406 119144 117814 119354
rect 117982 119144 118200 119354
rect 18 856 118200 119144
rect 18 734 4102 856
rect 4270 734 5206 856
rect 5374 734 6310 856
rect 6478 734 7414 856
rect 7582 734 8518 856
rect 8686 734 9622 856
rect 9790 734 10726 856
rect 10894 734 11830 856
rect 11998 734 12934 856
rect 13102 734 14038 856
rect 14206 734 15142 856
rect 15310 734 16246 856
rect 16414 734 17350 856
rect 17518 734 18454 856
rect 18622 734 19558 856
rect 19726 734 20662 856
rect 20830 734 21766 856
rect 21934 734 22870 856
rect 23038 734 23974 856
rect 24142 734 25078 856
rect 25246 734 26182 856
rect 26350 734 27286 856
rect 27454 734 28390 856
rect 28558 734 29494 856
rect 29662 734 30598 856
rect 30766 734 31702 856
rect 31870 734 32806 856
rect 32974 734 33910 856
rect 34078 734 35014 856
rect 35182 734 36118 856
rect 36286 734 37222 856
rect 37390 734 38326 856
rect 38494 734 39430 856
rect 39598 734 40534 856
rect 40702 734 41638 856
rect 41806 734 42742 856
rect 42910 734 43846 856
rect 44014 734 44950 856
rect 45118 734 46054 856
rect 46222 734 47158 856
rect 47326 734 48262 856
rect 48430 734 49366 856
rect 49534 734 50470 856
rect 50638 734 51574 856
rect 51742 734 52678 856
rect 52846 734 53782 856
rect 53950 734 54886 856
rect 55054 734 55990 856
rect 56158 734 57094 856
rect 57262 734 58198 856
rect 58366 734 59302 856
rect 59470 734 60406 856
rect 60574 734 61510 856
rect 61678 734 62614 856
rect 62782 734 63718 856
rect 63886 734 64822 856
rect 64990 734 65926 856
rect 66094 734 67030 856
rect 67198 734 68134 856
rect 68302 734 69238 856
rect 69406 734 70342 856
rect 70510 734 71446 856
rect 71614 734 72550 856
rect 72718 734 73654 856
rect 73822 734 74758 856
rect 74926 734 75862 856
rect 76030 734 76966 856
rect 77134 734 78070 856
rect 78238 734 79174 856
rect 79342 734 80278 856
rect 80446 734 81382 856
rect 81550 734 82486 856
rect 82654 734 83590 856
rect 83758 734 84694 856
rect 84862 734 85798 856
rect 85966 734 86902 856
rect 87070 734 88006 856
rect 88174 734 89110 856
rect 89278 734 90214 856
rect 90382 734 91318 856
rect 91486 734 92422 856
rect 92590 734 93526 856
rect 93694 734 94630 856
rect 94798 734 95734 856
rect 95902 734 96838 856
rect 97006 734 97942 856
rect 98110 734 99046 856
rect 99214 734 100150 856
rect 100318 734 101254 856
rect 101422 734 102358 856
rect 102526 734 103462 856
rect 103630 734 104566 856
rect 104734 734 105670 856
rect 105838 734 106774 856
rect 106942 734 107878 856
rect 108046 734 108982 856
rect 109150 734 110086 856
rect 110254 734 111190 856
rect 111358 734 112294 856
rect 112462 734 113398 856
rect 113566 734 114502 856
rect 114670 734 115606 856
rect 115774 734 118200 856
<< metal3 >>
rect 0 116968 800 117088
rect 0 114248 800 114368
rect 0 111528 800 111648
rect 0 108808 800 108928
rect 0 106088 800 106208
rect 0 103368 800 103488
rect 0 100648 800 100768
rect 0 97928 800 98048
rect 0 95208 800 95328
rect 0 92488 800 92608
rect 0 89768 800 89888
rect 0 87048 800 87168
rect 0 84328 800 84448
rect 0 81608 800 81728
rect 0 78888 800 79008
rect 0 76168 800 76288
rect 0 73448 800 73568
rect 0 70728 800 70848
rect 0 68008 800 68128
rect 0 65288 800 65408
rect 0 62568 800 62688
rect 0 59848 800 59968
rect 0 57128 800 57248
rect 0 54408 800 54528
rect 0 51688 800 51808
rect 0 48968 800 49088
rect 0 46248 800 46368
rect 0 43528 800 43648
rect 0 40808 800 40928
rect 0 38088 800 38208
rect 0 35368 800 35488
rect 0 32648 800 32768
rect 0 29928 800 30048
rect 0 27208 800 27328
rect 0 24488 800 24608
rect 0 21768 800 21888
rect 0 19048 800 19168
rect 0 16328 800 16448
rect 0 13608 800 13728
rect 0 10888 800 11008
rect 0 8168 800 8288
rect 0 5448 800 5568
rect 0 2728 800 2848
<< obsm3 >>
rect 13 117168 115079 117537
rect 880 116888 115079 117168
rect 13 114448 115079 116888
rect 880 114168 115079 114448
rect 13 111728 115079 114168
rect 880 111448 115079 111728
rect 13 109008 115079 111448
rect 880 108728 115079 109008
rect 13 106288 115079 108728
rect 880 106008 115079 106288
rect 13 103568 115079 106008
rect 880 103288 115079 103568
rect 13 100848 115079 103288
rect 880 100568 115079 100848
rect 13 98128 115079 100568
rect 880 97848 115079 98128
rect 13 95408 115079 97848
rect 880 95128 115079 95408
rect 13 92688 115079 95128
rect 880 92408 115079 92688
rect 13 89968 115079 92408
rect 880 89688 115079 89968
rect 13 87248 115079 89688
rect 880 86968 115079 87248
rect 13 84528 115079 86968
rect 880 84248 115079 84528
rect 13 81808 115079 84248
rect 880 81528 115079 81808
rect 13 79088 115079 81528
rect 880 78808 115079 79088
rect 13 76368 115079 78808
rect 880 76088 115079 76368
rect 13 73648 115079 76088
rect 880 73368 115079 73648
rect 13 70928 115079 73368
rect 880 70648 115079 70928
rect 13 68208 115079 70648
rect 880 67928 115079 68208
rect 13 65488 115079 67928
rect 880 65208 115079 65488
rect 13 62768 115079 65208
rect 880 62488 115079 62768
rect 13 60048 115079 62488
rect 880 59768 115079 60048
rect 13 57328 115079 59768
rect 880 57048 115079 57328
rect 13 54608 115079 57048
rect 880 54328 115079 54608
rect 13 51888 115079 54328
rect 880 51608 115079 51888
rect 13 49168 115079 51608
rect 880 48888 115079 49168
rect 13 46448 115079 48888
rect 880 46168 115079 46448
rect 13 43728 115079 46168
rect 880 43448 115079 43728
rect 13 41008 115079 43448
rect 880 40728 115079 41008
rect 13 38288 115079 40728
rect 880 38008 115079 38288
rect 13 35568 115079 38008
rect 880 35288 115079 35568
rect 13 32848 115079 35288
rect 880 32568 115079 32848
rect 13 30128 115079 32568
rect 880 29848 115079 30128
rect 13 27408 115079 29848
rect 880 27128 115079 27408
rect 13 24688 115079 27128
rect 880 24408 115079 24688
rect 13 21968 115079 24408
rect 880 21688 115079 21968
rect 13 19248 115079 21688
rect 880 18968 115079 19248
rect 13 16528 115079 18968
rect 880 16248 115079 16528
rect 13 13808 115079 16248
rect 880 13528 115079 13808
rect 13 11088 115079 13528
rect 880 10808 115079 11088
rect 13 8368 115079 10808
rect 880 8088 115079 8368
rect 13 5648 115079 8088
rect 880 5368 115079 5648
rect 13 2928 115079 5368
rect 880 2648 115079 2928
rect 13 2143 115079 2648
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
<< obsm4 >>
rect 1347 2619 4128 117197
rect 4608 2619 19488 117197
rect 19968 2619 34848 117197
rect 35328 2619 50208 117197
rect 50688 2619 65568 117197
rect 66048 2619 80928 117197
rect 81408 2619 95253 117197
<< labels >>
rlabel metal3 s 0 5448 800 5568 6 addr1[0]
port 1 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 addr1[1]
port 2 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 addr1[2]
port 3 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 addr1[3]
port 4 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 addr1[4]
port 5 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 addr1[5]
port 6 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 addr1[6]
port 7 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 addr1[7]
port 8 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 addr1[8]
port 9 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 addr1[9]
port 10 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 csb1
port 11 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 dout1[0]
port 12 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 dout1[10]
port 13 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 dout1[11]
port 14 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 dout1[12]
port 15 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 dout1[13]
port 16 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 dout1[14]
port 17 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 dout1[15]
port 18 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 dout1[16]
port 19 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 dout1[17]
port 20 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 dout1[18]
port 21 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 dout1[19]
port 22 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 dout1[1]
port 23 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 dout1[20]
port 24 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 dout1[21]
port 25 nsew signal input
rlabel metal3 s 0 92488 800 92608 6 dout1[22]
port 26 nsew signal input
rlabel metal3 s 0 95208 800 95328 6 dout1[23]
port 27 nsew signal input
rlabel metal3 s 0 97928 800 98048 6 dout1[24]
port 28 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 dout1[25]
port 29 nsew signal input
rlabel metal3 s 0 103368 800 103488 6 dout1[26]
port 30 nsew signal input
rlabel metal3 s 0 106088 800 106208 6 dout1[27]
port 31 nsew signal input
rlabel metal3 s 0 108808 800 108928 6 dout1[28]
port 32 nsew signal input
rlabel metal3 s 0 111528 800 111648 6 dout1[29]
port 33 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 dout1[2]
port 34 nsew signal input
rlabel metal3 s 0 114248 800 114368 6 dout1[30]
port 35 nsew signal input
rlabel metal3 s 0 116968 800 117088 6 dout1[31]
port 36 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 dout1[3]
port 37 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 dout1[4]
port 38 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 dout1[5]
port 39 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 dout1[6]
port 40 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 dout1[7]
port 41 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 dout1[8]
port 42 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 dout1[9]
port 43 nsew signal input
rlabel metal2 s 92110 119200 92166 120000 6 io_oeb[0]
port 44 nsew signal output
rlabel metal2 s 117870 119200 117926 120000 6 io_oeb[10]
port 45 nsew signal output
rlabel metal2 s 94686 119200 94742 120000 6 io_oeb[1]
port 46 nsew signal output
rlabel metal2 s 97262 119200 97318 120000 6 io_oeb[2]
port 47 nsew signal output
rlabel metal2 s 99838 119200 99894 120000 6 io_oeb[3]
port 48 nsew signal output
rlabel metal2 s 102414 119200 102470 120000 6 io_oeb[4]
port 49 nsew signal output
rlabel metal2 s 104990 119200 105046 120000 6 io_oeb[5]
port 50 nsew signal output
rlabel metal2 s 107566 119200 107622 120000 6 io_oeb[6]
port 51 nsew signal output
rlabel metal2 s 110142 119200 110198 120000 6 io_oeb[7]
port 52 nsew signal output
rlabel metal2 s 112718 119200 112774 120000 6 io_oeb[8]
port 53 nsew signal output
rlabel metal2 s 115294 119200 115350 120000 6 io_oeb[9]
port 54 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 io_wbs_ack
port 55 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 io_wbs_adr[0]
port 56 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 io_wbs_adr[10]
port 57 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 io_wbs_adr[11]
port 58 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 io_wbs_adr[12]
port 59 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 io_wbs_adr[13]
port 60 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 io_wbs_adr[14]
port 61 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 io_wbs_adr[15]
port 62 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 io_wbs_adr[16]
port 63 nsew signal input
rlabel metal2 s 67086 0 67142 800 6 io_wbs_adr[17]
port 64 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 io_wbs_adr[18]
port 65 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 io_wbs_adr[19]
port 66 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 io_wbs_adr[1]
port 67 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 io_wbs_adr[20]
port 68 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 io_wbs_adr[21]
port 69 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 io_wbs_adr[22]
port 70 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 io_wbs_adr[23]
port 71 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 io_wbs_adr[24]
port 72 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 io_wbs_adr[25]
port 73 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 io_wbs_adr[26]
port 74 nsew signal input
rlabel metal2 s 100206 0 100262 800 6 io_wbs_adr[27]
port 75 nsew signal input
rlabel metal2 s 103518 0 103574 800 6 io_wbs_adr[28]
port 76 nsew signal input
rlabel metal2 s 106830 0 106886 800 6 io_wbs_adr[29]
port 77 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 io_wbs_adr[2]
port 78 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 io_wbs_adr[30]
port 79 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 io_wbs_adr[31]
port 80 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 io_wbs_adr[3]
port 81 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 io_wbs_adr[4]
port 82 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 io_wbs_adr[5]
port 83 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 io_wbs_adr[6]
port 84 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 io_wbs_adr[7]
port 85 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 io_wbs_adr[8]
port 86 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 io_wbs_adr[9]
port 87 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 io_wbs_clk
port 88 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 io_wbs_cyc
port 89 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 io_wbs_datrd[0]
port 90 nsew signal output
rlabel metal2 s 45006 0 45062 800 6 io_wbs_datrd[10]
port 91 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 io_wbs_datrd[11]
port 92 nsew signal output
rlabel metal2 s 51630 0 51686 800 6 io_wbs_datrd[12]
port 93 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 io_wbs_datrd[13]
port 94 nsew signal output
rlabel metal2 s 58254 0 58310 800 6 io_wbs_datrd[14]
port 95 nsew signal output
rlabel metal2 s 61566 0 61622 800 6 io_wbs_datrd[15]
port 96 nsew signal output
rlabel metal2 s 64878 0 64934 800 6 io_wbs_datrd[16]
port 97 nsew signal output
rlabel metal2 s 68190 0 68246 800 6 io_wbs_datrd[17]
port 98 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 io_wbs_datrd[18]
port 99 nsew signal output
rlabel metal2 s 74814 0 74870 800 6 io_wbs_datrd[19]
port 100 nsew signal output
rlabel metal2 s 15198 0 15254 800 6 io_wbs_datrd[1]
port 101 nsew signal output
rlabel metal2 s 78126 0 78182 800 6 io_wbs_datrd[20]
port 102 nsew signal output
rlabel metal2 s 81438 0 81494 800 6 io_wbs_datrd[21]
port 103 nsew signal output
rlabel metal2 s 84750 0 84806 800 6 io_wbs_datrd[22]
port 104 nsew signal output
rlabel metal2 s 88062 0 88118 800 6 io_wbs_datrd[23]
port 105 nsew signal output
rlabel metal2 s 91374 0 91430 800 6 io_wbs_datrd[24]
port 106 nsew signal output
rlabel metal2 s 94686 0 94742 800 6 io_wbs_datrd[25]
port 107 nsew signal output
rlabel metal2 s 97998 0 98054 800 6 io_wbs_datrd[26]
port 108 nsew signal output
rlabel metal2 s 101310 0 101366 800 6 io_wbs_datrd[27]
port 109 nsew signal output
rlabel metal2 s 104622 0 104678 800 6 io_wbs_datrd[28]
port 110 nsew signal output
rlabel metal2 s 107934 0 107990 800 6 io_wbs_datrd[29]
port 111 nsew signal output
rlabel metal2 s 18510 0 18566 800 6 io_wbs_datrd[2]
port 112 nsew signal output
rlabel metal2 s 111246 0 111302 800 6 io_wbs_datrd[30]
port 113 nsew signal output
rlabel metal2 s 114558 0 114614 800 6 io_wbs_datrd[31]
port 114 nsew signal output
rlabel metal2 s 21822 0 21878 800 6 io_wbs_datrd[3]
port 115 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 io_wbs_datrd[4]
port 116 nsew signal output
rlabel metal2 s 28446 0 28502 800 6 io_wbs_datrd[5]
port 117 nsew signal output
rlabel metal2 s 31758 0 31814 800 6 io_wbs_datrd[6]
port 118 nsew signal output
rlabel metal2 s 35070 0 35126 800 6 io_wbs_datrd[7]
port 119 nsew signal output
rlabel metal2 s 38382 0 38438 800 6 io_wbs_datrd[8]
port 120 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 io_wbs_datrd[9]
port 121 nsew signal output
rlabel metal2 s 12990 0 13046 800 6 io_wbs_datwr[0]
port 122 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 io_wbs_datwr[10]
port 123 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 io_wbs_datwr[11]
port 124 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 io_wbs_datwr[12]
port 125 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 io_wbs_datwr[13]
port 126 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 io_wbs_datwr[14]
port 127 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 io_wbs_datwr[15]
port 128 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 io_wbs_datwr[16]
port 129 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 io_wbs_datwr[17]
port 130 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 io_wbs_datwr[18]
port 131 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 io_wbs_datwr[19]
port 132 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 io_wbs_datwr[1]
port 133 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 io_wbs_datwr[20]
port 134 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 io_wbs_datwr[21]
port 135 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 io_wbs_datwr[22]
port 136 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 io_wbs_datwr[23]
port 137 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 io_wbs_datwr[24]
port 138 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 io_wbs_datwr[25]
port 139 nsew signal input
rlabel metal2 s 99102 0 99158 800 6 io_wbs_datwr[26]
port 140 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 io_wbs_datwr[27]
port 141 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 io_wbs_datwr[28]
port 142 nsew signal input
rlabel metal2 s 109038 0 109094 800 6 io_wbs_datwr[29]
port 143 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 io_wbs_datwr[2]
port 144 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 io_wbs_datwr[30]
port 145 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 io_wbs_datwr[31]
port 146 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 io_wbs_datwr[3]
port 147 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 io_wbs_datwr[4]
port 148 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 io_wbs_datwr[5]
port 149 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 io_wbs_datwr[6]
port 150 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 io_wbs_datwr[7]
port 151 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 io_wbs_datwr[8]
port 152 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 io_wbs_datwr[9]
port 153 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 io_wbs_rst
port 154 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 io_wbs_stb
port 155 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 io_wbs_we
port 156 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 157 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 157 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 157 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 157 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 158 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 158 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 158 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 158 nsew ground bidirectional
rlabel metal2 s 9678 119200 9734 120000 6 wfg_drive_pat_dout_o[0]
port 159 nsew signal output
rlabel metal2 s 35438 119200 35494 120000 6 wfg_drive_pat_dout_o[10]
port 160 nsew signal output
rlabel metal2 s 38014 119200 38070 120000 6 wfg_drive_pat_dout_o[11]
port 161 nsew signal output
rlabel metal2 s 40590 119200 40646 120000 6 wfg_drive_pat_dout_o[12]
port 162 nsew signal output
rlabel metal2 s 43166 119200 43222 120000 6 wfg_drive_pat_dout_o[13]
port 163 nsew signal output
rlabel metal2 s 45742 119200 45798 120000 6 wfg_drive_pat_dout_o[14]
port 164 nsew signal output
rlabel metal2 s 48318 119200 48374 120000 6 wfg_drive_pat_dout_o[15]
port 165 nsew signal output
rlabel metal2 s 50894 119200 50950 120000 6 wfg_drive_pat_dout_o[16]
port 166 nsew signal output
rlabel metal2 s 53470 119200 53526 120000 6 wfg_drive_pat_dout_o[17]
port 167 nsew signal output
rlabel metal2 s 56046 119200 56102 120000 6 wfg_drive_pat_dout_o[18]
port 168 nsew signal output
rlabel metal2 s 58622 119200 58678 120000 6 wfg_drive_pat_dout_o[19]
port 169 nsew signal output
rlabel metal2 s 12254 119200 12310 120000 6 wfg_drive_pat_dout_o[1]
port 170 nsew signal output
rlabel metal2 s 61198 119200 61254 120000 6 wfg_drive_pat_dout_o[20]
port 171 nsew signal output
rlabel metal2 s 63774 119200 63830 120000 6 wfg_drive_pat_dout_o[21]
port 172 nsew signal output
rlabel metal2 s 66350 119200 66406 120000 6 wfg_drive_pat_dout_o[22]
port 173 nsew signal output
rlabel metal2 s 68926 119200 68982 120000 6 wfg_drive_pat_dout_o[23]
port 174 nsew signal output
rlabel metal2 s 71502 119200 71558 120000 6 wfg_drive_pat_dout_o[24]
port 175 nsew signal output
rlabel metal2 s 74078 119200 74134 120000 6 wfg_drive_pat_dout_o[25]
port 176 nsew signal output
rlabel metal2 s 76654 119200 76710 120000 6 wfg_drive_pat_dout_o[26]
port 177 nsew signal output
rlabel metal2 s 79230 119200 79286 120000 6 wfg_drive_pat_dout_o[27]
port 178 nsew signal output
rlabel metal2 s 81806 119200 81862 120000 6 wfg_drive_pat_dout_o[28]
port 179 nsew signal output
rlabel metal2 s 84382 119200 84438 120000 6 wfg_drive_pat_dout_o[29]
port 180 nsew signal output
rlabel metal2 s 14830 119200 14886 120000 6 wfg_drive_pat_dout_o[2]
port 181 nsew signal output
rlabel metal2 s 86958 119200 87014 120000 6 wfg_drive_pat_dout_o[30]
port 182 nsew signal output
rlabel metal2 s 89534 119200 89590 120000 6 wfg_drive_pat_dout_o[31]
port 183 nsew signal output
rlabel metal2 s 17406 119200 17462 120000 6 wfg_drive_pat_dout_o[3]
port 184 nsew signal output
rlabel metal2 s 19982 119200 20038 120000 6 wfg_drive_pat_dout_o[4]
port 185 nsew signal output
rlabel metal2 s 22558 119200 22614 120000 6 wfg_drive_pat_dout_o[5]
port 186 nsew signal output
rlabel metal2 s 25134 119200 25190 120000 6 wfg_drive_pat_dout_o[6]
port 187 nsew signal output
rlabel metal2 s 27710 119200 27766 120000 6 wfg_drive_pat_dout_o[7]
port 188 nsew signal output
rlabel metal2 s 30286 119200 30342 120000 6 wfg_drive_pat_dout_o[8]
port 189 nsew signal output
rlabel metal2 s 32862 119200 32918 120000 6 wfg_drive_pat_dout_o[9]
port 190 nsew signal output
rlabel metal2 s 1950 119200 2006 120000 6 wfg_drive_spi_cs_no
port 191 nsew signal output
rlabel metal2 s 4526 119200 4582 120000 6 wfg_drive_spi_sclk_o
port 192 nsew signal output
rlabel metal2 s 7102 119200 7158 120000 6 wfg_drive_spi_sdo_o
port 193 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 120000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 38057244
string GDS_FILE /home/leo/Dokumente/workspace-sky-mpw-7-redesign/caravel_wfg_sky130/openlane/wfg_top/runs/22_11_23_17_05/results/signoff/wfg_top.magic.gds
string GDS_START 1365564
<< end >>

