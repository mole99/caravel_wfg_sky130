magic
tech sky130A
magscale 1 2
timestamp 1669219296
<< viali >>
rect 2789 37417 2823 37451
rect 44465 37417 44499 37451
rect 45385 37417 45419 37451
rect 50353 37417 50387 37451
rect 54217 37417 54251 37451
rect 55597 37417 55631 37451
rect 58081 37417 58115 37451
rect 59369 37417 59403 37451
rect 80345 37417 80379 37451
rect 84025 37417 84059 37451
rect 89821 37417 89855 37451
rect 94237 37417 94271 37451
rect 95065 37417 95099 37451
rect 97549 37417 97583 37451
rect 99481 37417 99515 37451
rect 101965 37417 101999 37451
rect 103529 37417 103563 37451
rect 120089 37417 120123 37451
rect 121469 37417 121503 37451
rect 122573 37417 122607 37451
rect 125977 37417 126011 37451
rect 29193 37349 29227 37383
rect 59829 37349 59863 37383
rect 60841 37349 60875 37383
rect 67557 37349 67591 37383
rect 136189 37349 136223 37383
rect 138029 37349 138063 37383
rect 25053 37281 25087 37315
rect 27997 37281 28031 37315
rect 28089 37281 28123 37315
rect 30021 37281 30055 37315
rect 33609 37281 33643 37315
rect 35633 37281 35667 37315
rect 36829 37281 36863 37315
rect 38577 37281 38611 37315
rect 41337 37281 41371 37315
rect 42073 37281 42107 37315
rect 46213 37281 46247 37315
rect 47961 37281 47995 37315
rect 48145 37281 48179 37315
rect 51733 37281 51767 37315
rect 53021 37281 53055 37315
rect 57437 37281 57471 37315
rect 58633 37281 58667 37315
rect 61301 37281 61335 37315
rect 61485 37281 61519 37315
rect 63417 37281 63451 37315
rect 64613 37281 64647 37315
rect 64705 37281 64739 37315
rect 66361 37281 66395 37315
rect 68477 37281 68511 37315
rect 71053 37281 71087 37315
rect 72985 37281 73019 37315
rect 75561 37281 75595 37315
rect 77033 37281 77067 37315
rect 79517 37281 79551 37315
rect 79701 37281 79735 37315
rect 81449 37281 81483 37315
rect 81541 37281 81575 37315
rect 83013 37281 83047 37315
rect 105921 37281 105955 37315
rect 110337 37281 110371 37315
rect 116225 37281 116259 37315
rect 118065 37281 118099 37315
rect 120641 37281 120675 37315
rect 4905 37213 4939 37247
rect 5825 37213 5859 37247
rect 6745 37213 6779 37247
rect 7665 37213 7699 37247
rect 8585 37213 8619 37247
rect 9505 37213 9539 37247
rect 10149 37213 10183 37247
rect 11161 37213 11195 37247
rect 12265 37213 12299 37247
rect 13185 37213 13219 37247
rect 15025 37213 15059 37247
rect 15945 37213 15979 37247
rect 17141 37213 17175 37247
rect 17601 37213 17635 37247
rect 18705 37213 18739 37247
rect 19717 37213 19751 37247
rect 20545 37213 20579 37247
rect 21189 37213 21223 37247
rect 22385 37213 22419 37247
rect 23305 37213 23339 37247
rect 24041 37213 24075 37247
rect 26341 37213 26375 37247
rect 27353 37213 27387 37247
rect 29009 37213 29043 37247
rect 31585 37213 31619 37247
rect 32321 37213 32355 37247
rect 34345 37213 34379 37247
rect 38301 37213 38335 37247
rect 39405 37213 39439 37247
rect 40049 37213 40083 37247
rect 42993 37213 43027 37247
rect 44557 37213 44591 37247
rect 45293 37213 45327 37247
rect 46029 37213 46063 37247
rect 46949 37213 46983 37247
rect 49801 37213 49835 37247
rect 51181 37213 51215 37247
rect 52009 37213 52043 37247
rect 54953 37213 54987 37247
rect 56057 37213 56091 37247
rect 61209 37213 61243 37247
rect 62221 37213 62255 37247
rect 63509 37213 63543 37247
rect 64797 37213 64831 37247
rect 70225 37213 70259 37247
rect 72433 37213 72467 37247
rect 74641 37213 74675 37247
rect 77585 37213 77619 37247
rect 80437 37213 80471 37247
rect 82829 37213 82863 37247
rect 84853 37213 84887 37247
rect 85313 37213 85347 37247
rect 86693 37213 86727 37247
rect 87429 37213 87463 37247
rect 88165 37213 88199 37247
rect 89269 37213 89303 37247
rect 90741 37213 90775 37247
rect 91569 37213 91603 37247
rect 92305 37213 92339 37247
rect 93041 37213 93075 37247
rect 94329 37213 94363 37247
rect 95893 37213 95927 37247
rect 96997 37213 97031 37247
rect 98469 37213 98503 37247
rect 100033 37213 100067 37247
rect 100769 37213 100803 37247
rect 102885 37213 102919 37247
rect 104449 37213 104483 37247
rect 105185 37213 105219 37247
rect 107301 37213 107335 37247
rect 107761 37213 107795 37247
rect 108589 37213 108623 37247
rect 109601 37213 109635 37247
rect 111073 37213 111107 37247
rect 112177 37213 112211 37247
rect 112913 37213 112947 37247
rect 113649 37213 113683 37247
rect 114753 37213 114787 37247
rect 115489 37213 115523 37247
rect 116409 37213 116443 37247
rect 117329 37213 117363 37247
rect 119077 37213 119111 37247
rect 119905 37213 119939 37247
rect 121653 37213 121687 37247
rect 122757 37213 122791 37247
rect 123217 37213 123251 37247
rect 124229 37213 124263 37247
rect 125057 37213 125091 37247
rect 125793 37213 125827 37247
rect 126529 37213 126563 37247
rect 127633 37213 127667 37247
rect 128369 37213 128403 37247
rect 129105 37213 129139 37247
rect 130209 37213 130243 37247
rect 131221 37213 131255 37247
rect 131681 37213 131715 37247
rect 133061 37213 133095 37247
rect 133521 37213 133555 37247
rect 134349 37213 134383 37247
rect 135361 37213 135395 37247
rect 137109 37213 137143 37247
rect 138213 37213 138247 37247
rect 138949 37213 138983 37247
rect 139685 37213 139719 37247
rect 140513 37213 140547 37247
rect 141249 37213 141283 37247
rect 142261 37213 142295 37247
rect 143089 37213 143123 37247
rect 143825 37213 143859 37247
rect 144561 37213 144595 37247
rect 145665 37213 145699 37247
rect 146401 37213 146435 37247
rect 147229 37213 147263 37247
rect 25237 37145 25271 37179
rect 29837 37145 29871 37179
rect 30665 37145 30699 37179
rect 30849 37145 30883 37179
rect 33425 37145 33459 37179
rect 35357 37145 35391 37179
rect 35541 37145 35575 37179
rect 41153 37145 41187 37179
rect 43269 37145 43303 37179
rect 48237 37145 48271 37179
rect 53297 37145 53331 37179
rect 60013 37145 60047 37179
rect 62405 37145 62439 37179
rect 66269 37145 66303 37179
rect 66361 37145 66395 37179
rect 67741 37145 67775 37179
rect 68569 37145 68603 37179
rect 68753 37145 68787 37179
rect 71237 37145 71271 37179
rect 73629 37145 73663 37179
rect 73813 37145 73847 37179
rect 75377 37145 75411 37179
rect 76757 37145 76791 37179
rect 79425 37145 79459 37179
rect 81633 37145 81667 37179
rect 83933 37145 83967 37179
rect 89913 37145 89947 37179
rect 94973 37145 95007 37179
rect 97641 37145 97675 37179
rect 99389 37145 99423 37179
rect 102057 37145 102091 37179
rect 103437 37145 103471 37179
rect 106105 37145 106139 37179
rect 110521 37145 110555 37179
rect 118249 37145 118283 37179
rect 120825 37145 120859 37179
rect 136373 37145 136407 37179
rect 4721 37077 4755 37111
rect 5641 37077 5675 37111
rect 6561 37077 6595 37111
rect 7481 37077 7515 37111
rect 8401 37077 8435 37111
rect 9321 37077 9355 37111
rect 10333 37077 10367 37111
rect 10977 37077 11011 37111
rect 12081 37077 12115 37111
rect 13001 37077 13035 37111
rect 14841 37077 14875 37111
rect 15761 37077 15795 37111
rect 16957 37077 16991 37111
rect 17785 37077 17819 37111
rect 18521 37077 18555 37111
rect 19533 37077 19567 37111
rect 20361 37077 20395 37111
rect 21373 37077 21407 37111
rect 22201 37077 22235 37111
rect 23121 37077 23155 37111
rect 23857 37077 23891 37111
rect 24667 37077 24701 37111
rect 25145 37077 25179 37111
rect 25789 37077 25823 37111
rect 26525 37077 26559 37111
rect 27169 37077 27203 37111
rect 28181 37077 28215 37111
rect 28549 37077 28583 37111
rect 31401 37077 31435 37111
rect 32505 37077 32539 37111
rect 34161 37077 34195 37111
rect 35063 37077 35097 37111
rect 36185 37077 36219 37111
rect 36553 37077 36587 37111
rect 36645 37077 36679 37111
rect 37933 37077 37967 37111
rect 38393 37077 38427 37111
rect 39221 37077 39255 37111
rect 40233 37077 40267 37111
rect 40785 37077 40819 37111
rect 41245 37077 41279 37111
rect 43085 37077 43119 37111
rect 43555 37077 43589 37111
rect 47133 37077 47167 37111
rect 48605 37077 48639 37111
rect 49617 37077 49651 37111
rect 50997 37077 51031 37111
rect 51917 37077 51951 37111
rect 52377 37077 52411 37111
rect 53205 37077 53239 37111
rect 53665 37077 53699 37111
rect 54769 37077 54803 37111
rect 56241 37077 56275 37111
rect 56793 37077 56827 37111
rect 57161 37077 57195 37111
rect 57253 37077 57287 37111
rect 58449 37077 58483 37111
rect 58541 37077 58575 37111
rect 62037 37077 62071 37111
rect 63601 37077 63635 37111
rect 63969 37077 64003 37111
rect 65165 37077 65199 37111
rect 66831 37077 66865 37111
rect 69039 37077 69073 37111
rect 70041 37077 70075 37111
rect 71329 37077 71363 37111
rect 71697 37077 71731 37111
rect 72249 37077 72283 37111
rect 74457 37077 74491 37111
rect 76471 37077 76505 37111
rect 76941 37077 76975 37111
rect 77769 37077 77803 37111
rect 79057 37077 79091 37111
rect 82001 37077 82035 37111
rect 82461 37077 82495 37111
rect 82921 37077 82955 37111
rect 84669 37077 84703 37111
rect 85497 37077 85531 37111
rect 86509 37077 86543 37111
rect 87245 37077 87279 37111
rect 87981 37077 88015 37111
rect 89085 37077 89119 37111
rect 90557 37077 90591 37111
rect 91753 37077 91787 37111
rect 92489 37077 92523 37111
rect 93225 37077 93259 37111
rect 95709 37077 95743 37111
rect 96813 37077 96847 37111
rect 98285 37077 98319 37111
rect 100217 37077 100251 37111
rect 100953 37077 100987 37111
rect 102701 37077 102735 37111
rect 104633 37077 104667 37111
rect 105369 37077 105403 37111
rect 107117 37077 107151 37111
rect 107945 37077 107979 37111
rect 108773 37077 108807 37111
rect 109785 37077 109819 37111
rect 111257 37077 111291 37111
rect 112361 37077 112395 37111
rect 113097 37077 113131 37111
rect 113833 37077 113867 37111
rect 114937 37077 114971 37111
rect 115673 37077 115707 37111
rect 117513 37077 117547 37111
rect 118893 37077 118927 37111
rect 123401 37077 123435 37111
rect 124045 37077 124079 37111
rect 125241 37077 125275 37111
rect 126713 37077 126747 37111
rect 127817 37077 127851 37111
rect 128553 37077 128587 37111
rect 129289 37077 129323 37111
rect 130393 37077 130427 37111
rect 131037 37077 131071 37111
rect 131865 37077 131899 37111
rect 132877 37077 132911 37111
rect 133705 37077 133739 37111
rect 134533 37077 134567 37111
rect 135545 37077 135579 37111
rect 137293 37077 137327 37111
rect 139133 37077 139167 37111
rect 139869 37077 139903 37111
rect 140697 37077 140731 37111
rect 141433 37077 141467 37111
rect 142077 37077 142111 37111
rect 143273 37077 143307 37111
rect 144009 37077 144043 37111
rect 144745 37077 144779 37111
rect 145849 37077 145883 37111
rect 146585 37077 146619 37111
rect 147413 37077 147447 37111
rect 3801 36873 3835 36907
rect 4537 36873 4571 36907
rect 8217 36873 8251 36907
rect 9781 36873 9815 36907
rect 12449 36873 12483 36907
rect 17325 36873 17359 36907
rect 19073 36873 19107 36907
rect 20637 36873 20671 36907
rect 28365 36873 28399 36907
rect 28917 36873 28951 36907
rect 29653 36873 29687 36907
rect 30481 36873 30515 36907
rect 32321 36873 32355 36907
rect 33241 36873 33275 36907
rect 34253 36873 34287 36907
rect 36737 36873 36771 36907
rect 42625 36873 42659 36907
rect 42993 36873 43027 36907
rect 43913 36873 43947 36907
rect 58449 36873 58483 36907
rect 60289 36873 60323 36907
rect 62681 36873 62715 36907
rect 65441 36873 65475 36907
rect 66361 36873 66395 36907
rect 67373 36873 67407 36907
rect 72893 36873 72927 36907
rect 76573 36873 76607 36907
rect 77125 36873 77159 36907
rect 78781 36873 78815 36907
rect 80161 36873 80195 36907
rect 119905 36873 119939 36907
rect 124413 36873 124447 36907
rect 125057 36873 125091 36907
rect 125609 36873 125643 36907
rect 126529 36873 126563 36907
rect 127725 36873 127759 36907
rect 128369 36873 128403 36907
rect 128921 36873 128955 36907
rect 131497 36873 131531 36907
rect 132233 36873 132267 36907
rect 133245 36873 133279 36907
rect 134257 36873 134291 36907
rect 136005 36873 136039 36907
rect 137845 36873 137879 36907
rect 140513 36873 140547 36907
rect 141617 36873 141651 36907
rect 143825 36873 143859 36907
rect 145113 36873 145147 36907
rect 146309 36873 146343 36907
rect 147321 36873 147355 36907
rect 24501 36805 24535 36839
rect 37731 36805 37765 36839
rect 38669 36805 38703 36839
rect 41153 36805 41187 36839
rect 65349 36805 65383 36839
rect 87521 36805 87555 36839
rect 96997 36805 97031 36839
rect 99389 36805 99423 36839
rect 99849 36805 99883 36839
rect 103805 36805 103839 36839
rect 105369 36805 105403 36839
rect 105553 36805 105587 36839
rect 108037 36805 108071 36839
rect 108589 36805 108623 36839
rect 112637 36805 112671 36839
rect 113281 36805 113315 36839
rect 116225 36805 116259 36839
rect 142629 36805 142663 36839
rect 3985 36737 4019 36771
rect 6561 36737 6595 36771
rect 7205 36737 7239 36771
rect 8401 36737 8435 36771
rect 9965 36737 9999 36771
rect 13829 36737 13863 36771
rect 14473 36737 14507 36771
rect 17509 36737 17543 36771
rect 19257 36737 19291 36771
rect 19901 36737 19935 36771
rect 20821 36737 20855 36771
rect 21465 36737 21499 36771
rect 22017 36737 22051 36771
rect 22753 36737 22787 36771
rect 23305 36737 23339 36771
rect 25329 36737 25363 36771
rect 25789 36737 25823 36771
rect 27997 36737 28031 36771
rect 29101 36737 29135 36771
rect 30665 36737 30699 36771
rect 31125 36737 31159 36771
rect 31769 36737 31803 36771
rect 32505 36737 32539 36771
rect 33425 36737 33459 36771
rect 34069 36737 34103 36771
rect 35265 36737 35299 36771
rect 36001 36737 36035 36771
rect 36914 36737 36948 36771
rect 38853 36737 38887 36771
rect 39865 36737 39899 36771
rect 40601 36737 40635 36771
rect 41889 36737 41923 36771
rect 44097 36737 44131 36771
rect 44649 36737 44683 36771
rect 45293 36737 45327 36771
rect 46305 36737 46339 36771
rect 47225 36737 47259 36771
rect 48145 36737 48179 36771
rect 49065 36737 49099 36771
rect 50261 36737 50295 36771
rect 50445 36737 50479 36771
rect 51641 36737 51675 36771
rect 52101 36737 52135 36771
rect 52285 36737 52319 36771
rect 53573 36737 53607 36771
rect 54309 36737 54343 36771
rect 54953 36737 54987 36771
rect 55597 36737 55631 36771
rect 55781 36737 55815 36771
rect 56333 36737 56367 36771
rect 57161 36737 57195 36771
rect 59369 36737 59403 36771
rect 59553 36737 59587 36771
rect 60105 36737 60139 36771
rect 60933 36737 60967 36771
rect 61669 36737 61703 36771
rect 62497 36737 62531 36771
rect 63233 36737 63267 36771
rect 64245 36737 64279 36771
rect 64337 36737 64371 36771
rect 66545 36737 66579 36771
rect 67189 36737 67223 36771
rect 68661 36737 68695 36771
rect 68845 36737 68879 36771
rect 69489 36737 69523 36771
rect 69673 36737 69707 36771
rect 70409 36737 70443 36771
rect 70869 36737 70903 36771
rect 72249 36737 72283 36771
rect 72709 36737 72743 36771
rect 75285 36737 75319 36771
rect 76389 36737 76423 36771
rect 78965 36737 78999 36771
rect 80069 36737 80103 36771
rect 81265 36737 81299 36771
rect 82093 36737 82127 36771
rect 82277 36737 82311 36771
rect 83105 36737 83139 36771
rect 83841 36737 83875 36771
rect 84945 36737 84979 36771
rect 85129 36737 85163 36771
rect 86325 36737 86359 36771
rect 89269 36737 89303 36771
rect 90373 36737 90407 36771
rect 91017 36737 91051 36771
rect 93041 36737 93075 36771
rect 93225 36737 93259 36771
rect 95249 36737 95283 36771
rect 95985 36737 96019 36771
rect 98469 36737 98503 36771
rect 101229 36737 101263 36771
rect 103069 36737 103103 36771
rect 106381 36737 106415 36771
rect 106841 36737 106875 36771
rect 107485 36737 107519 36771
rect 110797 36737 110831 36771
rect 111441 36737 111475 36771
rect 112453 36737 112487 36771
rect 113741 36737 113775 36771
rect 113925 36737 113959 36771
rect 115029 36737 115063 36771
rect 115673 36737 115707 36771
rect 117145 36737 117179 36771
rect 117881 36737 117915 36771
rect 118065 36737 118099 36771
rect 118709 36737 118743 36771
rect 121009 36737 121043 36771
rect 121469 36737 121503 36771
rect 123217 36737 123251 36771
rect 123861 36737 123895 36771
rect 126713 36737 126747 36771
rect 129565 36737 129599 36771
rect 130485 36737 130519 36771
rect 132049 36737 132083 36771
rect 132693 36737 132727 36771
rect 135821 36737 135855 36771
rect 136465 36737 136499 36771
rect 137661 36737 137695 36771
rect 138305 36737 138339 36771
rect 141433 36737 141467 36771
rect 143641 36737 143675 36771
rect 144285 36737 144319 36771
rect 146125 36737 146159 36771
rect 146769 36737 146803 36771
rect 18521 36669 18555 36703
rect 24409 36669 24443 36703
rect 24593 36669 24627 36703
rect 27813 36669 27847 36703
rect 27905 36669 27939 36703
rect 43085 36669 43119 36703
rect 43177 36669 43211 36703
rect 47869 36669 47903 36703
rect 48053 36669 48087 36703
rect 58265 36669 58299 36703
rect 58357 36669 58391 36703
rect 61945 36669 61979 36703
rect 64521 36669 64555 36703
rect 65165 36669 65199 36703
rect 80345 36669 80379 36703
rect 80989 36669 81023 36703
rect 81173 36669 81207 36703
rect 85681 36669 85715 36703
rect 142077 36669 142111 36703
rect 6745 36601 6779 36635
rect 14013 36601 14047 36635
rect 19717 36601 19751 36635
rect 39681 36601 39715 36635
rect 40417 36601 40451 36635
rect 41337 36601 41371 36635
rect 44833 36601 44867 36635
rect 46121 36601 46155 36635
rect 48513 36601 48547 36635
rect 50997 36601 51031 36635
rect 53021 36601 53055 36635
rect 73629 36601 73663 36635
rect 74825 36601 74859 36635
rect 123401 36601 123435 36635
rect 8953 36533 8987 36567
rect 10517 36533 10551 36567
rect 16129 36533 16163 36567
rect 17969 36533 18003 36567
rect 21281 36533 21315 36567
rect 22201 36533 22235 36567
rect 23489 36533 23523 36567
rect 24041 36533 24075 36567
rect 25145 36533 25179 36567
rect 25973 36533 26007 36567
rect 26617 36533 26651 36567
rect 35357 36533 35391 36567
rect 36093 36533 36127 36567
rect 37841 36533 37875 36567
rect 41981 36533 42015 36567
rect 45477 36533 45511 36567
rect 47041 36533 47075 36567
rect 49157 36533 49191 36567
rect 51457 36533 51491 36567
rect 53665 36533 53699 36567
rect 54401 36533 54435 36567
rect 55137 36533 55171 36567
rect 56517 36533 56551 36567
rect 57069 36533 57103 36567
rect 58817 36533 58851 36567
rect 61025 36533 61059 36567
rect 63417 36533 63451 36567
rect 63877 36533 63911 36567
rect 65809 36533 65843 36567
rect 71053 36533 71087 36567
rect 71697 36533 71731 36567
rect 74089 36533 74123 36567
rect 75377 36533 75411 36567
rect 75745 36533 75779 36567
rect 77769 36533 77803 36567
rect 79701 36533 79735 36567
rect 81633 36533 81667 36567
rect 82921 36533 82955 36567
rect 84025 36533 84059 36567
rect 86417 36533 86451 36567
rect 86969 36533 87003 36567
rect 88073 36533 88107 36567
rect 89453 36533 89487 36567
rect 90465 36533 90499 36567
rect 91569 36533 91603 36567
rect 92121 36533 92155 36567
rect 94237 36533 94271 36567
rect 95065 36533 95099 36567
rect 95801 36533 95835 36567
rect 96445 36533 96479 36567
rect 98009 36533 98043 36567
rect 98653 36533 98687 36567
rect 100769 36533 100803 36567
rect 101413 36533 101447 36567
rect 102241 36533 102275 36567
rect 103253 36533 103287 36567
rect 104449 36533 104483 36567
rect 106197 36533 106231 36567
rect 107025 36533 107059 36567
rect 109601 36533 109635 36567
rect 110337 36533 110371 36567
rect 110981 36533 111015 36567
rect 115213 36533 115247 36567
rect 119169 36533 119203 36567
rect 121653 36533 121687 36567
rect 122757 36533 122791 36567
rect 127173 36533 127207 36567
rect 130301 36533 130335 36567
rect 130945 36533 130979 36567
rect 139501 36533 139535 36567
rect 10057 36329 10091 36363
rect 17417 36329 17451 36363
rect 22477 36329 22511 36363
rect 23489 36329 23523 36363
rect 24961 36329 24995 36363
rect 25881 36329 25915 36363
rect 27721 36329 27755 36363
rect 29745 36329 29779 36363
rect 30757 36329 30791 36363
rect 33793 36329 33827 36363
rect 39497 36329 39531 36363
rect 42441 36329 42475 36363
rect 43453 36329 43487 36363
rect 44281 36329 44315 36363
rect 53481 36329 53515 36363
rect 54217 36329 54251 36363
rect 54769 36329 54803 36363
rect 55873 36329 55907 36363
rect 59645 36329 59679 36363
rect 62681 36329 62715 36363
rect 64521 36329 64555 36363
rect 67097 36329 67131 36363
rect 68201 36329 68235 36363
rect 70409 36329 70443 36363
rect 72617 36329 72651 36363
rect 74089 36329 74123 36363
rect 74733 36329 74767 36363
rect 76297 36329 76331 36363
rect 80253 36329 80287 36363
rect 90741 36329 90775 36363
rect 93961 36329 93995 36363
rect 102977 36329 103011 36363
rect 103437 36329 103471 36363
rect 105001 36329 105035 36363
rect 106381 36329 106415 36363
rect 107117 36329 107151 36363
rect 107669 36329 107703 36363
rect 110889 36329 110923 36363
rect 115305 36329 115339 36363
rect 117881 36329 117915 36363
rect 136097 36329 136131 36363
rect 138029 36329 138063 36363
rect 143641 36329 143675 36363
rect 24041 36261 24075 36295
rect 34253 36261 34287 36295
rect 36093 36261 36127 36295
rect 37289 36261 37323 36295
rect 37933 36261 37967 36295
rect 41613 36261 41647 36295
rect 49525 36261 49559 36295
rect 50813 36261 50847 36295
rect 52193 36261 52227 36295
rect 60841 36261 60875 36295
rect 69213 36261 69247 36295
rect 70961 36261 70995 36295
rect 78689 36261 78723 36295
rect 121101 36261 121135 36295
rect 126437 36261 126471 36295
rect 46489 36193 46523 36227
rect 48145 36193 48179 36227
rect 67649 36193 67683 36227
rect 81357 36193 81391 36227
rect 82461 36193 82495 36227
rect 105829 36193 105863 36227
rect 20177 36125 20211 36159
rect 21189 36125 21223 36159
rect 21833 36125 21867 36159
rect 25145 36125 25179 36159
rect 26065 36125 26099 36159
rect 26709 36125 26743 36159
rect 27905 36125 27939 36159
rect 31769 36125 31803 36159
rect 32229 36125 32263 36159
rect 35909 36125 35943 36159
rect 36737 36125 36771 36159
rect 37749 36125 37783 36159
rect 40049 36125 40083 36159
rect 40969 36125 41003 36159
rect 41429 36125 41463 36159
rect 42625 36125 42659 36159
rect 43637 36125 43671 36159
rect 44097 36125 44131 36159
rect 45937 36125 45971 36159
rect 46949 36125 46983 36159
rect 49341 36125 49375 36159
rect 50629 36125 50663 36159
rect 52009 36125 52043 36159
rect 53665 36125 53699 36159
rect 57989 36125 58023 36159
rect 59829 36125 59863 36159
rect 60657 36125 60691 36159
rect 61393 36125 61427 36159
rect 62865 36125 62899 36159
rect 64705 36125 64739 36159
rect 68385 36125 68419 36159
rect 69029 36125 69063 36159
rect 69673 36125 69707 36159
rect 74549 36125 74583 36159
rect 76113 36125 76147 36159
rect 77309 36125 77343 36159
rect 80069 36125 80103 36159
rect 81633 36125 81667 36159
rect 6929 36057 6963 36091
rect 19625 36057 19659 36091
rect 48605 36057 48639 36091
rect 48789 36057 48823 36091
rect 52745 36057 52779 36091
rect 52929 36057 52963 36091
rect 56977 36057 57011 36091
rect 57161 36057 57195 36091
rect 58909 36057 58943 36091
rect 59093 36057 59127 36091
rect 61761 36057 61795 36091
rect 63693 36057 63727 36091
rect 63877 36057 63911 36091
rect 65901 36057 65935 36091
rect 66085 36057 66119 36091
rect 77953 36057 77987 36091
rect 78505 36057 78539 36091
rect 95433 36057 95467 36091
rect 9229 35989 9263 36023
rect 20637 35989 20671 36023
rect 21373 35989 21407 36023
rect 26893 35989 26927 36023
rect 28641 35989 28675 36023
rect 32413 35989 32447 36023
rect 33149 35989 33183 36023
rect 35449 35989 35483 36023
rect 36553 35989 36587 36023
rect 38945 35989 38979 36023
rect 40233 35989 40267 36023
rect 45293 35989 45327 36023
rect 47133 35989 47167 36023
rect 51549 35989 51583 36023
rect 56425 35989 56459 36023
rect 58173 35989 58207 36023
rect 65165 35989 65199 36023
rect 75193 35989 75227 36023
rect 79149 35989 79183 36023
rect 81541 35989 81575 36023
rect 82001 35989 82035 36023
rect 83105 35989 83139 36023
rect 83657 35989 83691 36023
rect 84117 35989 84151 36023
rect 84761 35989 84795 36023
rect 85405 35989 85439 36023
rect 86417 35989 86451 36023
rect 89085 35989 89119 36023
rect 89637 35989 89671 36023
rect 90189 35989 90223 36023
rect 92857 35989 92891 36023
rect 94697 35989 94731 36023
rect 95893 35989 95927 36023
rect 97825 35989 97859 36023
rect 98377 35989 98411 36023
rect 100585 35989 100619 36023
rect 112177 35989 112211 36023
rect 112729 35989 112763 36023
rect 113465 35989 113499 36023
rect 114201 35989 114235 36023
rect 114753 35989 114787 36023
rect 121561 35989 121595 36023
rect 123125 35989 123159 36023
rect 19901 35785 19935 35819
rect 21097 35785 21131 35819
rect 25237 35785 25271 35819
rect 26617 35785 26651 35819
rect 28549 35785 28583 35819
rect 29193 35785 29227 35819
rect 31769 35785 31803 35819
rect 35265 35785 35299 35819
rect 36369 35785 36403 35819
rect 37657 35785 37691 35819
rect 38669 35785 38703 35819
rect 39313 35785 39347 35819
rect 42717 35785 42751 35819
rect 44005 35785 44039 35819
rect 45109 35785 45143 35819
rect 46121 35785 46155 35819
rect 46673 35785 46707 35819
rect 49157 35785 49191 35819
rect 50537 35785 50571 35819
rect 51273 35785 51307 35819
rect 52285 35785 52319 35819
rect 55045 35785 55079 35819
rect 57529 35785 57563 35819
rect 58173 35785 58207 35819
rect 59921 35785 59955 35819
rect 60381 35785 60415 35819
rect 61025 35785 61059 35819
rect 62681 35785 62715 35819
rect 64337 35785 64371 35819
rect 64889 35785 64923 35819
rect 66637 35785 66671 35819
rect 67281 35785 67315 35819
rect 68477 35785 68511 35819
rect 81173 35785 81207 35819
rect 81725 35785 81759 35819
rect 82369 35785 82403 35819
rect 83841 35785 83875 35819
rect 85221 35785 85255 35819
rect 34529 35717 34563 35751
rect 62129 35717 62163 35751
rect 63785 35649 63819 35683
rect 65349 35649 65383 35683
rect 65993 35649 66027 35683
rect 80437 35649 80471 35683
rect 80989 35649 81023 35683
rect 78965 35581 78999 35615
rect 25789 35513 25823 35547
rect 28089 35513 28123 35547
rect 35817 35513 35851 35547
rect 40877 35513 40911 35547
rect 59369 35513 59403 35547
rect 65533 35513 65567 35547
rect 24225 35445 24259 35479
rect 24777 35445 24811 35479
rect 30941 35445 30975 35479
rect 33149 35445 33183 35479
rect 36921 35445 36955 35479
rect 38117 35445 38151 35479
rect 39865 35445 39899 35479
rect 40417 35445 40451 35479
rect 41429 35445 41463 35479
rect 42073 35445 42107 35479
rect 43453 35445 43487 35479
rect 44465 35445 44499 35479
rect 47133 35445 47167 35479
rect 48145 35445 48179 35479
rect 48605 35445 48639 35479
rect 49893 35445 49927 35479
rect 51825 35445 51859 35479
rect 53113 35445 53147 35479
rect 54033 35445 54067 35479
rect 56057 35445 56091 35479
rect 56977 35445 57011 35479
rect 58725 35445 58759 35479
rect 61577 35445 61611 35479
rect 69213 35445 69247 35479
rect 69765 35445 69799 35479
rect 75101 35445 75135 35479
rect 79977 35445 80011 35479
rect 82921 35445 82955 35479
rect 84393 35445 84427 35479
rect 21005 35241 21039 35275
rect 24777 35241 24811 35275
rect 25973 35241 26007 35275
rect 28733 35241 28767 35275
rect 79517 35241 79551 35275
rect 80069 35241 80103 35275
rect 80621 35241 80655 35275
rect 81357 35241 81391 35275
rect 81817 35241 81851 35275
rect 82369 35241 82403 35275
rect 36001 35173 36035 35207
rect 37565 35173 37599 35207
rect 41705 35173 41739 35207
rect 43453 35173 43487 35207
rect 44189 35173 44223 35207
rect 58909 35105 58943 35139
rect 59921 35105 59955 35139
rect 62313 35105 62347 35139
rect 62957 35105 62991 35139
rect 64245 35105 64279 35139
rect 65901 35105 65935 35139
rect 69213 35105 69247 35139
rect 37013 35037 37047 35071
rect 65257 35037 65291 35071
rect 47685 34969 47719 35003
rect 48605 34969 48639 35003
rect 50353 34969 50387 35003
rect 51273 34969 51307 35003
rect 53849 34969 53883 35003
rect 25513 34901 25547 34935
rect 38853 34901 38887 34935
rect 40693 34901 40727 34935
rect 42809 34901 42843 34935
rect 45661 34901 45695 34935
rect 60749 34901 60783 34935
rect 61209 34901 61243 34935
rect 61853 34901 61887 34935
rect 63693 34901 63727 34935
rect 43821 34629 43855 34663
rect 64061 5865 64095 5899
rect 65809 5865 65843 5899
rect 80069 5865 80103 5899
rect 65165 5525 65199 5559
rect 69489 5525 69523 5559
rect 79057 5525 79091 5559
rect 79517 5525 79551 5559
rect 80621 5525 80655 5559
rect 28365 5321 28399 5355
rect 36093 5321 36127 5355
rect 38301 5321 38335 5355
rect 53481 5321 53515 5355
rect 63693 5321 63727 5355
rect 65993 5321 66027 5355
rect 69029 5321 69063 5355
rect 69673 5321 69707 5355
rect 78781 5321 78815 5355
rect 67097 5253 67131 5287
rect 79333 5185 79367 5219
rect 80161 5185 80195 5219
rect 80805 5185 80839 5219
rect 81449 5185 81483 5219
rect 36737 5049 36771 5083
rect 37565 5049 37599 5083
rect 60841 5049 60875 5083
rect 62589 5049 62623 5083
rect 66545 5049 66579 5083
rect 78137 5049 78171 5083
rect 82553 5049 82587 5083
rect 35633 4981 35667 5015
rect 42717 4981 42751 5015
rect 47133 4981 47167 5015
rect 48145 4981 48179 5015
rect 48605 4981 48639 5015
rect 49157 4981 49191 5015
rect 53021 4981 53055 5015
rect 58081 4981 58115 5015
rect 58725 4981 58759 5015
rect 61853 4981 61887 5015
rect 64337 4981 64371 5015
rect 64889 4981 64923 5015
rect 65349 4981 65383 5015
rect 68477 4981 68511 5015
rect 70133 4981 70167 5015
rect 70685 4981 70719 5015
rect 79425 4981 79459 5015
rect 79977 4981 80011 5015
rect 80621 4981 80655 5015
rect 81357 4981 81391 5015
rect 82001 4981 82035 5015
rect 83013 4981 83047 5015
rect 40601 4777 40635 4811
rect 45293 4777 45327 4811
rect 48329 4777 48363 4811
rect 48973 4777 49007 4811
rect 49525 4777 49559 4811
rect 53849 4777 53883 4811
rect 57989 4777 58023 4811
rect 59093 4777 59127 4811
rect 61117 4777 61151 4811
rect 67649 4777 67683 4811
rect 68201 4777 68235 4811
rect 78229 4777 78263 4811
rect 83105 4777 83139 4811
rect 43453 4709 43487 4743
rect 66085 4709 66119 4743
rect 66729 4709 66763 4743
rect 80621 4709 80655 4743
rect 33701 4641 33735 4675
rect 34345 4641 34379 4675
rect 47501 4641 47535 4675
rect 47593 4641 47627 4675
rect 62957 4641 62991 4675
rect 79793 4641 79827 4675
rect 28181 4573 28215 4607
rect 29101 4573 29135 4607
rect 35357 4573 35391 4607
rect 35817 4573 35851 4607
rect 38025 4573 38059 4607
rect 40049 4573 40083 4607
rect 41981 4573 42015 4607
rect 42441 4573 42475 4607
rect 47409 4573 47443 4607
rect 51641 4573 51675 4607
rect 57069 4573 57103 4607
rect 62221 4573 62255 4607
rect 65073 4573 65107 4607
rect 69857 4573 69891 4607
rect 70961 4573 70995 4607
rect 79701 4573 79735 4607
rect 80437 4573 80471 4607
rect 81449 4573 81483 4607
rect 82093 4573 82127 4607
rect 29745 4505 29779 4539
rect 36829 4505 36863 4539
rect 48421 4505 48455 4539
rect 58449 4505 58483 4539
rect 64153 4505 64187 4539
rect 71513 4505 71547 4539
rect 82645 4505 82679 4539
rect 6377 4437 6411 4471
rect 22661 4437 22695 4471
rect 23857 4437 23891 4471
rect 27629 4437 27663 4471
rect 30389 4437 30423 4471
rect 31953 4437 31987 4471
rect 32781 4437 32815 4471
rect 35909 4437 35943 4471
rect 37289 4437 37323 4471
rect 38761 4437 38795 4471
rect 39497 4437 39531 4471
rect 41245 4437 41279 4471
rect 42533 4437 42567 4471
rect 46489 4437 46523 4471
rect 47041 4437 47075 4471
rect 50445 4437 50479 4471
rect 51733 4437 51767 4471
rect 52745 4437 52779 4471
rect 54309 4437 54343 4471
rect 56057 4437 56091 4471
rect 56609 4437 56643 4471
rect 57253 4437 57287 4471
rect 61669 4437 61703 4471
rect 62313 4437 62347 4471
rect 63509 4437 63543 4471
rect 64429 4437 64463 4471
rect 65257 4437 65291 4471
rect 68661 4437 68695 4471
rect 69213 4437 69247 4471
rect 70041 4437 70075 4471
rect 75009 4437 75043 4471
rect 77677 4437 77711 4471
rect 78689 4437 78723 4471
rect 79241 4437 79275 4471
rect 79609 4437 79643 4471
rect 81357 4437 81391 4471
rect 81909 4437 81943 4471
rect 83657 4437 83691 4471
rect 67189 4233 67223 4267
rect 81449 4233 81483 4267
rect 81817 4233 81851 4267
rect 26617 4165 26651 4199
rect 35817 4165 35851 4199
rect 37565 4165 37599 4199
rect 44281 4165 44315 4199
rect 48145 4165 48179 4199
rect 53021 4165 53055 4199
rect 56517 4165 56551 4199
rect 64705 4165 64739 4199
rect 79425 4165 79459 4199
rect 6561 4097 6595 4131
rect 22477 4097 22511 4131
rect 23581 4097 23615 4131
rect 27353 4097 27387 4131
rect 27997 4097 28031 4131
rect 29009 4097 29043 4131
rect 32781 4097 32815 4131
rect 33241 4097 33275 4131
rect 34069 4097 34103 4131
rect 34989 4097 35023 4131
rect 36001 4097 36035 4131
rect 36461 4097 36495 4131
rect 37749 4097 37783 4131
rect 38209 4097 38243 4131
rect 39405 4097 39439 4131
rect 39865 4097 39899 4131
rect 42073 4097 42107 4131
rect 42993 4097 43027 4131
rect 44465 4097 44499 4131
rect 46305 4097 46339 4131
rect 47041 4097 47075 4131
rect 48237 4097 48271 4131
rect 49065 4097 49099 4131
rect 49617 4097 49651 4131
rect 49801 4097 49835 4131
rect 51089 4097 51123 4131
rect 51733 4097 51767 4131
rect 52377 4097 52411 4131
rect 53205 4097 53239 4131
rect 55137 4097 55171 4131
rect 55873 4097 55907 4131
rect 56701 4097 56735 4131
rect 57345 4097 57379 4131
rect 58081 4097 58115 4131
rect 60105 4097 60139 4131
rect 60657 4097 60691 4131
rect 60841 4097 60875 4131
rect 61485 4097 61519 4131
rect 62313 4097 62347 4131
rect 63325 4097 63359 4131
rect 65717 4097 65751 4131
rect 66545 4097 66579 4131
rect 68753 4097 68787 4131
rect 71789 4097 71823 4131
rect 75745 4097 75779 4131
rect 77953 4097 77987 4131
rect 81909 4097 81943 4131
rect 83841 4097 83875 4131
rect 29653 4029 29687 4063
rect 48329 4029 48363 4063
rect 64429 4029 64463 4063
rect 64613 4029 64647 4063
rect 69397 4029 69431 4063
rect 69673 4029 69707 4063
rect 72341 4029 72375 4063
rect 79149 4029 79183 4063
rect 82001 4029 82035 4063
rect 83197 4029 83231 4063
rect 7205 3961 7239 3995
rect 24685 3961 24719 3995
rect 28549 3961 28583 3995
rect 41429 3961 41463 3995
rect 58173 3961 58207 3995
rect 62405 3961 62439 3995
rect 65073 3961 65107 3995
rect 68937 3961 68971 3995
rect 73537 3961 73571 3995
rect 77125 3961 77159 3995
rect 80897 3961 80931 3995
rect 82737 3961 82771 3995
rect 6009 3893 6043 3927
rect 6745 3893 6779 3927
rect 8033 3893 8067 3927
rect 22293 3893 22327 3927
rect 23397 3893 23431 3927
rect 24133 3893 24167 3927
rect 25973 3893 26007 3927
rect 27169 3893 27203 3927
rect 27905 3893 27939 3927
rect 30481 3893 30515 3927
rect 31677 3893 31711 3927
rect 33333 3893 33367 3927
rect 33885 3893 33919 3927
rect 35173 3893 35207 3927
rect 36645 3893 36679 3927
rect 38301 3893 38335 3927
rect 39221 3893 39255 3927
rect 39957 3893 39991 3927
rect 40877 3893 40911 3927
rect 41889 3893 41923 3927
rect 42809 3893 42843 3927
rect 43729 3893 43763 3927
rect 45109 3893 45143 3927
rect 45569 3893 45603 3927
rect 46213 3893 46247 3927
rect 46857 3893 46891 3927
rect 47777 3893 47811 3927
rect 50445 3893 50479 3927
rect 50905 3893 50939 3927
rect 51549 3893 51583 3927
rect 52285 3893 52319 3927
rect 54033 3893 54067 3927
rect 54585 3893 54619 3927
rect 55229 3893 55263 3927
rect 57161 3893 57195 3927
rect 59185 3893 59219 3927
rect 61393 3893 61427 3927
rect 63509 3893 63543 3927
rect 65533 3893 65567 3927
rect 66453 3893 66487 3927
rect 67833 3893 67867 3927
rect 71145 3893 71179 3927
rect 74641 3893 74675 3927
rect 76573 3893 76607 3927
rect 78137 3893 78171 3927
rect 84393 3893 84427 3927
rect 8585 3689 8619 3723
rect 22753 3689 22787 3723
rect 23949 3689 23983 3723
rect 24685 3689 24719 3723
rect 30205 3689 30239 3723
rect 33149 3689 33183 3723
rect 40233 3689 40267 3723
rect 40969 3689 41003 3723
rect 43821 3689 43855 3723
rect 51917 3689 51951 3723
rect 57437 3689 57471 3723
rect 65257 3689 65291 3723
rect 68845 3689 68879 3723
rect 70041 3689 70075 3723
rect 81265 3689 81299 3723
rect 82461 3689 82495 3723
rect 84761 3689 84795 3723
rect 29009 3621 29043 3655
rect 36921 3621 36955 3655
rect 43361 3621 43395 3655
rect 53941 3621 53975 3655
rect 63325 3621 63359 3655
rect 23397 3553 23431 3587
rect 26249 3553 26283 3587
rect 26525 3553 26559 3587
rect 35725 3553 35759 3587
rect 35817 3553 35851 3587
rect 41613 3553 41647 3587
rect 41889 3553 41923 3587
rect 44281 3553 44315 3587
rect 44373 3553 44407 3587
rect 52377 3553 52411 3587
rect 52561 3553 52595 3587
rect 56425 3553 56459 3587
rect 56517 3553 56551 3587
rect 57989 3553 58023 3587
rect 61117 3553 61151 3587
rect 61209 3553 61243 3587
rect 63785 3553 63819 3587
rect 63877 3553 63911 3587
rect 64613 3553 64647 3587
rect 64797 3553 64831 3587
rect 66453 3553 66487 3587
rect 68293 3553 68327 3587
rect 69397 3553 69431 3587
rect 71421 3553 71455 3587
rect 71605 3553 71639 3587
rect 75377 3553 75411 3587
rect 77861 3553 77895 3587
rect 78505 3553 78539 3587
rect 78781 3553 78815 3587
rect 80253 3553 80287 3587
rect 81909 3553 81943 3587
rect 83013 3553 83047 3587
rect 4905 3485 4939 3519
rect 5365 3485 5399 3519
rect 6285 3485 6319 3519
rect 6929 3485 6963 3519
rect 8033 3485 8067 3519
rect 21465 3485 21499 3519
rect 22109 3485 22143 3519
rect 28825 3485 28859 3519
rect 30757 3485 30791 3519
rect 34161 3485 34195 3519
rect 38669 3485 38703 3519
rect 45201 3485 45235 3519
rect 46213 3485 46247 3519
rect 46859 3485 46893 3519
rect 49065 3485 49099 3519
rect 49341 3485 49375 3519
rect 50905 3485 50939 3519
rect 52285 3485 52319 3519
rect 54953 3485 54987 3519
rect 59185 3485 59219 3519
rect 60105 3485 60139 3519
rect 62037 3485 62071 3519
rect 62497 3485 62531 3519
rect 63693 3485 63727 3519
rect 64889 3485 64923 3519
rect 66269 3485 66303 3519
rect 67373 3485 67407 3519
rect 68385 3485 68419 3519
rect 68477 3485 68511 3519
rect 69581 3485 69615 3519
rect 69673 3485 69707 3519
rect 73537 3485 73571 3519
rect 74089 3485 74123 3519
rect 74181 3485 74215 3519
rect 75285 3485 75319 3519
rect 76113 3485 76147 3519
rect 76849 3485 76883 3519
rect 77769 3485 77803 3519
rect 81633 3485 81667 3519
rect 82921 3485 82955 3519
rect 6193 3417 6227 3451
rect 31953 3417 31987 3451
rect 33057 3417 33091 3451
rect 35633 3417 35667 3451
rect 38209 3417 38243 3451
rect 40141 3417 40175 3451
rect 41061 3417 41095 3451
rect 44189 3417 44223 3451
rect 53205 3417 53239 3451
rect 53757 3417 53791 3451
rect 57897 3417 57931 3451
rect 61025 3417 61059 3451
rect 81725 3417 81759 3451
rect 84209 3417 84243 3451
rect 5549 3349 5583 3383
rect 6745 3349 6779 3383
rect 7941 3349 7975 3383
rect 9229 3349 9263 3383
rect 20453 3349 20487 3383
rect 21005 3349 21039 3383
rect 21649 3349 21683 3383
rect 22201 3349 22235 3383
rect 23121 3349 23155 3383
rect 23213 3349 23247 3383
rect 25145 3349 25179 3383
rect 25789 3349 25823 3383
rect 27997 3349 28031 3383
rect 30849 3349 30883 3383
rect 32413 3349 32447 3383
rect 34345 3349 34379 3383
rect 35265 3349 35299 3383
rect 38853 3349 38887 3383
rect 39497 3349 39531 3383
rect 45293 3349 45327 3383
rect 46397 3349 46431 3383
rect 48145 3349 48179 3383
rect 50353 3349 50387 3383
rect 51089 3349 51123 3383
rect 54769 3349 54803 3383
rect 55965 3349 55999 3383
rect 56333 3349 56367 3383
rect 57805 3349 57839 3383
rect 58725 3349 58759 3383
rect 59369 3349 59403 3383
rect 59921 3349 59955 3383
rect 60657 3349 60691 3383
rect 61853 3349 61887 3383
rect 62681 3349 62715 3383
rect 67281 3349 67315 3383
rect 70961 3349 70995 3383
rect 71329 3349 71363 3383
rect 72249 3349 72283 3383
rect 72985 3349 73019 3383
rect 74825 3349 74859 3383
rect 75193 3349 75227 3383
rect 76665 3349 76699 3383
rect 77309 3349 77343 3383
rect 77677 3349 77711 3383
rect 82829 3349 82863 3383
rect 83657 3349 83691 3383
rect 85405 3349 85439 3383
rect 5733 3145 5767 3179
rect 5825 3145 5859 3179
rect 8125 3145 8159 3179
rect 9413 3145 9447 3179
rect 24225 3145 24259 3179
rect 24685 3145 24719 3179
rect 27353 3145 27387 3179
rect 27721 3145 27755 3179
rect 28549 3145 28583 3179
rect 29009 3145 29043 3179
rect 30849 3145 30883 3179
rect 33793 3145 33827 3179
rect 34161 3145 34195 3179
rect 34253 3145 34287 3179
rect 37473 3145 37507 3179
rect 37933 3145 37967 3179
rect 45017 3145 45051 3179
rect 57345 3145 57379 3179
rect 68937 3145 68971 3179
rect 71881 3145 71915 3179
rect 73721 3145 73755 3179
rect 77217 3145 77251 3179
rect 78045 3145 78079 3179
rect 81725 3145 81759 3179
rect 82185 3145 82219 3179
rect 83013 3145 83047 3179
rect 145941 3145 145975 3179
rect 5273 3077 5307 3111
rect 6009 3077 6043 3111
rect 21373 3077 21407 3111
rect 23489 3077 23523 3111
rect 27813 3077 27847 3111
rect 28917 3077 28951 3111
rect 29837 3077 29871 3111
rect 30757 3077 30791 3111
rect 31493 3077 31527 3111
rect 31677 3077 31711 3111
rect 32413 3077 32447 3111
rect 36921 3077 36955 3111
rect 39221 3077 39255 3111
rect 41613 3077 41647 3111
rect 41705 3077 41739 3111
rect 45937 3077 45971 3111
rect 47777 3077 47811 3111
rect 49525 3077 49559 3111
rect 50905 3077 50939 3111
rect 53297 3077 53331 3111
rect 53389 3077 53423 3111
rect 54585 3077 54619 3111
rect 57437 3077 57471 3111
rect 58541 3077 58575 3111
rect 60013 3077 60047 3111
rect 62221 3077 62255 3111
rect 63693 3077 63727 3111
rect 64613 3077 64647 3111
rect 64797 3077 64831 3111
rect 65533 3077 65567 3111
rect 70409 3077 70443 3111
rect 78689 3077 78723 3111
rect 84577 3077 84611 3111
rect 6745 3009 6779 3043
rect 7021 3009 7055 3043
rect 8309 3009 8343 3043
rect 9229 3009 9263 3043
rect 9413 3009 9447 3043
rect 20821 3009 20855 3043
rect 21281 3009 21315 3043
rect 23765 3009 23799 3043
rect 24593 3009 24627 3043
rect 25789 3009 25823 3043
rect 26433 3009 26467 3043
rect 32873 3009 32907 3043
rect 37841 3009 37875 3043
rect 38945 3009 38979 3043
rect 42717 3009 42751 3043
rect 43729 3009 43763 3043
rect 46121 3009 46155 3043
rect 46765 3009 46799 3043
rect 50169 3009 50203 3043
rect 50629 3009 50663 3043
rect 54309 3009 54343 3043
rect 56609 3009 56643 3043
rect 58449 3009 58483 3043
rect 59737 3009 59771 3043
rect 61945 3009 61979 3043
rect 63601 3009 63635 3043
rect 65257 3009 65291 3043
rect 67557 3009 67591 3043
rect 68845 3009 68879 3043
rect 69489 3009 69523 3043
rect 70133 3009 70167 3043
rect 72433 3009 72467 3043
rect 73629 3009 73663 3043
rect 74457 3009 74491 3043
rect 75101 3009 75135 3043
rect 75745 3009 75779 3043
rect 77309 3009 77343 3043
rect 77861 3009 77895 3043
rect 81265 3009 81299 3043
rect 82093 3009 82127 3043
rect 83105 3009 83139 3043
rect 84025 3009 84059 3043
rect 86141 3009 86175 3043
rect 104541 3009 104575 3043
rect 20269 2941 20303 2975
rect 22017 2941 22051 2975
rect 24777 2941 24811 2975
rect 27905 2941 27939 2975
rect 29101 2941 29135 2975
rect 30113 2941 30147 2975
rect 33149 2941 33183 2975
rect 34437 2941 34471 2975
rect 35173 2941 35207 2975
rect 38025 2941 38059 2975
rect 41429 2941 41463 2975
rect 52377 2941 52411 2975
rect 53573 2941 53607 2975
rect 58633 2941 58667 2975
rect 61485 2941 61519 2975
rect 63877 2941 63911 2975
rect 79241 2941 79275 2975
rect 79517 2941 79551 2975
rect 82277 2941 82311 2975
rect 85037 2941 85071 2975
rect 5273 2873 5307 2907
rect 52929 2873 52963 2907
rect 58081 2873 58115 2907
rect 63233 2873 63267 2907
rect 72617 2873 72651 2907
rect 75193 2873 75227 2907
rect 4721 2805 4755 2839
rect 15025 2805 15059 2839
rect 25973 2805 26007 2839
rect 26525 2805 26559 2839
rect 40693 2805 40727 2839
rect 42073 2805 42107 2839
rect 43177 2805 43211 2839
rect 46949 2805 46983 2839
rect 50077 2805 50111 2839
rect 56057 2805 56091 2839
rect 56701 2805 56735 2839
rect 67005 2805 67039 2839
rect 67741 2805 67775 2839
rect 69673 2805 69707 2839
rect 74273 2805 74307 2839
rect 75929 2805 75963 2839
rect 76481 2805 76515 2839
rect 83933 2805 83967 2839
rect 85681 2805 85715 2839
rect 97733 2805 97767 2839
rect 101873 2805 101907 2839
rect 110245 2805 110279 2839
rect 118433 2805 118467 2839
rect 122573 2805 122607 2839
rect 125333 2805 125367 2839
rect 130853 2805 130887 2839
rect 143273 2805 143307 2839
rect 4261 2601 4295 2635
rect 9505 2601 9539 2635
rect 14473 2601 14507 2635
rect 15393 2601 15427 2635
rect 21281 2601 21315 2635
rect 24777 2601 24811 2635
rect 25697 2601 25731 2635
rect 26525 2601 26559 2635
rect 28917 2601 28951 2635
rect 34069 2601 34103 2635
rect 36645 2601 36679 2635
rect 39221 2601 39255 2635
rect 40049 2601 40083 2635
rect 41337 2601 41371 2635
rect 44373 2601 44407 2635
rect 47225 2601 47259 2635
rect 49525 2601 49559 2635
rect 62681 2601 62715 2635
rect 64981 2601 65015 2635
rect 69029 2601 69063 2635
rect 85497 2601 85531 2635
rect 89729 2601 89763 2635
rect 94329 2601 94363 2635
rect 98009 2601 98043 2635
rect 102149 2601 102183 2635
rect 106289 2601 106323 2635
rect 110521 2601 110555 2635
rect 114937 2601 114971 2635
rect 118709 2601 118743 2635
rect 122849 2601 122883 2635
rect 126989 2601 127023 2635
rect 131129 2601 131163 2635
rect 137293 2601 137327 2635
rect 139409 2601 139443 2635
rect 143549 2601 143583 2635
rect 147321 2601 147355 2635
rect 19717 2533 19751 2567
rect 20729 2533 20763 2567
rect 52377 2533 52411 2567
rect 53573 2533 53607 2567
rect 69673 2533 69707 2567
rect 109785 2533 109819 2567
rect 129565 2533 129599 2567
rect 135545 2533 135579 2567
rect 6009 2465 6043 2499
rect 6561 2465 6595 2499
rect 22017 2465 22051 2499
rect 27169 2465 27203 2499
rect 29929 2465 29963 2499
rect 32321 2465 32355 2499
rect 34897 2465 34931 2499
rect 37473 2465 37507 2499
rect 40601 2465 40635 2499
rect 42625 2465 42659 2499
rect 45477 2465 45511 2499
rect 45753 2465 45787 2499
rect 47777 2465 47811 2499
rect 50629 2465 50663 2499
rect 50905 2465 50939 2499
rect 54217 2465 54251 2499
rect 55689 2465 55723 2499
rect 58081 2465 58115 2499
rect 60933 2465 60967 2499
rect 63233 2465 63267 2499
rect 65809 2465 65843 2499
rect 70961 2465 70995 2499
rect 73537 2465 73571 2499
rect 76113 2465 76147 2499
rect 78689 2465 78723 2499
rect 78965 2465 78999 2499
rect 81265 2465 81299 2499
rect 86509 2465 86543 2499
rect 120733 2465 120767 2499
rect 2881 2397 2915 2431
rect 9689 2397 9723 2431
rect 10149 2397 10183 2431
rect 12541 2397 12575 2431
rect 15209 2397 15243 2431
rect 18061 2397 18095 2431
rect 21465 2397 21499 2431
rect 30297 2397 30331 2431
rect 31769 2397 31803 2431
rect 40417 2397 40451 2431
rect 41797 2397 41831 2431
rect 53389 2397 53423 2431
rect 54493 2397 54527 2431
rect 69581 2397 69615 2431
rect 70225 2397 70259 2431
rect 75561 2397 75595 2431
rect 84301 2397 84335 2431
rect 84945 2397 84979 2431
rect 88165 2397 88199 2431
rect 92305 2397 92339 2431
rect 96721 2397 96755 2431
rect 100585 2397 100619 2431
rect 104725 2397 104759 2431
rect 109601 2397 109635 2431
rect 113005 2397 113039 2431
rect 117329 2397 117363 2431
rect 121285 2397 121319 2431
rect 125425 2397 125459 2431
rect 130209 2397 130243 2431
rect 133153 2397 133187 2431
rect 133705 2397 133739 2431
rect 135361 2397 135395 2431
rect 137937 2397 137971 2431
rect 138765 2397 138799 2431
rect 139225 2397 139259 2431
rect 141985 2397 142019 2431
rect 146125 2397 146159 2431
rect 5733 2329 5767 2363
rect 6837 2329 6871 2363
rect 8585 2329 8619 2363
rect 14381 2329 14415 2363
rect 19533 2329 19567 2363
rect 20545 2329 20579 2363
rect 22293 2329 22327 2363
rect 24869 2329 24903 2363
rect 25789 2329 25823 2363
rect 26433 2329 26467 2363
rect 27445 2329 27479 2363
rect 32597 2329 32631 2363
rect 35173 2329 35207 2363
rect 37749 2329 37783 2363
rect 40509 2329 40543 2363
rect 42901 2329 42935 2363
rect 48053 2329 48087 2363
rect 55965 2329 55999 2363
rect 58357 2329 58391 2363
rect 61209 2329 61243 2363
rect 63509 2329 63543 2363
rect 66085 2329 66119 2363
rect 68937 2329 68971 2363
rect 71237 2329 71271 2363
rect 73813 2329 73847 2363
rect 76389 2329 76423 2363
rect 78137 2329 78171 2363
rect 80713 2329 80747 2363
rect 81541 2329 81575 2363
rect 84853 2329 84887 2363
rect 85589 2329 85623 2363
rect 86969 2329 87003 2363
rect 89085 2329 89119 2363
rect 89637 2329 89671 2363
rect 94237 2329 94271 2363
rect 97917 2329 97951 2363
rect 102057 2329 102091 2363
rect 105645 2329 105679 2363
rect 106197 2329 106231 2363
rect 110429 2329 110463 2363
rect 114845 2329 114879 2363
rect 118617 2329 118651 2363
rect 122757 2329 122791 2363
rect 126345 2329 126379 2363
rect 126897 2329 126931 2363
rect 131037 2329 131071 2363
rect 143457 2329 143491 2363
rect 147597 2329 147631 2363
rect 148241 2329 148275 2363
rect 2697 2261 2731 2295
rect 3433 2261 3467 2295
rect 12357 2261 12391 2295
rect 13645 2261 13679 2295
rect 17877 2261 17911 2295
rect 18889 2261 18923 2295
rect 23765 2261 23799 2295
rect 41981 2261 42015 2295
rect 57437 2261 57471 2295
rect 59829 2261 59863 2295
rect 67557 2261 67591 2295
rect 70317 2261 70351 2295
rect 72709 2261 72743 2295
rect 83013 2261 83047 2295
rect 84117 2261 84151 2295
rect 87613 2261 87647 2295
rect 88349 2261 88383 2295
rect 91753 2261 91787 2295
rect 92489 2261 92523 2295
rect 93593 2261 93627 2295
rect 96077 2261 96111 2295
rect 96905 2261 96939 2295
rect 100033 2261 100067 2295
rect 100769 2261 100803 2295
rect 104909 2261 104943 2295
rect 109049 2261 109083 2295
rect 112453 2261 112487 2295
rect 113189 2261 113223 2295
rect 114201 2261 114235 2295
rect 116685 2261 116719 2295
rect 117513 2261 117547 2295
rect 121469 2261 121503 2295
rect 125609 2261 125643 2295
rect 130393 2261 130427 2295
rect 133889 2261 133923 2295
rect 134809 2261 134843 2295
rect 138121 2261 138155 2295
rect 141433 2261 141467 2295
rect 142169 2261 142203 2295
rect 146309 2261 146343 2295
<< metal1 >>
rect 42610 39312 42616 39364
rect 42668 39352 42674 39364
rect 73614 39352 73620 39364
rect 42668 39324 73620 39352
rect 42668 39312 42674 39324
rect 73614 39312 73620 39324
rect 73672 39312 73678 39364
rect 39390 39244 39396 39296
rect 39448 39284 39454 39296
rect 68646 39284 68652 39296
rect 39448 39256 68652 39284
rect 39448 39244 39454 39256
rect 68646 39244 68652 39256
rect 68704 39244 68710 39296
rect 84930 39284 84936 39296
rect 70366 39256 84936 39284
rect 46290 39176 46296 39228
rect 46348 39216 46354 39228
rect 70366 39216 70394 39256
rect 84930 39244 84936 39256
rect 84988 39244 84994 39296
rect 83826 39216 83832 39228
rect 46348 39188 70394 39216
rect 73632 39188 83832 39216
rect 46348 39176 46354 39188
rect 22186 39108 22192 39160
rect 22244 39148 22250 39160
rect 73632 39148 73660 39188
rect 83826 39176 83832 39188
rect 83884 39176 83890 39228
rect 22244 39120 73660 39148
rect 22244 39108 22250 39120
rect 75178 39108 75184 39160
rect 75236 39148 75242 39160
rect 85298 39148 85304 39160
rect 75236 39120 85304 39148
rect 75236 39108 75242 39120
rect 85298 39108 85304 39120
rect 85356 39108 85362 39160
rect 63494 39040 63500 39092
rect 63552 39080 63558 39092
rect 118050 39080 118056 39092
rect 63552 39052 118056 39080
rect 63552 39040 63558 39052
rect 118050 39040 118056 39052
rect 118108 39040 118114 39092
rect 43990 38972 43996 39024
rect 44048 39012 44054 39024
rect 82078 39012 82084 39024
rect 44048 38984 82084 39012
rect 44048 38972 44054 38984
rect 82078 38972 82084 38984
rect 82136 38972 82142 39024
rect 46934 38904 46940 38956
rect 46992 38944 46998 38956
rect 89806 38944 89812 38956
rect 46992 38916 89812 38944
rect 46992 38904 46998 38916
rect 89806 38904 89812 38916
rect 89864 38904 89870 38956
rect 49786 38836 49792 38888
rect 49844 38876 49850 38888
rect 93026 38876 93032 38888
rect 49844 38848 93032 38876
rect 49844 38836 49850 38848
rect 93026 38836 93032 38848
rect 93084 38836 93090 38888
rect 95050 38836 95056 38888
rect 95108 38876 95114 38888
rect 123110 38876 123116 38888
rect 95108 38848 123116 38876
rect 95108 38836 95114 38848
rect 123110 38836 123116 38848
rect 123168 38836 123174 38888
rect 35526 38768 35532 38820
rect 35584 38808 35590 38820
rect 94222 38808 94228 38820
rect 35584 38780 94228 38808
rect 35584 38768 35590 38780
rect 94222 38768 94228 38780
rect 94280 38768 94286 38820
rect 54938 38700 54944 38752
rect 54996 38740 55002 38752
rect 105262 38740 105268 38752
rect 54996 38712 105268 38740
rect 54996 38700 55002 38712
rect 105262 38700 105268 38712
rect 105320 38700 105326 38752
rect 59906 38632 59912 38684
rect 59964 38672 59970 38684
rect 113726 38672 113732 38684
rect 59964 38644 113732 38672
rect 59964 38632 59970 38644
rect 113726 38632 113732 38644
rect 113784 38632 113790 38684
rect 60090 38564 60096 38616
rect 60148 38604 60154 38616
rect 117866 38604 117872 38616
rect 60148 38576 117872 38604
rect 60148 38564 60154 38576
rect 117866 38564 117872 38576
rect 117924 38564 117930 38616
rect 61286 38496 61292 38548
rect 61344 38536 61350 38548
rect 120074 38536 120080 38548
rect 61344 38508 120080 38536
rect 61344 38496 61350 38508
rect 120074 38496 120080 38508
rect 120132 38496 120138 38548
rect 62850 38428 62856 38480
rect 62908 38468 62914 38480
rect 122558 38468 122564 38480
rect 62908 38440 122564 38468
rect 62908 38428 62914 38440
rect 122558 38428 122564 38440
rect 122616 38428 122622 38480
rect 53190 38360 53196 38412
rect 53248 38400 53254 38412
rect 112990 38400 112996 38412
rect 53248 38372 112996 38400
rect 53248 38360 53254 38372
rect 112990 38360 112996 38372
rect 113048 38360 113054 38412
rect 64690 38292 64696 38344
rect 64748 38332 64754 38344
rect 126514 38332 126520 38344
rect 64748 38304 126520 38332
rect 64748 38292 64754 38304
rect 126514 38292 126520 38304
rect 126572 38292 126578 38344
rect 48038 38224 48044 38276
rect 48096 38264 48102 38276
rect 111242 38264 111248 38276
rect 48096 38236 111248 38264
rect 48096 38224 48102 38236
rect 111242 38224 111248 38236
rect 111300 38224 111306 38276
rect 58526 38156 58532 38208
rect 58584 38196 58590 38208
rect 121454 38196 121460 38208
rect 58584 38168 121460 38196
rect 58584 38156 58590 38168
rect 121454 38156 121460 38168
rect 121512 38156 121518 38208
rect 66530 38088 66536 38140
rect 66588 38128 66594 38140
rect 130286 38128 130292 38140
rect 66588 38100 130292 38128
rect 66588 38088 66594 38100
rect 130286 38088 130292 38100
rect 130344 38088 130350 38140
rect 58710 38020 58716 38072
rect 58768 38060 58774 38072
rect 125870 38060 125876 38072
rect 58768 38032 125876 38060
rect 58768 38020 58774 38032
rect 125870 38020 125876 38032
rect 125928 38020 125934 38072
rect 51166 37952 51172 38004
rect 51224 37992 51230 38004
rect 97534 37992 97540 38004
rect 51224 37964 97540 37992
rect 51224 37952 51230 37964
rect 97534 37952 97540 37964
rect 97592 37952 97598 38004
rect 54294 37884 54300 37936
rect 54352 37924 54358 37936
rect 101950 37924 101956 37936
rect 54352 37896 101956 37924
rect 54352 37884 54358 37896
rect 101950 37884 101956 37896
rect 102008 37884 102014 37936
rect 33594 37816 33600 37868
rect 33652 37856 33658 37868
rect 75178 37856 75184 37868
rect 33652 37828 75184 37856
rect 33652 37816 33658 37828
rect 75178 37816 75184 37828
rect 75236 37816 75242 37868
rect 75914 37816 75920 37868
rect 75972 37856 75978 37868
rect 79318 37856 79324 37868
rect 75972 37828 79324 37856
rect 75972 37816 75978 37828
rect 79318 37816 79324 37828
rect 79376 37816 79382 37868
rect 80238 37816 80244 37868
rect 80296 37856 80302 37868
rect 83182 37856 83188 37868
rect 80296 37828 83188 37856
rect 80296 37816 80302 37828
rect 83182 37816 83188 37828
rect 83240 37816 83246 37868
rect 99466 37816 99472 37868
rect 99524 37856 99530 37868
rect 124950 37856 124956 37868
rect 99524 37828 124956 37856
rect 99524 37816 99530 37828
rect 124950 37816 124956 37828
rect 125008 37816 125014 37868
rect 45370 37748 45376 37800
rect 45428 37788 45434 37800
rect 62666 37788 62672 37800
rect 45428 37760 62672 37788
rect 45428 37748 45434 37760
rect 62666 37748 62672 37760
rect 62724 37748 62730 37800
rect 64414 37748 64420 37800
rect 64472 37788 64478 37800
rect 116210 37788 116216 37800
rect 64472 37760 116216 37788
rect 64472 37748 64478 37760
rect 116210 37748 116216 37760
rect 116268 37748 116274 37800
rect 40034 37680 40040 37732
rect 40092 37720 40098 37732
rect 67542 37720 67548 37732
rect 40092 37692 67548 37720
rect 40092 37680 40098 37692
rect 67542 37680 67548 37692
rect 67600 37680 67606 37732
rect 68370 37680 68376 37732
rect 68428 37720 68434 37732
rect 120626 37720 120632 37732
rect 68428 37692 120632 37720
rect 68428 37680 68434 37692
rect 120626 37680 120632 37692
rect 120684 37680 120690 37732
rect 19426 37612 19432 37664
rect 19484 37652 19490 37664
rect 25130 37652 25136 37664
rect 19484 37624 25136 37652
rect 19484 37612 19490 37624
rect 25130 37612 25136 37624
rect 25188 37612 25194 37664
rect 29086 37612 29092 37664
rect 29144 37652 29150 37664
rect 31018 37652 31024 37664
rect 29144 37624 31024 37652
rect 29144 37612 29150 37624
rect 31018 37612 31024 37624
rect 31076 37612 31082 37664
rect 33410 37612 33416 37664
rect 33468 37652 33474 37664
rect 53558 37652 53564 37664
rect 33468 37624 53564 37652
rect 33468 37612 33474 37624
rect 53558 37612 53564 37624
rect 53616 37612 53622 37664
rect 55214 37612 55220 37664
rect 55272 37652 55278 37664
rect 56134 37652 56140 37664
rect 55272 37624 56140 37652
rect 55272 37612 55278 37624
rect 56134 37612 56140 37624
rect 56192 37652 56198 37664
rect 110230 37652 110236 37664
rect 56192 37624 110236 37652
rect 56192 37612 56198 37624
rect 110230 37612 110236 37624
rect 110288 37612 110294 37664
rect 119890 37612 119896 37664
rect 119948 37652 119954 37664
rect 126422 37652 126428 37664
rect 119948 37624 126428 37652
rect 119948 37612 119954 37624
rect 126422 37612 126428 37624
rect 126480 37612 126486 37664
rect 1104 37562 148856 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 65654 37562
rect 65706 37510 65718 37562
rect 65770 37510 65782 37562
rect 65834 37510 65846 37562
rect 65898 37510 65910 37562
rect 65962 37510 96374 37562
rect 96426 37510 96438 37562
rect 96490 37510 96502 37562
rect 96554 37510 96566 37562
rect 96618 37510 96630 37562
rect 96682 37510 127094 37562
rect 127146 37510 127158 37562
rect 127210 37510 127222 37562
rect 127274 37510 127286 37562
rect 127338 37510 127350 37562
rect 127402 37510 148856 37562
rect 1104 37488 148856 37510
rect 2774 37448 2780 37460
rect 2735 37420 2780 37448
rect 2774 37408 2780 37420
rect 2832 37408 2838 37460
rect 6886 37420 30972 37448
rect 4522 37340 4528 37392
rect 4580 37380 4586 37392
rect 6886 37380 6914 37420
rect 29086 37380 29092 37392
rect 4580 37352 6914 37380
rect 22388 37352 29092 37380
rect 4580 37340 4586 37352
rect 4890 37244 4896 37256
rect 4851 37216 4896 37244
rect 4890 37204 4896 37216
rect 4948 37204 4954 37256
rect 5813 37247 5871 37253
rect 5813 37213 5825 37247
rect 5859 37244 5871 37247
rect 6733 37247 6791 37253
rect 5859 37216 6592 37244
rect 5859 37213 5871 37216
rect 5813 37207 5871 37213
rect 4614 37068 4620 37120
rect 4672 37108 4678 37120
rect 4709 37111 4767 37117
rect 4709 37108 4721 37111
rect 4672 37080 4721 37108
rect 4672 37068 4678 37080
rect 4709 37077 4721 37080
rect 4755 37077 4767 37111
rect 4709 37071 4767 37077
rect 5534 37068 5540 37120
rect 5592 37108 5598 37120
rect 6564 37117 6592 37216
rect 6733 37213 6745 37247
rect 6779 37244 6791 37247
rect 6914 37244 6920 37256
rect 6779 37216 6920 37244
rect 6779 37213 6791 37216
rect 6733 37207 6791 37213
rect 6914 37204 6920 37216
rect 6972 37204 6978 37256
rect 7653 37247 7711 37253
rect 7653 37213 7665 37247
rect 7699 37244 7711 37247
rect 8202 37244 8208 37256
rect 7699 37216 8208 37244
rect 7699 37213 7711 37216
rect 7653 37207 7711 37213
rect 8202 37204 8208 37216
rect 8260 37204 8266 37256
rect 8570 37244 8576 37256
rect 8531 37216 8576 37244
rect 8570 37204 8576 37216
rect 8628 37204 8634 37256
rect 9493 37247 9551 37253
rect 9493 37213 9505 37247
rect 9539 37244 9551 37247
rect 9766 37244 9772 37256
rect 9539 37216 9772 37244
rect 9539 37213 9551 37216
rect 9493 37207 9551 37213
rect 9766 37204 9772 37216
rect 9824 37204 9830 37256
rect 10042 37204 10048 37256
rect 10100 37244 10106 37256
rect 10137 37247 10195 37253
rect 10137 37244 10149 37247
rect 10100 37216 10149 37244
rect 10100 37204 10106 37216
rect 10137 37213 10149 37216
rect 10183 37213 10195 37247
rect 10137 37207 10195 37213
rect 11149 37247 11207 37253
rect 11149 37213 11161 37247
rect 11195 37213 11207 37247
rect 12250 37244 12256 37256
rect 12211 37216 12256 37244
rect 11149 37207 11207 37213
rect 11164 37176 11192 37207
rect 12250 37204 12256 37216
rect 12308 37204 12314 37256
rect 13170 37244 13176 37256
rect 13131 37216 13176 37244
rect 13170 37204 13176 37216
rect 13228 37204 13234 37256
rect 15013 37247 15071 37253
rect 15013 37213 15025 37247
rect 15059 37213 15071 37247
rect 15930 37244 15936 37256
rect 15891 37216 15936 37244
rect 15013 37207 15071 37213
rect 15028 37176 15056 37207
rect 15930 37204 15936 37216
rect 15988 37204 15994 37256
rect 17129 37247 17187 37253
rect 17129 37213 17141 37247
rect 17175 37244 17187 37247
rect 17310 37244 17316 37256
rect 17175 37216 17316 37244
rect 17175 37213 17187 37216
rect 17129 37207 17187 37213
rect 17310 37204 17316 37216
rect 17368 37204 17374 37256
rect 17402 37204 17408 37256
rect 17460 37244 17466 37256
rect 17589 37247 17647 37253
rect 17589 37244 17601 37247
rect 17460 37216 17601 37244
rect 17460 37204 17466 37216
rect 17589 37213 17601 37216
rect 17635 37213 17647 37247
rect 17589 37207 17647 37213
rect 18693 37247 18751 37253
rect 18693 37213 18705 37247
rect 18739 37244 18751 37247
rect 19058 37244 19064 37256
rect 18739 37216 19064 37244
rect 18739 37213 18751 37216
rect 18693 37207 18751 37213
rect 19058 37204 19064 37216
rect 19116 37204 19122 37256
rect 19702 37244 19708 37256
rect 19663 37216 19708 37244
rect 19702 37204 19708 37216
rect 19760 37204 19766 37256
rect 20533 37247 20591 37253
rect 20533 37213 20545 37247
rect 20579 37244 20591 37247
rect 20622 37244 20628 37256
rect 20579 37216 20628 37244
rect 20579 37213 20591 37216
rect 20533 37207 20591 37213
rect 20622 37204 20628 37216
rect 20680 37204 20686 37256
rect 20714 37204 20720 37256
rect 20772 37244 20778 37256
rect 21177 37247 21235 37253
rect 21177 37244 21189 37247
rect 20772 37216 21189 37244
rect 20772 37204 20778 37216
rect 21177 37213 21189 37216
rect 21223 37213 21235 37247
rect 22278 37244 22284 37256
rect 21177 37207 21235 37213
rect 21284 37216 22284 37244
rect 21284 37176 21312 37216
rect 22278 37204 22284 37216
rect 22336 37204 22342 37256
rect 22388 37253 22416 37352
rect 29086 37340 29092 37352
rect 29144 37340 29150 37392
rect 29181 37383 29239 37389
rect 29181 37349 29193 37383
rect 29227 37380 29239 37383
rect 29638 37380 29644 37392
rect 29227 37352 29644 37380
rect 29227 37349 29239 37352
rect 29181 37343 29239 37349
rect 29638 37340 29644 37352
rect 29696 37340 29702 37392
rect 30944 37380 30972 37420
rect 31018 37408 31024 37460
rect 31076 37448 31082 37460
rect 44453 37451 44511 37457
rect 44453 37448 44465 37451
rect 31076 37420 44465 37448
rect 31076 37408 31082 37420
rect 44453 37417 44465 37420
rect 44499 37417 44511 37451
rect 45370 37448 45376 37460
rect 45331 37420 45376 37448
rect 44453 37411 44511 37417
rect 45370 37408 45376 37420
rect 45428 37408 45434 37460
rect 47854 37408 47860 37460
rect 47912 37448 47918 37460
rect 50341 37451 50399 37457
rect 50341 37448 50353 37451
rect 47912 37420 50353 37448
rect 47912 37408 47918 37420
rect 50341 37417 50353 37420
rect 50387 37448 50399 37451
rect 51718 37448 51724 37460
rect 50387 37420 51724 37448
rect 50387 37417 50399 37420
rect 50341 37411 50399 37417
rect 51718 37408 51724 37420
rect 51776 37408 51782 37460
rect 54205 37451 54263 37457
rect 54205 37417 54217 37451
rect 54251 37448 54263 37451
rect 55214 37448 55220 37460
rect 54251 37420 55220 37448
rect 54251 37417 54263 37420
rect 54205 37411 54263 37417
rect 55214 37408 55220 37420
rect 55272 37408 55278 37460
rect 55585 37451 55643 37457
rect 55585 37417 55597 37451
rect 55631 37448 55643 37451
rect 57514 37448 57520 37460
rect 55631 37420 57520 37448
rect 55631 37417 55643 37420
rect 55585 37411 55643 37417
rect 57514 37408 57520 37420
rect 57572 37408 57578 37460
rect 58069 37451 58127 37457
rect 58069 37417 58081 37451
rect 58115 37448 58127 37451
rect 58158 37448 58164 37460
rect 58115 37420 58164 37448
rect 58115 37417 58127 37420
rect 58069 37411 58127 37417
rect 58158 37408 58164 37420
rect 58216 37408 58222 37460
rect 59357 37451 59415 37457
rect 59357 37417 59369 37451
rect 59403 37448 59415 37451
rect 62390 37448 62396 37460
rect 59403 37420 62396 37448
rect 59403 37417 59415 37420
rect 59357 37411 59415 37417
rect 62390 37408 62396 37420
rect 62448 37408 62454 37460
rect 72326 37408 72332 37460
rect 72384 37448 72390 37460
rect 72384 37420 79272 37448
rect 72384 37408 72390 37420
rect 58342 37380 58348 37392
rect 30944 37352 58348 37380
rect 58342 37340 58348 37352
rect 58400 37340 58406 37392
rect 59814 37380 59820 37392
rect 59775 37352 59820 37380
rect 59814 37340 59820 37352
rect 59872 37340 59878 37392
rect 60829 37383 60887 37389
rect 60829 37349 60841 37383
rect 60875 37380 60887 37383
rect 61102 37380 61108 37392
rect 60875 37352 61108 37380
rect 60875 37349 60887 37352
rect 60829 37343 60887 37349
rect 61102 37340 61108 37352
rect 61160 37340 61166 37392
rect 65058 37380 65064 37392
rect 64616 37352 65064 37380
rect 25041 37315 25099 37321
rect 25041 37312 25053 37315
rect 23952 37284 25053 37312
rect 22373 37247 22431 37253
rect 22373 37213 22385 37247
rect 22419 37244 22431 37247
rect 22462 37244 22468 37256
rect 22419 37216 22468 37244
rect 22419 37213 22431 37216
rect 22373 37207 22431 37213
rect 22462 37204 22468 37216
rect 22520 37204 22526 37256
rect 23290 37244 23296 37256
rect 23251 37216 23296 37244
rect 23290 37204 23296 37216
rect 23348 37204 23354 37256
rect 23382 37204 23388 37256
rect 23440 37244 23446 37256
rect 23952 37244 23980 37284
rect 25041 37281 25053 37284
rect 25087 37281 25099 37315
rect 25041 37275 25099 37281
rect 25130 37272 25136 37324
rect 25188 37312 25194 37324
rect 27982 37312 27988 37324
rect 25188 37284 26464 37312
rect 27943 37284 27988 37312
rect 25188 37272 25194 37284
rect 23440 37216 23980 37244
rect 24029 37247 24087 37253
rect 23440 37204 23446 37216
rect 24029 37213 24041 37247
rect 24075 37244 24087 37247
rect 24670 37244 24676 37256
rect 24075 37216 24676 37244
rect 24075 37213 24087 37216
rect 24029 37207 24087 37213
rect 24670 37204 24676 37216
rect 24728 37204 24734 37256
rect 25866 37244 25872 37256
rect 24780 37216 25872 37244
rect 11164 37148 14964 37176
rect 15028 37148 21312 37176
rect 5629 37111 5687 37117
rect 5629 37108 5641 37111
rect 5592 37080 5641 37108
rect 5592 37068 5598 37080
rect 5629 37077 5641 37080
rect 5675 37077 5687 37111
rect 5629 37071 5687 37077
rect 6549 37111 6607 37117
rect 6549 37077 6561 37111
rect 6595 37077 6607 37111
rect 6549 37071 6607 37077
rect 7282 37068 7288 37120
rect 7340 37108 7346 37120
rect 7469 37111 7527 37117
rect 7469 37108 7481 37111
rect 7340 37080 7481 37108
rect 7340 37068 7346 37080
rect 7469 37077 7481 37080
rect 7515 37077 7527 37111
rect 7469 37071 7527 37077
rect 8294 37068 8300 37120
rect 8352 37108 8358 37120
rect 8389 37111 8447 37117
rect 8389 37108 8401 37111
rect 8352 37080 8401 37108
rect 8352 37068 8358 37080
rect 8389 37077 8401 37080
rect 8435 37077 8447 37111
rect 8389 37071 8447 37077
rect 9122 37068 9128 37120
rect 9180 37108 9186 37120
rect 9309 37111 9367 37117
rect 9309 37108 9321 37111
rect 9180 37080 9321 37108
rect 9180 37068 9186 37080
rect 9309 37077 9321 37080
rect 9355 37077 9367 37111
rect 10318 37108 10324 37120
rect 10279 37080 10324 37108
rect 9309 37071 9367 37077
rect 10318 37068 10324 37080
rect 10376 37068 10382 37120
rect 10962 37108 10968 37120
rect 10923 37080 10968 37108
rect 10962 37068 10968 37080
rect 11020 37068 11026 37120
rect 11882 37068 11888 37120
rect 11940 37108 11946 37120
rect 12069 37111 12127 37117
rect 12069 37108 12081 37111
rect 11940 37080 12081 37108
rect 11940 37068 11946 37080
rect 12069 37077 12081 37080
rect 12115 37077 12127 37111
rect 12069 37071 12127 37077
rect 12802 37068 12808 37120
rect 12860 37108 12866 37120
rect 12989 37111 13047 37117
rect 12989 37108 13001 37111
rect 12860 37080 13001 37108
rect 12860 37068 12866 37080
rect 12989 37077 13001 37080
rect 13035 37077 13047 37111
rect 12989 37071 13047 37077
rect 14642 37068 14648 37120
rect 14700 37108 14706 37120
rect 14829 37111 14887 37117
rect 14829 37108 14841 37111
rect 14700 37080 14841 37108
rect 14700 37068 14706 37080
rect 14829 37077 14841 37080
rect 14875 37077 14887 37111
rect 14936 37108 14964 37148
rect 21542 37136 21548 37188
rect 21600 37176 21606 37188
rect 21600 37148 23888 37176
rect 21600 37136 21606 37148
rect 15470 37108 15476 37120
rect 14936 37080 15476 37108
rect 14829 37071 14887 37077
rect 15470 37068 15476 37080
rect 15528 37068 15534 37120
rect 15562 37068 15568 37120
rect 15620 37108 15626 37120
rect 15749 37111 15807 37117
rect 15749 37108 15761 37111
rect 15620 37080 15761 37108
rect 15620 37068 15626 37080
rect 15749 37077 15761 37080
rect 15795 37077 15807 37111
rect 15749 37071 15807 37077
rect 16574 37068 16580 37120
rect 16632 37108 16638 37120
rect 16945 37111 17003 37117
rect 16945 37108 16957 37111
rect 16632 37080 16957 37108
rect 16632 37068 16638 37080
rect 16945 37077 16957 37080
rect 16991 37077 17003 37111
rect 17770 37108 17776 37120
rect 17731 37080 17776 37108
rect 16945 37071 17003 37077
rect 17770 37068 17776 37080
rect 17828 37068 17834 37120
rect 18322 37068 18328 37120
rect 18380 37108 18386 37120
rect 18509 37111 18567 37117
rect 18509 37108 18521 37111
rect 18380 37080 18521 37108
rect 18380 37068 18386 37080
rect 18509 37077 18521 37080
rect 18555 37077 18567 37111
rect 18509 37071 18567 37077
rect 19334 37068 19340 37120
rect 19392 37108 19398 37120
rect 19521 37111 19579 37117
rect 19521 37108 19533 37111
rect 19392 37080 19533 37108
rect 19392 37068 19398 37080
rect 19521 37077 19533 37080
rect 19567 37077 19579 37111
rect 19521 37071 19579 37077
rect 20162 37068 20168 37120
rect 20220 37108 20226 37120
rect 20349 37111 20407 37117
rect 20349 37108 20361 37111
rect 20220 37080 20361 37108
rect 20220 37068 20226 37080
rect 20349 37077 20361 37080
rect 20395 37077 20407 37111
rect 21358 37108 21364 37120
rect 21319 37080 21364 37108
rect 20349 37071 20407 37077
rect 21358 37068 21364 37080
rect 21416 37068 21422 37120
rect 22094 37068 22100 37120
rect 22152 37108 22158 37120
rect 22189 37111 22247 37117
rect 22189 37108 22201 37111
rect 22152 37080 22201 37108
rect 22152 37068 22158 37080
rect 22189 37077 22201 37080
rect 22235 37077 22247 37111
rect 22189 37071 22247 37077
rect 22922 37068 22928 37120
rect 22980 37108 22986 37120
rect 23860 37117 23888 37148
rect 23934 37136 23940 37188
rect 23992 37176 23998 37188
rect 24780 37176 24808 37216
rect 25866 37204 25872 37216
rect 25924 37204 25930 37256
rect 26329 37247 26387 37253
rect 26329 37244 26341 37247
rect 26206 37216 26341 37244
rect 23992 37148 24808 37176
rect 23992 37136 23998 37148
rect 25038 37136 25044 37188
rect 25096 37176 25102 37188
rect 25225 37179 25283 37185
rect 25225 37176 25237 37179
rect 25096 37148 25237 37176
rect 25096 37136 25102 37148
rect 25225 37145 25237 37148
rect 25271 37176 25283 37179
rect 25498 37176 25504 37188
rect 25271 37148 25504 37176
rect 25271 37145 25283 37148
rect 25225 37139 25283 37145
rect 25498 37136 25504 37148
rect 25556 37176 25562 37188
rect 25958 37176 25964 37188
rect 25556 37148 25964 37176
rect 25556 37136 25562 37148
rect 25958 37136 25964 37148
rect 26016 37136 26022 37188
rect 23109 37111 23167 37117
rect 23109 37108 23121 37111
rect 22980 37080 23121 37108
rect 22980 37068 22986 37080
rect 23109 37077 23121 37080
rect 23155 37077 23167 37111
rect 23109 37071 23167 37077
rect 23845 37111 23903 37117
rect 23845 37077 23857 37111
rect 23891 37077 23903 37111
rect 23845 37071 23903 37077
rect 24026 37068 24032 37120
rect 24084 37108 24090 37120
rect 24655 37111 24713 37117
rect 24655 37108 24667 37111
rect 24084 37080 24667 37108
rect 24084 37068 24090 37080
rect 24655 37077 24667 37080
rect 24701 37077 24713 37111
rect 25130 37108 25136 37120
rect 25091 37080 25136 37108
rect 24655 37071 24713 37077
rect 25130 37068 25136 37080
rect 25188 37068 25194 37120
rect 25314 37068 25320 37120
rect 25372 37108 25378 37120
rect 25777 37111 25835 37117
rect 25777 37108 25789 37111
rect 25372 37080 25789 37108
rect 25372 37068 25378 37080
rect 25777 37077 25789 37080
rect 25823 37108 25835 37111
rect 26206 37108 26234 37216
rect 26329 37213 26341 37216
rect 26375 37213 26387 37247
rect 26436 37244 26464 37284
rect 27982 37272 27988 37284
rect 28040 37272 28046 37324
rect 28077 37315 28135 37321
rect 28077 37281 28089 37315
rect 28123 37281 28135 37315
rect 30006 37312 30012 37324
rect 29967 37284 30012 37312
rect 28077 37275 28135 37281
rect 27338 37244 27344 37256
rect 26436 37216 27200 37244
rect 27299 37216 27344 37244
rect 26329 37207 26387 37213
rect 26510 37108 26516 37120
rect 25823 37080 26234 37108
rect 26471 37080 26516 37108
rect 25823 37077 25835 37080
rect 25777 37071 25835 37077
rect 26510 37068 26516 37080
rect 26568 37068 26574 37120
rect 27172 37117 27200 37216
rect 27338 37204 27344 37216
rect 27396 37204 27402 37256
rect 28092 37244 28120 37275
rect 30006 37272 30012 37284
rect 30064 37272 30070 37324
rect 33594 37312 33600 37324
rect 33555 37284 33600 37312
rect 33594 37272 33600 37284
rect 33652 37272 33658 37324
rect 35621 37315 35679 37321
rect 35621 37281 35633 37315
rect 35667 37312 35679 37315
rect 36817 37315 36875 37321
rect 36817 37312 36829 37315
rect 35667 37284 36829 37312
rect 35667 37281 35679 37284
rect 35621 37275 35679 37281
rect 36817 37281 36829 37284
rect 36863 37312 36875 37315
rect 37550 37312 37556 37324
rect 36863 37284 37556 37312
rect 36863 37281 36875 37284
rect 36817 37275 36875 37281
rect 37550 37272 37556 37284
rect 37608 37312 37614 37324
rect 38565 37315 38623 37321
rect 38565 37312 38577 37315
rect 37608 37284 38577 37312
rect 37608 37272 37614 37284
rect 38565 37281 38577 37284
rect 38611 37312 38623 37315
rect 40862 37312 40868 37324
rect 38611 37284 40868 37312
rect 38611 37281 38623 37284
rect 38565 37275 38623 37281
rect 40862 37272 40868 37284
rect 40920 37312 40926 37324
rect 41325 37315 41383 37321
rect 41325 37312 41337 37315
rect 40920 37284 41337 37312
rect 40920 37272 40926 37284
rect 41325 37281 41337 37284
rect 41371 37281 41383 37315
rect 41325 37275 41383 37281
rect 42061 37315 42119 37321
rect 42061 37281 42073 37315
rect 42107 37312 42119 37315
rect 46198 37312 46204 37324
rect 42107 37284 44588 37312
rect 46159 37284 46204 37312
rect 42107 37281 42119 37284
rect 42061 37275 42119 37281
rect 28718 37244 28724 37256
rect 28092 37216 28724 37244
rect 28718 37204 28724 37216
rect 28776 37244 28782 37256
rect 28902 37244 28908 37256
rect 28776 37216 28908 37244
rect 28776 37204 28782 37216
rect 28902 37204 28908 37216
rect 28960 37204 28966 37256
rect 28997 37247 29055 37253
rect 28997 37213 29009 37247
rect 29043 37213 29055 37247
rect 28997 37207 29055 37213
rect 27246 37136 27252 37188
rect 27304 37176 27310 37188
rect 29012 37176 29040 37207
rect 31294 37204 31300 37256
rect 31352 37244 31358 37256
rect 31573 37247 31631 37253
rect 31573 37244 31585 37247
rect 31352 37216 31585 37244
rect 31352 37204 31358 37216
rect 31573 37213 31585 37216
rect 31619 37213 31631 37247
rect 31573 37207 31631 37213
rect 32309 37247 32367 37253
rect 32309 37213 32321 37247
rect 32355 37213 32367 37247
rect 34330 37244 34336 37256
rect 34291 37216 34336 37244
rect 32309 37207 32367 37213
rect 29362 37176 29368 37188
rect 27304 37148 28856 37176
rect 29012 37148 29368 37176
rect 27304 37136 27310 37148
rect 27157 37111 27215 37117
rect 27157 37077 27169 37111
rect 27203 37077 27215 37111
rect 28166 37108 28172 37120
rect 28127 37080 28172 37108
rect 27157 37071 27215 37077
rect 28166 37068 28172 37080
rect 28224 37068 28230 37120
rect 28537 37111 28595 37117
rect 28537 37077 28549 37111
rect 28583 37108 28595 37111
rect 28626 37108 28632 37120
rect 28583 37080 28632 37108
rect 28583 37077 28595 37080
rect 28537 37071 28595 37077
rect 28626 37068 28632 37080
rect 28684 37068 28690 37120
rect 28828 37108 28856 37148
rect 29362 37136 29368 37148
rect 29420 37136 29426 37188
rect 29822 37176 29828 37188
rect 29783 37148 29828 37176
rect 29822 37136 29828 37148
rect 29880 37136 29886 37188
rect 30653 37179 30711 37185
rect 30653 37145 30665 37179
rect 30699 37176 30711 37179
rect 30742 37176 30748 37188
rect 30699 37148 30748 37176
rect 30699 37145 30711 37148
rect 30653 37139 30711 37145
rect 30742 37136 30748 37148
rect 30800 37136 30806 37188
rect 30837 37179 30895 37185
rect 30837 37145 30849 37179
rect 30883 37176 30895 37179
rect 31754 37176 31760 37188
rect 30883 37148 31760 37176
rect 30883 37145 30895 37148
rect 30837 37139 30895 37145
rect 31754 37136 31760 37148
rect 31812 37136 31818 37188
rect 31110 37108 31116 37120
rect 28828 37080 31116 37108
rect 31110 37068 31116 37080
rect 31168 37068 31174 37120
rect 31202 37068 31208 37120
rect 31260 37108 31266 37120
rect 31389 37111 31447 37117
rect 31389 37108 31401 37111
rect 31260 37080 31401 37108
rect 31260 37068 31266 37080
rect 31389 37077 31401 37080
rect 31435 37077 31447 37111
rect 31389 37071 31447 37077
rect 31478 37068 31484 37120
rect 31536 37108 31542 37120
rect 32324 37108 32352 37207
rect 34330 37204 34336 37216
rect 34388 37204 34394 37256
rect 34698 37204 34704 37256
rect 34756 37244 34762 37256
rect 38289 37247 38347 37253
rect 38289 37244 38301 37247
rect 34756 37216 38301 37244
rect 34756 37204 34762 37216
rect 38289 37213 38301 37216
rect 38335 37213 38347 37247
rect 39390 37244 39396 37256
rect 39351 37216 39396 37244
rect 38289 37207 38347 37213
rect 39390 37204 39396 37216
rect 39448 37204 39454 37256
rect 40034 37244 40040 37256
rect 39995 37216 40040 37244
rect 40034 37204 40040 37216
rect 40092 37204 40098 37256
rect 40126 37204 40132 37256
rect 40184 37244 40190 37256
rect 42702 37244 42708 37256
rect 40184 37216 42708 37244
rect 40184 37204 40190 37216
rect 42702 37204 42708 37216
rect 42760 37204 42766 37256
rect 42794 37204 42800 37256
rect 42852 37244 42858 37256
rect 44560 37253 44588 37284
rect 46198 37272 46204 37284
rect 46256 37272 46262 37324
rect 46860 37284 47164 37312
rect 42981 37247 43039 37253
rect 42981 37244 42993 37247
rect 42852 37216 42993 37244
rect 42852 37204 42858 37216
rect 42981 37213 42993 37216
rect 43027 37213 43039 37247
rect 42981 37207 43039 37213
rect 44545 37247 44603 37253
rect 44545 37213 44557 37247
rect 44591 37244 44603 37247
rect 45281 37247 45339 37253
rect 45281 37244 45293 37247
rect 44591 37216 45293 37244
rect 44591 37213 44603 37216
rect 44545 37207 44603 37213
rect 45281 37213 45293 37216
rect 45327 37213 45339 37247
rect 45281 37207 45339 37213
rect 32950 37136 32956 37188
rect 33008 37176 33014 37188
rect 33413 37179 33471 37185
rect 33413 37176 33425 37179
rect 33008 37148 33425 37176
rect 33008 37136 33014 37148
rect 33413 37145 33425 37148
rect 33459 37145 33471 37179
rect 33413 37139 33471 37145
rect 33594 37136 33600 37188
rect 33652 37176 33658 37188
rect 35345 37179 35403 37185
rect 35345 37176 35357 37179
rect 33652 37148 35357 37176
rect 33652 37136 33658 37148
rect 35345 37145 35357 37148
rect 35391 37145 35403 37179
rect 35526 37176 35532 37188
rect 35487 37148 35532 37176
rect 35345 37139 35403 37145
rect 35526 37136 35532 37148
rect 35584 37136 35590 37188
rect 35710 37136 35716 37188
rect 35768 37176 35774 37188
rect 41141 37179 41199 37185
rect 41141 37176 41153 37179
rect 35768 37148 41153 37176
rect 35768 37136 35774 37148
rect 41141 37145 41153 37148
rect 41187 37145 41199 37179
rect 43257 37179 43315 37185
rect 43257 37176 43269 37179
rect 41141 37139 41199 37145
rect 42996 37148 43269 37176
rect 32490 37108 32496 37120
rect 31536 37080 32352 37108
rect 32451 37080 32496 37108
rect 31536 37068 31542 37080
rect 32490 37068 32496 37080
rect 32548 37068 32554 37120
rect 34149 37111 34207 37117
rect 34149 37077 34161 37111
rect 34195 37108 34207 37111
rect 34422 37108 34428 37120
rect 34195 37080 34428 37108
rect 34195 37077 34207 37080
rect 34149 37071 34207 37077
rect 34422 37068 34428 37080
rect 34480 37068 34486 37120
rect 34790 37068 34796 37120
rect 34848 37108 34854 37120
rect 35051 37111 35109 37117
rect 35051 37108 35063 37111
rect 34848 37080 35063 37108
rect 34848 37068 34854 37080
rect 35051 37077 35063 37080
rect 35097 37077 35109 37111
rect 35051 37071 35109 37077
rect 36078 37068 36084 37120
rect 36136 37108 36142 37120
rect 36173 37111 36231 37117
rect 36173 37108 36185 37111
rect 36136 37080 36185 37108
rect 36136 37068 36142 37080
rect 36173 37077 36185 37080
rect 36219 37077 36231 37111
rect 36538 37108 36544 37120
rect 36499 37080 36544 37108
rect 36173 37071 36231 37077
rect 36538 37068 36544 37080
rect 36596 37068 36602 37120
rect 36630 37068 36636 37120
rect 36688 37108 36694 37120
rect 37921 37111 37979 37117
rect 36688 37080 36733 37108
rect 36688 37068 36694 37080
rect 37921 37077 37933 37111
rect 37967 37108 37979 37111
rect 38194 37108 38200 37120
rect 37967 37080 38200 37108
rect 37967 37077 37979 37080
rect 37921 37071 37979 37077
rect 38194 37068 38200 37080
rect 38252 37068 38258 37120
rect 38381 37111 38439 37117
rect 38381 37077 38393 37111
rect 38427 37108 38439 37111
rect 38470 37108 38476 37120
rect 38427 37080 38476 37108
rect 38427 37077 38439 37080
rect 38381 37071 38439 37077
rect 38470 37068 38476 37080
rect 38528 37068 38534 37120
rect 38654 37068 38660 37120
rect 38712 37108 38718 37120
rect 39209 37111 39267 37117
rect 39209 37108 39221 37111
rect 38712 37080 39221 37108
rect 38712 37068 38718 37080
rect 39209 37077 39221 37080
rect 39255 37077 39267 37111
rect 39209 37071 39267 37077
rect 40221 37111 40279 37117
rect 40221 37077 40233 37111
rect 40267 37108 40279 37111
rect 40402 37108 40408 37120
rect 40267 37080 40408 37108
rect 40267 37077 40279 37080
rect 40221 37071 40279 37077
rect 40402 37068 40408 37080
rect 40460 37068 40466 37120
rect 40586 37068 40592 37120
rect 40644 37108 40650 37120
rect 40773 37111 40831 37117
rect 40773 37108 40785 37111
rect 40644 37080 40785 37108
rect 40644 37068 40650 37080
rect 40773 37077 40785 37080
rect 40819 37077 40831 37111
rect 40773 37071 40831 37077
rect 41230 37068 41236 37120
rect 41288 37108 41294 37120
rect 41288 37080 41333 37108
rect 41288 37068 41294 37080
rect 41506 37068 41512 37120
rect 41564 37108 41570 37120
rect 42996 37108 43024 37148
rect 43257 37145 43269 37148
rect 43303 37145 43315 37179
rect 43806 37176 43812 37188
rect 43257 37139 43315 37145
rect 43364 37148 43812 37176
rect 41564 37080 43024 37108
rect 43073 37111 43131 37117
rect 41564 37068 41570 37080
rect 43073 37077 43085 37111
rect 43119 37108 43131 37111
rect 43364 37108 43392 37148
rect 43806 37136 43812 37148
rect 43864 37136 43870 37188
rect 45296 37176 45324 37207
rect 45370 37204 45376 37256
rect 45428 37244 45434 37256
rect 46017 37247 46075 37253
rect 46017 37244 46029 37247
rect 45428 37216 46029 37244
rect 45428 37204 45434 37216
rect 46017 37213 46029 37216
rect 46063 37213 46075 37247
rect 46860 37244 46888 37284
rect 46017 37207 46075 37213
rect 46124 37216 46888 37244
rect 45646 37176 45652 37188
rect 45296 37148 45652 37176
rect 45646 37136 45652 37148
rect 45704 37136 45710 37188
rect 45830 37136 45836 37188
rect 45888 37176 45894 37188
rect 46124 37176 46152 37216
rect 46934 37204 46940 37256
rect 46992 37244 46998 37256
rect 47136 37244 47164 37284
rect 47854 37272 47860 37324
rect 47912 37312 47918 37324
rect 47949 37315 48007 37321
rect 47949 37312 47961 37315
rect 47912 37284 47961 37312
rect 47912 37272 47918 37284
rect 47949 37281 47961 37284
rect 47995 37281 48007 37315
rect 48130 37312 48136 37324
rect 48091 37284 48136 37312
rect 47949 37275 48007 37281
rect 48130 37272 48136 37284
rect 48188 37272 48194 37324
rect 51718 37312 51724 37324
rect 49712 37284 50016 37312
rect 46992 37216 47037 37244
rect 47136 37216 48360 37244
rect 46992 37204 46998 37216
rect 48225 37179 48283 37185
rect 48225 37176 48237 37179
rect 45888 37148 46152 37176
rect 46216 37148 48237 37176
rect 45888 37136 45894 37148
rect 43119 37080 43392 37108
rect 43119 37077 43131 37080
rect 43073 37071 43131 37077
rect 43438 37068 43444 37120
rect 43496 37108 43502 37120
rect 43543 37111 43601 37117
rect 43543 37108 43555 37111
rect 43496 37080 43555 37108
rect 43496 37068 43502 37080
rect 43543 37077 43555 37080
rect 43589 37077 43601 37111
rect 43543 37071 43601 37077
rect 43714 37068 43720 37120
rect 43772 37108 43778 37120
rect 46216 37108 46244 37148
rect 48225 37145 48237 37148
rect 48271 37145 48283 37179
rect 48332 37176 48360 37216
rect 48498 37204 48504 37256
rect 48556 37244 48562 37256
rect 49712 37244 49740 37284
rect 48556 37216 49740 37244
rect 48556 37204 48562 37216
rect 49786 37204 49792 37256
rect 49844 37244 49850 37256
rect 49988 37244 50016 37284
rect 51092 37284 51396 37312
rect 51679 37284 51724 37312
rect 51092 37244 51120 37284
rect 49844 37216 49889 37244
rect 49988 37216 51120 37244
rect 49844 37204 49850 37216
rect 51166 37204 51172 37256
rect 51224 37244 51230 37256
rect 51368 37244 51396 37284
rect 51718 37272 51724 37284
rect 51776 37312 51782 37324
rect 53009 37315 53067 37321
rect 53009 37312 53021 37315
rect 51776 37284 53021 37312
rect 51776 37272 51782 37284
rect 53009 37281 53021 37284
rect 53055 37281 53067 37315
rect 53009 37275 53067 37281
rect 57425 37315 57483 37321
rect 57425 37281 57437 37315
rect 57471 37312 57483 37315
rect 58250 37312 58256 37324
rect 57471 37284 58256 37312
rect 57471 37281 57483 37284
rect 57425 37275 57483 37281
rect 58250 37272 58256 37284
rect 58308 37272 58314 37324
rect 58618 37312 58624 37324
rect 58579 37284 58624 37312
rect 58618 37272 58624 37284
rect 58676 37272 58682 37324
rect 61286 37312 61292 37324
rect 61247 37284 61292 37312
rect 61286 37272 61292 37284
rect 61344 37272 61350 37324
rect 61378 37272 61384 37324
rect 61436 37312 61442 37324
rect 64616 37321 64644 37352
rect 65058 37340 65064 37352
rect 65116 37380 65122 37392
rect 66254 37380 66260 37392
rect 65116 37352 66260 37380
rect 65116 37340 65122 37352
rect 66254 37340 66260 37352
rect 66312 37380 66318 37392
rect 67542 37380 67548 37392
rect 66312 37352 66484 37380
rect 67503 37352 67548 37380
rect 66312 37340 66318 37352
rect 61473 37315 61531 37321
rect 61473 37312 61485 37315
rect 61436 37284 61485 37312
rect 61436 37272 61442 37284
rect 61473 37281 61485 37284
rect 61519 37312 61531 37315
rect 63405 37315 63463 37321
rect 63405 37312 63417 37315
rect 61519 37284 63417 37312
rect 61519 37281 61531 37284
rect 61473 37275 61531 37281
rect 63405 37281 63417 37284
rect 63451 37312 63463 37315
rect 64601 37315 64659 37321
rect 64601 37312 64613 37315
rect 63451 37284 64613 37312
rect 63451 37281 63463 37284
rect 63405 37275 63463 37281
rect 64601 37281 64613 37284
rect 64647 37281 64659 37315
rect 64601 37275 64659 37281
rect 64693 37315 64751 37321
rect 64693 37281 64705 37315
rect 64739 37312 64751 37315
rect 65150 37312 65156 37324
rect 64739 37284 65156 37312
rect 64739 37281 64751 37284
rect 64693 37275 64751 37281
rect 65150 37272 65156 37284
rect 65208 37272 65214 37324
rect 65426 37272 65432 37324
rect 65484 37312 65490 37324
rect 66349 37315 66407 37321
rect 66349 37312 66361 37315
rect 65484 37284 66361 37312
rect 65484 37272 65490 37284
rect 66349 37281 66361 37284
rect 66395 37281 66407 37315
rect 66456 37312 66484 37352
rect 67542 37340 67548 37352
rect 67600 37340 67606 37392
rect 67818 37340 67824 37392
rect 67876 37380 67882 37392
rect 79134 37380 79140 37392
rect 67876 37352 79140 37380
rect 67876 37340 67882 37352
rect 79134 37340 79140 37352
rect 79192 37340 79198 37392
rect 79244 37380 79272 37420
rect 79318 37408 79324 37460
rect 79376 37448 79382 37460
rect 80333 37451 80391 37457
rect 80333 37448 80345 37451
rect 79376 37420 80345 37448
rect 79376 37408 79382 37420
rect 80333 37417 80345 37420
rect 80379 37417 80391 37451
rect 80333 37411 80391 37417
rect 81342 37408 81348 37460
rect 81400 37448 81406 37460
rect 84013 37451 84071 37457
rect 81400 37420 83044 37448
rect 81400 37408 81406 37420
rect 81618 37380 81624 37392
rect 79244 37352 81624 37380
rect 81618 37340 81624 37352
rect 81676 37340 81682 37392
rect 68465 37315 68523 37321
rect 68465 37312 68477 37315
rect 66456 37284 68477 37312
rect 66349 37275 66407 37281
rect 68465 37281 68477 37284
rect 68511 37281 68523 37315
rect 68465 37275 68523 37281
rect 70854 37272 70860 37324
rect 70912 37312 70918 37324
rect 71041 37315 71099 37321
rect 71041 37312 71053 37315
rect 70912 37284 71053 37312
rect 70912 37272 70918 37284
rect 71041 37281 71053 37284
rect 71087 37312 71099 37315
rect 72973 37315 73031 37321
rect 71087 37284 72924 37312
rect 71087 37281 71099 37284
rect 71041 37275 71099 37281
rect 51997 37247 52055 37253
rect 51997 37244 52009 37247
rect 51224 37216 51269 37244
rect 51368 37216 52009 37244
rect 51224 37204 51230 37216
rect 51997 37213 52009 37216
rect 52043 37213 52055 37247
rect 51997 37207 52055 37213
rect 54938 37204 54944 37256
rect 54996 37244 55002 37256
rect 56045 37247 56103 37253
rect 54996 37216 55041 37244
rect 54996 37204 55002 37216
rect 56045 37213 56057 37247
rect 56091 37244 56103 37247
rect 56134 37244 56140 37256
rect 56091 37216 56140 37244
rect 56091 37213 56103 37216
rect 56045 37207 56103 37213
rect 56134 37204 56140 37216
rect 56192 37204 56198 37256
rect 56686 37204 56692 37256
rect 56744 37244 56750 37256
rect 58342 37244 58348 37256
rect 56744 37216 58348 37244
rect 56744 37204 56750 37216
rect 58342 37204 58348 37216
rect 58400 37204 58406 37256
rect 60706 37216 60964 37244
rect 53285 37179 53343 37185
rect 53285 37176 53297 37179
rect 48332 37148 53297 37176
rect 48225 37139 48283 37145
rect 53285 37145 53297 37148
rect 53331 37145 53343 37179
rect 53285 37139 53343 37145
rect 53558 37136 53564 37188
rect 53616 37176 53622 37188
rect 55582 37176 55588 37188
rect 53616 37148 55588 37176
rect 53616 37136 53622 37148
rect 55582 37136 55588 37148
rect 55640 37136 55646 37188
rect 55674 37136 55680 37188
rect 55732 37176 55738 37188
rect 59814 37176 59820 37188
rect 55732 37148 59820 37176
rect 55732 37136 55738 37148
rect 59814 37136 59820 37148
rect 59872 37136 59878 37188
rect 60001 37179 60059 37185
rect 60001 37145 60013 37179
rect 60047 37176 60059 37179
rect 60706 37176 60734 37216
rect 60047 37148 60734 37176
rect 60047 37145 60059 37148
rect 60001 37139 60059 37145
rect 43772 37080 46244 37108
rect 47121 37111 47179 37117
rect 43772 37068 43778 37080
rect 47121 37077 47133 37111
rect 47167 37108 47179 37111
rect 47762 37108 47768 37120
rect 47167 37080 47768 37108
rect 47167 37077 47179 37080
rect 47121 37071 47179 37077
rect 47762 37068 47768 37080
rect 47820 37068 47826 37120
rect 48593 37111 48651 37117
rect 48593 37077 48605 37111
rect 48639 37108 48651 37111
rect 48958 37108 48964 37120
rect 48639 37080 48964 37108
rect 48639 37077 48651 37080
rect 48593 37071 48651 37077
rect 48958 37068 48964 37080
rect 49016 37068 49022 37120
rect 49602 37108 49608 37120
rect 49563 37080 49608 37108
rect 49602 37068 49608 37080
rect 49660 37068 49666 37120
rect 50985 37111 51043 37117
rect 50985 37077 50997 37111
rect 51031 37108 51043 37111
rect 51442 37108 51448 37120
rect 51031 37080 51448 37108
rect 51031 37077 51043 37080
rect 50985 37071 51043 37077
rect 51442 37068 51448 37080
rect 51500 37068 51506 37120
rect 51534 37068 51540 37120
rect 51592 37108 51598 37120
rect 51905 37111 51963 37117
rect 51905 37108 51917 37111
rect 51592 37080 51917 37108
rect 51592 37068 51598 37080
rect 51905 37077 51917 37080
rect 51951 37077 51963 37111
rect 52362 37108 52368 37120
rect 52323 37080 52368 37108
rect 51905 37071 51963 37077
rect 52362 37068 52368 37080
rect 52420 37068 52426 37120
rect 53190 37108 53196 37120
rect 53151 37080 53196 37108
rect 53190 37068 53196 37080
rect 53248 37068 53254 37120
rect 53650 37108 53656 37120
rect 53611 37080 53656 37108
rect 53650 37068 53656 37080
rect 53708 37068 53714 37120
rect 54757 37111 54815 37117
rect 54757 37077 54769 37111
rect 54803 37108 54815 37111
rect 55122 37108 55128 37120
rect 54803 37080 55128 37108
rect 54803 37077 54815 37080
rect 54757 37071 54815 37077
rect 55122 37068 55128 37080
rect 55180 37068 55186 37120
rect 56229 37111 56287 37117
rect 56229 37077 56241 37111
rect 56275 37108 56287 37111
rect 56502 37108 56508 37120
rect 56275 37080 56508 37108
rect 56275 37077 56287 37080
rect 56229 37071 56287 37077
rect 56502 37068 56508 37080
rect 56560 37068 56566 37120
rect 56778 37108 56784 37120
rect 56739 37080 56784 37108
rect 56778 37068 56784 37080
rect 56836 37068 56842 37120
rect 57146 37108 57152 37120
rect 57107 37080 57152 37108
rect 57146 37068 57152 37080
rect 57204 37068 57210 37120
rect 57241 37111 57299 37117
rect 57241 37077 57253 37111
rect 57287 37108 57299 37111
rect 57514 37108 57520 37120
rect 57287 37080 57520 37108
rect 57287 37077 57299 37080
rect 57241 37071 57299 37077
rect 57514 37068 57520 37080
rect 57572 37068 57578 37120
rect 57974 37068 57980 37120
rect 58032 37108 58038 37120
rect 58437 37111 58495 37117
rect 58437 37108 58449 37111
rect 58032 37080 58449 37108
rect 58032 37068 58038 37080
rect 58437 37077 58449 37080
rect 58483 37077 58495 37111
rect 58437 37071 58495 37077
rect 58529 37111 58587 37117
rect 58529 37077 58541 37111
rect 58575 37108 58587 37111
rect 58618 37108 58624 37120
rect 58575 37080 58624 37108
rect 58575 37077 58587 37080
rect 58529 37071 58587 37077
rect 58618 37068 58624 37080
rect 58676 37068 58682 37120
rect 58710 37068 58716 37120
rect 58768 37108 58774 37120
rect 60734 37108 60740 37120
rect 58768 37080 60740 37108
rect 58768 37068 58774 37080
rect 60734 37068 60740 37080
rect 60792 37068 60798 37120
rect 60936 37108 60964 37216
rect 61010 37204 61016 37256
rect 61068 37244 61074 37256
rect 61197 37247 61255 37253
rect 61197 37244 61209 37247
rect 61068 37216 61209 37244
rect 61068 37204 61074 37216
rect 61197 37213 61209 37216
rect 61243 37213 61255 37247
rect 61197 37207 61255 37213
rect 61746 37204 61752 37256
rect 61804 37244 61810 37256
rect 62209 37247 62267 37253
rect 62209 37244 62221 37247
rect 61804 37216 62221 37244
rect 61804 37204 61810 37216
rect 62209 37213 62221 37216
rect 62255 37213 62267 37247
rect 63494 37244 63500 37256
rect 63455 37216 63500 37244
rect 62209 37207 62267 37213
rect 63494 37204 63500 37216
rect 63552 37244 63558 37256
rect 64138 37244 64144 37256
rect 63552 37216 64144 37244
rect 63552 37204 63558 37216
rect 64138 37204 64144 37216
rect 64196 37204 64202 37256
rect 64782 37244 64788 37256
rect 64743 37216 64788 37244
rect 64782 37204 64788 37216
rect 64840 37204 64846 37256
rect 64874 37204 64880 37256
rect 64932 37244 64938 37256
rect 65518 37244 65524 37256
rect 64932 37216 65524 37244
rect 64932 37204 64938 37216
rect 65518 37204 65524 37216
rect 65576 37204 65582 37256
rect 67266 37244 67272 37256
rect 66364 37216 67272 37244
rect 62390 37136 62396 37188
rect 62448 37176 62454 37188
rect 62448 37148 62493 37176
rect 62448 37136 62454 37148
rect 62574 37136 62580 37188
rect 62632 37176 62638 37188
rect 66254 37176 66260 37188
rect 62632 37148 66116 37176
rect 66215 37148 66260 37176
rect 62632 37136 62638 37148
rect 62025 37111 62083 37117
rect 62025 37108 62037 37111
rect 60936 37080 62037 37108
rect 62025 37077 62037 37080
rect 62071 37077 62083 37111
rect 62025 37071 62083 37077
rect 63586 37068 63592 37120
rect 63644 37108 63650 37120
rect 63957 37111 64015 37117
rect 63644 37080 63689 37108
rect 63644 37068 63650 37080
rect 63957 37077 63969 37111
rect 64003 37108 64015 37111
rect 64046 37108 64052 37120
rect 64003 37080 64052 37108
rect 64003 37077 64015 37080
rect 63957 37071 64015 37077
rect 64046 37068 64052 37080
rect 64104 37068 64110 37120
rect 65153 37111 65211 37117
rect 65153 37077 65165 37111
rect 65199 37108 65211 37111
rect 65978 37108 65984 37120
rect 65199 37080 65984 37108
rect 65199 37077 65211 37080
rect 65153 37071 65211 37077
rect 65978 37068 65984 37080
rect 66036 37068 66042 37120
rect 66088 37108 66116 37148
rect 66254 37136 66260 37148
rect 66312 37136 66318 37188
rect 66364 37185 66392 37216
rect 67266 37204 67272 37216
rect 67324 37244 67330 37256
rect 70213 37247 70271 37253
rect 67324 37216 68876 37244
rect 67324 37204 67330 37216
rect 66349 37179 66407 37185
rect 66349 37145 66361 37179
rect 66395 37145 66407 37179
rect 67726 37176 67732 37188
rect 66349 37139 66407 37145
rect 66456 37148 66944 37176
rect 67687 37148 67732 37176
rect 66456 37108 66484 37148
rect 66806 37108 66812 37120
rect 66864 37117 66870 37120
rect 66864 37111 66877 37117
rect 66088 37080 66484 37108
rect 66777 37080 66812 37108
rect 66806 37068 66812 37080
rect 66865 37077 66877 37111
rect 66916 37108 66944 37148
rect 67726 37136 67732 37148
rect 67784 37136 67790 37188
rect 68554 37136 68560 37188
rect 68612 37176 68618 37188
rect 68741 37179 68799 37185
rect 68612 37148 68657 37176
rect 68612 37136 68618 37148
rect 68741 37145 68753 37179
rect 68787 37145 68799 37179
rect 68848 37176 68876 37216
rect 70213 37213 70225 37247
rect 70259 37244 70271 37247
rect 70486 37244 70492 37256
rect 70259 37216 70492 37244
rect 70259 37213 70271 37216
rect 70213 37207 70271 37213
rect 70486 37204 70492 37216
rect 70544 37204 70550 37256
rect 72421 37247 72479 37253
rect 72421 37213 72433 37247
rect 72467 37244 72479 37247
rect 72510 37244 72516 37256
rect 72467 37216 72516 37244
rect 72467 37213 72479 37216
rect 72421 37207 72479 37213
rect 72510 37204 72516 37216
rect 72568 37204 72574 37256
rect 72896 37244 72924 37284
rect 72973 37281 72985 37315
rect 73019 37312 73031 37315
rect 75549 37315 75607 37321
rect 73019 37284 74672 37312
rect 73019 37281 73031 37284
rect 72973 37275 73031 37281
rect 74534 37244 74540 37256
rect 72896 37216 74540 37244
rect 74534 37204 74540 37216
rect 74592 37204 74598 37256
rect 74644 37253 74672 37284
rect 75549 37281 75561 37315
rect 75595 37312 75607 37315
rect 75822 37312 75828 37324
rect 75595 37284 75828 37312
rect 75595 37281 75607 37284
rect 75549 37275 75607 37281
rect 75822 37272 75828 37284
rect 75880 37272 75886 37324
rect 76190 37272 76196 37324
rect 76248 37312 76254 37324
rect 77018 37312 77024 37324
rect 76248 37284 77024 37312
rect 76248 37272 76254 37284
rect 77018 37272 77024 37284
rect 77076 37312 77082 37324
rect 79502 37312 79508 37324
rect 77076 37284 77708 37312
rect 79463 37284 79508 37312
rect 77076 37272 77082 37284
rect 74629 37247 74687 37253
rect 74629 37213 74641 37247
rect 74675 37213 74687 37247
rect 74629 37207 74687 37213
rect 71130 37176 71136 37188
rect 68848 37148 71136 37176
rect 68741 37139 68799 37145
rect 68756 37108 68784 37139
rect 71130 37136 71136 37148
rect 71188 37136 71194 37188
rect 71225 37179 71283 37185
rect 71225 37145 71237 37179
rect 71271 37176 71283 37179
rect 71590 37176 71596 37188
rect 71271 37148 71596 37176
rect 71271 37145 71283 37148
rect 71225 37139 71283 37145
rect 71590 37136 71596 37148
rect 71648 37136 71654 37188
rect 73614 37176 73620 37188
rect 73575 37148 73620 37176
rect 73614 37136 73620 37148
rect 73672 37136 73678 37188
rect 73798 37176 73804 37188
rect 73759 37148 73804 37176
rect 73798 37136 73804 37148
rect 73856 37136 73862 37188
rect 69014 37108 69020 37120
rect 69072 37117 69078 37120
rect 69072 37111 69085 37117
rect 66916 37080 68784 37108
rect 68985 37080 69020 37108
rect 66864 37071 66877 37077
rect 66864 37068 66870 37071
rect 69014 37068 69020 37080
rect 69073 37077 69085 37111
rect 69072 37071 69085 37077
rect 69072 37068 69078 37071
rect 69842 37068 69848 37120
rect 69900 37108 69906 37120
rect 70029 37111 70087 37117
rect 70029 37108 70041 37111
rect 69900 37080 70041 37108
rect 69900 37068 69906 37080
rect 70029 37077 70041 37080
rect 70075 37077 70087 37111
rect 70029 37071 70087 37077
rect 71314 37068 71320 37120
rect 71372 37108 71378 37120
rect 71372 37080 71417 37108
rect 71372 37068 71378 37080
rect 71498 37068 71504 37120
rect 71556 37108 71562 37120
rect 71685 37111 71743 37117
rect 71685 37108 71697 37111
rect 71556 37080 71697 37108
rect 71556 37068 71562 37080
rect 71685 37077 71697 37080
rect 71731 37077 71743 37111
rect 71685 37071 71743 37077
rect 71774 37068 71780 37120
rect 71832 37108 71838 37120
rect 72237 37111 72295 37117
rect 72237 37108 72249 37111
rect 71832 37080 72249 37108
rect 71832 37068 71838 37080
rect 72237 37077 72249 37080
rect 72283 37077 72295 37111
rect 72237 37071 72295 37077
rect 73522 37068 73528 37120
rect 73580 37108 73586 37120
rect 74445 37111 74503 37117
rect 74445 37108 74457 37111
rect 73580 37080 74457 37108
rect 73580 37068 73586 37080
rect 74445 37077 74457 37080
rect 74491 37077 74503 37111
rect 74644 37108 74672 37207
rect 74718 37204 74724 37256
rect 74776 37244 74782 37256
rect 74776 37216 77156 37244
rect 74776 37204 74782 37216
rect 75086 37136 75092 37188
rect 75144 37176 75150 37188
rect 75365 37179 75423 37185
rect 75365 37176 75377 37179
rect 75144 37148 75377 37176
rect 75144 37136 75150 37148
rect 75365 37145 75377 37148
rect 75411 37145 75423 37179
rect 75365 37139 75423 37145
rect 75546 37136 75552 37188
rect 75604 37176 75610 37188
rect 76745 37179 76803 37185
rect 76745 37176 76757 37179
rect 75604 37148 76757 37176
rect 75604 37136 75610 37148
rect 76745 37145 76757 37148
rect 76791 37145 76803 37179
rect 77128 37176 77156 37216
rect 77386 37204 77392 37256
rect 77444 37244 77450 37256
rect 77573 37247 77631 37253
rect 77573 37244 77585 37247
rect 77444 37216 77585 37244
rect 77444 37204 77450 37216
rect 77573 37213 77585 37216
rect 77619 37213 77631 37247
rect 77680 37244 77708 37284
rect 79502 37272 79508 37284
rect 79560 37272 79566 37324
rect 79689 37315 79747 37321
rect 79689 37281 79701 37315
rect 79735 37312 79747 37315
rect 79735 37284 79824 37312
rect 79735 37281 79747 37284
rect 79689 37275 79747 37281
rect 79796 37244 79824 37284
rect 80790 37272 80796 37324
rect 80848 37312 80854 37324
rect 81342 37312 81348 37324
rect 80848 37284 81348 37312
rect 80848 37272 80854 37284
rect 81342 37272 81348 37284
rect 81400 37312 81406 37324
rect 81437 37315 81495 37321
rect 81437 37312 81449 37315
rect 81400 37284 81449 37312
rect 81400 37272 81406 37284
rect 81437 37281 81449 37284
rect 81483 37281 81495 37315
rect 81437 37275 81495 37281
rect 81529 37315 81587 37321
rect 81529 37281 81541 37315
rect 81575 37312 81587 37315
rect 81575 37284 81848 37312
rect 81575 37281 81587 37284
rect 81529 37275 81587 37281
rect 77680 37216 79824 37244
rect 77573 37207 77631 37213
rect 79413 37179 79471 37185
rect 79413 37176 79425 37179
rect 77128 37148 79425 37176
rect 76745 37139 76803 37145
rect 79413 37145 79425 37148
rect 79459 37145 79471 37179
rect 79413 37139 79471 37145
rect 75730 37108 75736 37120
rect 74644 37080 75736 37108
rect 74445 37071 74503 37077
rect 75730 37068 75736 37080
rect 75788 37068 75794 37120
rect 76466 37117 76472 37120
rect 76459 37111 76472 37117
rect 76459 37077 76471 37111
rect 76524 37108 76530 37120
rect 76929 37111 76987 37117
rect 76524 37080 76559 37108
rect 76459 37071 76472 37077
rect 76466 37068 76472 37071
rect 76524 37068 76530 37080
rect 76929 37077 76941 37111
rect 76975 37108 76987 37111
rect 77110 37108 77116 37120
rect 76975 37080 77116 37108
rect 76975 37077 76987 37080
rect 76929 37071 76987 37077
rect 77110 37068 77116 37080
rect 77168 37068 77174 37120
rect 77294 37068 77300 37120
rect 77352 37108 77358 37120
rect 77757 37111 77815 37117
rect 77757 37108 77769 37111
rect 77352 37080 77769 37108
rect 77352 37068 77358 37080
rect 77757 37077 77769 37080
rect 77803 37077 77815 37111
rect 79042 37108 79048 37120
rect 79003 37080 79048 37108
rect 77757 37071 77815 37077
rect 79042 37068 79048 37080
rect 79100 37068 79106 37120
rect 79796 37108 79824 37216
rect 80422 37204 80428 37256
rect 80480 37244 80486 37256
rect 81820 37244 81848 37284
rect 82722 37272 82728 37324
rect 82780 37312 82786 37324
rect 83016 37321 83044 37420
rect 84013 37417 84025 37451
rect 84059 37448 84071 37451
rect 89714 37448 89720 37460
rect 84059 37420 89720 37448
rect 84059 37417 84071 37420
rect 84013 37411 84071 37417
rect 89714 37408 89720 37420
rect 89772 37408 89778 37460
rect 89806 37408 89812 37460
rect 89864 37448 89870 37460
rect 94222 37448 94228 37460
rect 89864 37420 89909 37448
rect 94183 37420 94228 37448
rect 89864 37408 89870 37420
rect 94222 37408 94228 37420
rect 94280 37408 94286 37460
rect 95050 37448 95056 37460
rect 95011 37420 95056 37448
rect 95050 37408 95056 37420
rect 95108 37408 95114 37460
rect 97534 37448 97540 37460
rect 97495 37420 97540 37448
rect 97534 37408 97540 37420
rect 97592 37408 97598 37460
rect 99466 37448 99472 37460
rect 99427 37420 99472 37448
rect 99466 37408 99472 37420
rect 99524 37408 99530 37460
rect 101950 37448 101956 37460
rect 101911 37420 101956 37448
rect 101950 37408 101956 37420
rect 102008 37408 102014 37460
rect 103517 37451 103575 37457
rect 103517 37417 103529 37451
rect 103563 37448 103575 37451
rect 119890 37448 119896 37460
rect 103563 37420 119896 37448
rect 103563 37417 103575 37420
rect 103517 37411 103575 37417
rect 119890 37408 119896 37420
rect 119948 37408 119954 37460
rect 120074 37448 120080 37460
rect 120035 37420 120080 37448
rect 120074 37408 120080 37420
rect 120132 37408 120138 37460
rect 120442 37408 120448 37460
rect 120500 37448 120506 37460
rect 121457 37451 121515 37457
rect 121457 37448 121469 37451
rect 120500 37420 121469 37448
rect 120500 37408 120506 37420
rect 121457 37417 121469 37420
rect 121503 37417 121515 37451
rect 122558 37448 122564 37460
rect 122519 37420 122564 37448
rect 121457 37411 121515 37417
rect 122558 37408 122564 37420
rect 122616 37408 122622 37460
rect 125870 37408 125876 37460
rect 125928 37448 125934 37460
rect 125965 37451 126023 37457
rect 125965 37448 125977 37451
rect 125928 37420 125977 37448
rect 125928 37408 125934 37420
rect 125965 37417 125977 37420
rect 126011 37417 126023 37451
rect 125965 37411 126023 37417
rect 83182 37340 83188 37392
rect 83240 37380 83246 37392
rect 136177 37383 136235 37389
rect 136177 37380 136189 37383
rect 83240 37352 136189 37380
rect 83240 37340 83246 37352
rect 136177 37349 136189 37352
rect 136223 37349 136235 37383
rect 136177 37343 136235 37349
rect 138017 37383 138075 37389
rect 138017 37349 138029 37383
rect 138063 37349 138075 37383
rect 138017 37343 138075 37349
rect 83001 37315 83059 37321
rect 82780 37284 82952 37312
rect 82780 37272 82786 37284
rect 82630 37244 82636 37256
rect 80480 37216 80525 37244
rect 81820 37216 82636 37244
rect 80480 37204 80486 37216
rect 82630 37204 82636 37216
rect 82688 37204 82694 37256
rect 82814 37244 82820 37256
rect 82775 37216 82820 37244
rect 82814 37204 82820 37216
rect 82872 37204 82878 37256
rect 82924 37244 82952 37284
rect 83001 37281 83013 37315
rect 83047 37281 83059 37315
rect 83001 37275 83059 37281
rect 83090 37272 83096 37324
rect 83148 37312 83154 37324
rect 84194 37312 84200 37324
rect 83148 37284 84200 37312
rect 83148 37272 83154 37284
rect 84194 37272 84200 37284
rect 84252 37272 84258 37324
rect 89714 37272 89720 37324
rect 89772 37312 89778 37324
rect 99466 37312 99472 37324
rect 89772 37284 99472 37312
rect 89772 37272 89778 37284
rect 99466 37272 99472 37284
rect 99524 37272 99530 37324
rect 102042 37272 102048 37324
rect 102100 37312 102106 37324
rect 105906 37312 105912 37324
rect 102100 37284 102916 37312
rect 105867 37284 105912 37312
rect 102100 37272 102106 37284
rect 102888 37256 102916 37284
rect 105906 37272 105912 37284
rect 105964 37272 105970 37324
rect 110230 37272 110236 37324
rect 110288 37312 110294 37324
rect 110325 37315 110383 37321
rect 110325 37312 110337 37315
rect 110288 37284 110337 37312
rect 110288 37272 110294 37284
rect 110325 37281 110337 37284
rect 110371 37281 110383 37315
rect 116210 37312 116216 37324
rect 116171 37284 116216 37312
rect 110325 37275 110383 37281
rect 116210 37272 116216 37284
rect 116268 37272 116274 37324
rect 118050 37312 118056 37324
rect 118011 37284 118056 37312
rect 118050 37272 118056 37284
rect 118108 37272 118114 37324
rect 120626 37312 120632 37324
rect 120587 37284 120632 37312
rect 120626 37272 120632 37284
rect 120684 37272 120690 37324
rect 123478 37272 123484 37324
rect 123536 37312 123542 37324
rect 138032 37312 138060 37343
rect 123536 37284 138060 37312
rect 139596 37284 140636 37312
rect 123536 37272 123542 37284
rect 84838 37244 84844 37256
rect 82924 37216 84844 37244
rect 84838 37204 84844 37216
rect 84896 37204 84902 37256
rect 85298 37244 85304 37256
rect 85259 37216 85304 37244
rect 85298 37204 85304 37216
rect 85356 37204 85362 37256
rect 86681 37247 86739 37253
rect 86681 37213 86693 37247
rect 86727 37244 86739 37247
rect 86770 37244 86776 37256
rect 86727 37216 86776 37244
rect 86727 37213 86739 37216
rect 86681 37207 86739 37213
rect 86770 37204 86776 37216
rect 86828 37204 86834 37256
rect 86954 37204 86960 37256
rect 87012 37244 87018 37256
rect 87417 37247 87475 37253
rect 87417 37244 87429 37247
rect 87012 37216 87429 37244
rect 87012 37204 87018 37216
rect 87417 37213 87429 37216
rect 87463 37244 87475 37247
rect 87506 37244 87512 37256
rect 87463 37216 87512 37244
rect 87463 37213 87475 37216
rect 87417 37207 87475 37213
rect 87506 37204 87512 37216
rect 87564 37204 87570 37256
rect 88058 37204 88064 37256
rect 88116 37244 88122 37256
rect 88153 37247 88211 37253
rect 88153 37244 88165 37247
rect 88116 37216 88165 37244
rect 88116 37204 88122 37216
rect 88153 37213 88165 37216
rect 88199 37213 88211 37247
rect 88153 37207 88211 37213
rect 89257 37247 89315 37253
rect 89257 37213 89269 37247
rect 89303 37244 89315 37247
rect 89622 37244 89628 37256
rect 89303 37216 89628 37244
rect 89303 37213 89315 37216
rect 89257 37207 89315 37213
rect 89622 37204 89628 37216
rect 89680 37204 89686 37256
rect 90082 37204 90088 37256
rect 90140 37244 90146 37256
rect 90726 37244 90732 37256
rect 90140 37216 90732 37244
rect 90140 37204 90146 37216
rect 90726 37204 90732 37216
rect 90784 37204 90790 37256
rect 91554 37244 91560 37256
rect 91515 37216 91560 37244
rect 91554 37204 91560 37216
rect 91612 37204 91618 37256
rect 92106 37204 92112 37256
rect 92164 37244 92170 37256
rect 92293 37247 92351 37253
rect 92293 37244 92305 37247
rect 92164 37216 92305 37244
rect 92164 37204 92170 37216
rect 92293 37213 92305 37216
rect 92339 37213 92351 37247
rect 92293 37207 92351 37213
rect 92934 37204 92940 37256
rect 92992 37244 92998 37256
rect 93029 37247 93087 37253
rect 93029 37244 93041 37247
rect 92992 37216 93041 37244
rect 92992 37204 92998 37216
rect 93029 37213 93041 37216
rect 93075 37213 93087 37247
rect 93029 37207 93087 37213
rect 93854 37204 93860 37256
rect 93912 37244 93918 37256
rect 94317 37247 94375 37253
rect 94317 37244 94329 37247
rect 93912 37216 94329 37244
rect 93912 37204 93918 37216
rect 94317 37213 94329 37216
rect 94363 37213 94375 37247
rect 94317 37207 94375 37213
rect 95881 37247 95939 37253
rect 95881 37213 95893 37247
rect 95927 37244 95939 37247
rect 96154 37244 96160 37256
rect 95927 37216 96160 37244
rect 95927 37213 95939 37216
rect 95881 37207 95939 37213
rect 96154 37204 96160 37216
rect 96212 37204 96218 37256
rect 96706 37204 96712 37256
rect 96764 37244 96770 37256
rect 96985 37247 97043 37253
rect 96985 37244 96997 37247
rect 96764 37216 96997 37244
rect 96764 37204 96770 37216
rect 96985 37213 96997 37216
rect 97031 37213 97043 37247
rect 98454 37244 98460 37256
rect 98415 37216 98460 37244
rect 96985 37207 97043 37213
rect 98454 37204 98460 37216
rect 98512 37204 98518 37256
rect 99282 37204 99288 37256
rect 99340 37244 99346 37256
rect 99834 37244 99840 37256
rect 99340 37216 99840 37244
rect 99340 37204 99346 37216
rect 99834 37204 99840 37216
rect 99892 37244 99898 37256
rect 100021 37247 100079 37253
rect 100021 37244 100033 37247
rect 99892 37216 100033 37244
rect 99892 37204 99898 37216
rect 100021 37213 100033 37216
rect 100067 37213 100079 37247
rect 100021 37207 100079 37213
rect 100570 37204 100576 37256
rect 100628 37244 100634 37256
rect 100757 37247 100815 37253
rect 100757 37244 100769 37247
rect 100628 37216 100769 37244
rect 100628 37204 100634 37216
rect 100757 37213 100769 37216
rect 100803 37213 100815 37247
rect 102778 37244 102784 37256
rect 100757 37207 100815 37213
rect 100864 37216 102784 37244
rect 81434 37136 81440 37188
rect 81492 37176 81498 37188
rect 81621 37179 81679 37185
rect 81621 37176 81633 37179
rect 81492 37148 81633 37176
rect 81492 37136 81498 37148
rect 81621 37145 81633 37148
rect 81667 37145 81679 37179
rect 81621 37139 81679 37145
rect 82262 37136 82268 37188
rect 82320 37176 82326 37188
rect 83918 37176 83924 37188
rect 82320 37148 83924 37176
rect 82320 37136 82326 37148
rect 83918 37136 83924 37148
rect 83976 37136 83982 37188
rect 84562 37136 84568 37188
rect 84620 37176 84626 37188
rect 89901 37179 89959 37185
rect 84620 37148 85528 37176
rect 84620 37136 84626 37148
rect 80790 37108 80796 37120
rect 79796 37080 80796 37108
rect 80790 37068 80796 37080
rect 80848 37068 80854 37120
rect 81802 37068 81808 37120
rect 81860 37108 81866 37120
rect 81989 37111 82047 37117
rect 81989 37108 82001 37111
rect 81860 37080 82001 37108
rect 81860 37068 81866 37080
rect 81989 37077 82001 37080
rect 82035 37077 82047 37111
rect 82446 37108 82452 37120
rect 82407 37080 82452 37108
rect 81989 37071 82047 37077
rect 82446 37068 82452 37080
rect 82504 37068 82510 37120
rect 82909 37111 82967 37117
rect 82909 37077 82921 37111
rect 82955 37108 82967 37111
rect 83090 37108 83096 37120
rect 82955 37080 83096 37108
rect 82955 37077 82967 37080
rect 82909 37071 82967 37077
rect 83090 37068 83096 37080
rect 83148 37068 83154 37120
rect 84654 37108 84660 37120
rect 84615 37080 84660 37108
rect 84654 37068 84660 37080
rect 84712 37068 84718 37120
rect 85500 37117 85528 37148
rect 89901 37145 89913 37179
rect 89947 37176 89959 37179
rect 90358 37176 90364 37188
rect 89947 37148 90364 37176
rect 89947 37145 89959 37148
rect 89901 37139 89959 37145
rect 90358 37136 90364 37148
rect 90416 37136 90422 37188
rect 94961 37179 95019 37185
rect 94961 37176 94973 37179
rect 94332 37148 94973 37176
rect 94332 37120 94360 37148
rect 94961 37145 94973 37148
rect 95007 37145 95019 37179
rect 94961 37139 95019 37145
rect 97629 37179 97687 37185
rect 97629 37145 97641 37179
rect 97675 37176 97687 37179
rect 97810 37176 97816 37188
rect 97675 37148 97816 37176
rect 97675 37145 97687 37148
rect 97629 37139 97687 37145
rect 97810 37136 97816 37148
rect 97868 37176 97874 37188
rect 98730 37176 98736 37188
rect 97868 37148 98736 37176
rect 97868 37136 97874 37148
rect 98730 37136 98736 37148
rect 98788 37136 98794 37188
rect 99374 37176 99380 37188
rect 99335 37148 99380 37176
rect 99374 37136 99380 37148
rect 99432 37136 99438 37188
rect 100864 37176 100892 37216
rect 102778 37204 102784 37216
rect 102836 37204 102842 37256
rect 102870 37204 102876 37256
rect 102928 37244 102934 37256
rect 104434 37244 104440 37256
rect 102928 37216 103021 37244
rect 104395 37216 104440 37244
rect 102928 37204 102934 37216
rect 104434 37204 104440 37216
rect 104492 37204 104498 37256
rect 104894 37204 104900 37256
rect 104952 37244 104958 37256
rect 105173 37247 105231 37253
rect 105173 37244 105185 37247
rect 104952 37216 105185 37244
rect 104952 37204 104958 37216
rect 105173 37213 105185 37216
rect 105219 37213 105231 37247
rect 105173 37207 105231 37213
rect 105280 37216 106228 37244
rect 99484 37148 100892 37176
rect 102045 37179 102103 37185
rect 85485 37111 85543 37117
rect 85485 37077 85497 37111
rect 85531 37077 85543 37111
rect 85485 37071 85543 37077
rect 85574 37068 85580 37120
rect 85632 37108 85638 37120
rect 86497 37111 86555 37117
rect 86497 37108 86509 37111
rect 85632 37080 86509 37108
rect 85632 37068 85638 37080
rect 86497 37077 86509 37080
rect 86543 37077 86555 37111
rect 87230 37108 87236 37120
rect 87191 37080 87236 37108
rect 86497 37071 86555 37077
rect 87230 37068 87236 37080
rect 87288 37068 87294 37120
rect 87322 37068 87328 37120
rect 87380 37108 87386 37120
rect 87969 37111 88027 37117
rect 87969 37108 87981 37111
rect 87380 37080 87981 37108
rect 87380 37068 87386 37080
rect 87969 37077 87981 37080
rect 88015 37077 88027 37111
rect 87969 37071 88027 37077
rect 88334 37068 88340 37120
rect 88392 37108 88398 37120
rect 89073 37111 89131 37117
rect 89073 37108 89085 37111
rect 88392 37080 89085 37108
rect 88392 37068 88398 37080
rect 89073 37077 89085 37080
rect 89119 37077 89131 37111
rect 89073 37071 89131 37077
rect 89254 37068 89260 37120
rect 89312 37108 89318 37120
rect 90545 37111 90603 37117
rect 90545 37108 90557 37111
rect 89312 37080 90557 37108
rect 89312 37068 89318 37080
rect 90545 37077 90557 37080
rect 90591 37077 90603 37111
rect 90545 37071 90603 37077
rect 91094 37068 91100 37120
rect 91152 37108 91158 37120
rect 91741 37111 91799 37117
rect 91741 37108 91753 37111
rect 91152 37080 91753 37108
rect 91152 37068 91158 37080
rect 91741 37077 91753 37080
rect 91787 37077 91799 37111
rect 91741 37071 91799 37077
rect 91922 37068 91928 37120
rect 91980 37108 91986 37120
rect 92477 37111 92535 37117
rect 92477 37108 92489 37111
rect 91980 37080 92489 37108
rect 91980 37068 91986 37080
rect 92477 37077 92489 37080
rect 92523 37077 92535 37111
rect 92477 37071 92535 37077
rect 92842 37068 92848 37120
rect 92900 37108 92906 37120
rect 93213 37111 93271 37117
rect 93213 37108 93225 37111
rect 92900 37080 93225 37108
rect 92900 37068 92906 37080
rect 93213 37077 93225 37080
rect 93259 37077 93271 37111
rect 93213 37071 93271 37077
rect 94314 37068 94320 37120
rect 94372 37068 94378 37120
rect 95234 37068 95240 37120
rect 95292 37108 95298 37120
rect 95697 37111 95755 37117
rect 95697 37108 95709 37111
rect 95292 37080 95709 37108
rect 95292 37068 95298 37080
rect 95697 37077 95709 37080
rect 95743 37077 95755 37111
rect 96798 37108 96804 37120
rect 96759 37080 96804 37108
rect 95697 37071 95755 37077
rect 96798 37068 96804 37080
rect 96856 37068 96862 37120
rect 97994 37068 98000 37120
rect 98052 37108 98058 37120
rect 98273 37111 98331 37117
rect 98273 37108 98285 37111
rect 98052 37080 98285 37108
rect 98052 37068 98058 37080
rect 98273 37077 98285 37080
rect 98319 37077 98331 37111
rect 98273 37071 98331 37077
rect 98546 37068 98552 37120
rect 98604 37108 98610 37120
rect 99484 37108 99512 37148
rect 102045 37145 102057 37179
rect 102091 37176 102103 37179
rect 102134 37176 102140 37188
rect 102091 37148 102140 37176
rect 102091 37145 102103 37148
rect 102045 37139 102103 37145
rect 102134 37136 102140 37148
rect 102192 37176 102198 37188
rect 103422 37176 103428 37188
rect 102192 37148 103428 37176
rect 102192 37136 102198 37148
rect 103422 37136 103428 37148
rect 103480 37136 103486 37188
rect 105280 37176 105308 37216
rect 103808 37148 105308 37176
rect 106093 37179 106151 37185
rect 100202 37108 100208 37120
rect 98604 37080 99512 37108
rect 100163 37080 100208 37108
rect 98604 37068 98610 37080
rect 100202 37068 100208 37080
rect 100260 37068 100266 37120
rect 100754 37068 100760 37120
rect 100812 37108 100818 37120
rect 100941 37111 100999 37117
rect 100941 37108 100953 37111
rect 100812 37080 100953 37108
rect 100812 37068 100818 37080
rect 100941 37077 100953 37080
rect 100987 37077 100999 37111
rect 102686 37108 102692 37120
rect 102647 37080 102692 37108
rect 100941 37071 100999 37077
rect 102686 37068 102692 37080
rect 102744 37068 102750 37120
rect 102778 37068 102784 37120
rect 102836 37108 102842 37120
rect 103808 37108 103836 37148
rect 106093 37145 106105 37179
rect 106139 37145 106151 37179
rect 106200 37176 106228 37216
rect 106642 37204 106648 37256
rect 106700 37244 106706 37256
rect 107286 37244 107292 37256
rect 106700 37216 107292 37244
rect 106700 37204 106706 37216
rect 107286 37204 107292 37216
rect 107344 37204 107350 37256
rect 107746 37244 107752 37256
rect 107707 37216 107752 37244
rect 107746 37204 107752 37216
rect 107804 37204 107810 37256
rect 108482 37204 108488 37256
rect 108540 37244 108546 37256
rect 108577 37247 108635 37253
rect 108577 37244 108589 37247
rect 108540 37216 108589 37244
rect 108540 37204 108546 37216
rect 108577 37213 108589 37216
rect 108623 37213 108635 37247
rect 109586 37244 109592 37256
rect 109547 37216 109592 37244
rect 108577 37207 108635 37213
rect 109586 37204 109592 37216
rect 109644 37204 109650 37256
rect 110432 37216 110644 37244
rect 110432 37176 110460 37216
rect 106200 37148 110460 37176
rect 110509 37179 110567 37185
rect 106093 37139 106151 37145
rect 110509 37145 110521 37179
rect 110555 37145 110567 37179
rect 110616 37176 110644 37216
rect 110690 37204 110696 37256
rect 110748 37244 110754 37256
rect 111061 37247 111119 37253
rect 111061 37244 111073 37247
rect 110748 37216 111073 37244
rect 110748 37204 110754 37216
rect 111061 37213 111073 37216
rect 111107 37213 111119 37247
rect 112162 37244 112168 37256
rect 112123 37216 112168 37244
rect 111061 37207 111119 37213
rect 112162 37204 112168 37216
rect 112220 37204 112226 37256
rect 112254 37204 112260 37256
rect 112312 37244 112318 37256
rect 112714 37244 112720 37256
rect 112312 37216 112720 37244
rect 112312 37204 112318 37216
rect 112714 37204 112720 37216
rect 112772 37244 112778 37256
rect 112901 37247 112959 37253
rect 112901 37244 112913 37247
rect 112772 37216 112913 37244
rect 112772 37204 112778 37216
rect 112901 37213 112913 37216
rect 112947 37213 112959 37247
rect 112901 37207 112959 37213
rect 113450 37204 113456 37256
rect 113508 37244 113514 37256
rect 113637 37247 113695 37253
rect 113637 37244 113649 37247
rect 113508 37216 113649 37244
rect 113508 37204 113514 37216
rect 113637 37213 113649 37216
rect 113683 37213 113695 37247
rect 113637 37207 113695 37213
rect 114002 37204 114008 37256
rect 114060 37244 114066 37256
rect 114741 37247 114799 37253
rect 114741 37244 114753 37247
rect 114060 37216 114753 37244
rect 114060 37204 114066 37216
rect 114741 37213 114753 37216
rect 114787 37244 114799 37247
rect 114830 37244 114836 37256
rect 114787 37216 114836 37244
rect 114787 37213 114799 37216
rect 114741 37207 114799 37213
rect 114830 37204 114836 37216
rect 114888 37204 114894 37256
rect 115474 37244 115480 37256
rect 115435 37216 115480 37244
rect 115474 37204 115480 37216
rect 115532 37204 115538 37256
rect 115934 37204 115940 37256
rect 115992 37244 115998 37256
rect 116118 37244 116124 37256
rect 115992 37216 116124 37244
rect 115992 37204 115998 37216
rect 116118 37204 116124 37216
rect 116176 37244 116182 37256
rect 116397 37247 116455 37253
rect 116397 37244 116409 37247
rect 116176 37216 116409 37244
rect 116176 37204 116182 37216
rect 116397 37213 116409 37216
rect 116443 37213 116455 37247
rect 116397 37207 116455 37213
rect 117130 37204 117136 37256
rect 117188 37244 117194 37256
rect 117317 37247 117375 37253
rect 117317 37244 117329 37247
rect 117188 37216 117329 37244
rect 117188 37204 117194 37216
rect 117317 37213 117329 37216
rect 117363 37213 117375 37247
rect 119065 37247 119123 37253
rect 117317 37207 117375 37213
rect 117424 37216 118694 37244
rect 117424 37176 117452 37216
rect 110616 37148 117452 37176
rect 110509 37139 110567 37145
rect 102836 37080 103836 37108
rect 102836 37068 102842 37080
rect 103882 37068 103888 37120
rect 103940 37108 103946 37120
rect 104621 37111 104679 37117
rect 104621 37108 104633 37111
rect 103940 37080 104633 37108
rect 103940 37068 103946 37080
rect 104621 37077 104633 37080
rect 104667 37077 104679 37111
rect 105354 37108 105360 37120
rect 105315 37080 105360 37108
rect 104621 37071 104679 37077
rect 105354 37068 105360 37080
rect 105412 37068 105418 37120
rect 106108 37108 106136 37139
rect 106550 37108 106556 37120
rect 106108 37080 106556 37108
rect 106550 37068 106556 37080
rect 106608 37068 106614 37120
rect 107102 37108 107108 37120
rect 107063 37080 107108 37108
rect 107102 37068 107108 37080
rect 107160 37068 107166 37120
rect 107654 37068 107660 37120
rect 107712 37108 107718 37120
rect 107933 37111 107991 37117
rect 107933 37108 107945 37111
rect 107712 37080 107945 37108
rect 107712 37068 107718 37080
rect 107933 37077 107945 37080
rect 107979 37077 107991 37111
rect 108758 37108 108764 37120
rect 108719 37080 108764 37108
rect 107933 37071 107991 37077
rect 108758 37068 108764 37080
rect 108816 37068 108822 37120
rect 109402 37068 109408 37120
rect 109460 37108 109466 37120
rect 109773 37111 109831 37117
rect 109773 37108 109785 37111
rect 109460 37080 109785 37108
rect 109460 37068 109466 37080
rect 109773 37077 109785 37080
rect 109819 37077 109831 37111
rect 109773 37071 109831 37077
rect 110414 37068 110420 37120
rect 110472 37108 110478 37120
rect 110522 37108 110550 37139
rect 117682 37136 117688 37188
rect 117740 37176 117746 37188
rect 118237 37179 118295 37185
rect 118237 37176 118249 37179
rect 117740 37148 118249 37176
rect 117740 37136 117746 37148
rect 118237 37145 118249 37148
rect 118283 37145 118295 37179
rect 118666 37176 118694 37216
rect 119065 37213 119077 37247
rect 119111 37244 119123 37247
rect 119154 37244 119160 37256
rect 119111 37216 119160 37244
rect 119111 37213 119123 37216
rect 119065 37207 119123 37213
rect 119154 37204 119160 37216
rect 119212 37204 119218 37256
rect 119522 37204 119528 37256
rect 119580 37244 119586 37256
rect 119890 37244 119896 37256
rect 119580 37216 119896 37244
rect 119580 37204 119586 37216
rect 119890 37204 119896 37216
rect 119948 37204 119954 37256
rect 121641 37247 121699 37253
rect 120000 37216 121592 37244
rect 120000 37176 120028 37216
rect 120810 37176 120816 37188
rect 118666 37148 120028 37176
rect 120771 37148 120816 37176
rect 118237 37139 118295 37145
rect 120810 37136 120816 37148
rect 120868 37136 120874 37188
rect 121564 37176 121592 37216
rect 121641 37213 121653 37247
rect 121687 37244 121699 37247
rect 121730 37244 121736 37256
rect 121687 37216 121736 37244
rect 121687 37213 121699 37216
rect 121641 37207 121699 37213
rect 121730 37204 121736 37216
rect 121788 37204 121794 37256
rect 122745 37247 122803 37253
rect 122745 37213 122757 37247
rect 122791 37244 122803 37247
rect 122926 37244 122932 37256
rect 122791 37216 122932 37244
rect 122791 37213 122803 37216
rect 122745 37207 122803 37213
rect 122926 37204 122932 37216
rect 122984 37204 122990 37256
rect 123110 37204 123116 37256
rect 123168 37244 123174 37256
rect 123205 37247 123263 37253
rect 123205 37244 123217 37247
rect 123168 37216 123217 37244
rect 123168 37204 123174 37216
rect 123205 37213 123217 37216
rect 123251 37213 123263 37247
rect 123205 37207 123263 37213
rect 123294 37204 123300 37256
rect 123352 37244 123358 37256
rect 124217 37247 124275 37253
rect 124217 37244 124229 37247
rect 123352 37216 124229 37244
rect 123352 37204 123358 37216
rect 124217 37213 124229 37216
rect 124263 37244 124275 37247
rect 124398 37244 124404 37256
rect 124263 37216 124404 37244
rect 124263 37213 124275 37216
rect 124217 37207 124275 37213
rect 124398 37204 124404 37216
rect 124456 37204 124462 37256
rect 124950 37204 124956 37256
rect 125008 37244 125014 37256
rect 125045 37247 125103 37253
rect 125045 37244 125057 37247
rect 125008 37216 125057 37244
rect 125008 37204 125014 37216
rect 125045 37213 125057 37216
rect 125091 37213 125103 37247
rect 125045 37207 125103 37213
rect 125134 37204 125140 37256
rect 125192 37244 125198 37256
rect 125594 37244 125600 37256
rect 125192 37216 125600 37244
rect 125192 37204 125198 37216
rect 125594 37204 125600 37216
rect 125652 37244 125658 37256
rect 125781 37247 125839 37253
rect 125781 37244 125793 37247
rect 125652 37216 125793 37244
rect 125652 37204 125658 37216
rect 125781 37213 125793 37216
rect 125827 37213 125839 37247
rect 125781 37207 125839 37213
rect 126422 37204 126428 37256
rect 126480 37244 126486 37256
rect 126517 37247 126575 37253
rect 126517 37244 126529 37247
rect 126480 37216 126529 37244
rect 126480 37204 126486 37216
rect 126517 37213 126529 37216
rect 126563 37213 126575 37247
rect 126517 37207 126575 37213
rect 126974 37204 126980 37256
rect 127032 37244 127038 37256
rect 127621 37247 127679 37253
rect 127621 37244 127633 37247
rect 127032 37216 127633 37244
rect 127032 37204 127038 37216
rect 127621 37213 127633 37216
rect 127667 37244 127679 37247
rect 127710 37244 127716 37256
rect 127667 37216 127716 37244
rect 127667 37213 127679 37216
rect 127621 37207 127679 37213
rect 127710 37204 127716 37216
rect 127768 37204 127774 37256
rect 128357 37247 128415 37253
rect 128357 37213 128369 37247
rect 128403 37244 128415 37247
rect 128446 37244 128452 37256
rect 128403 37216 128452 37244
rect 128403 37213 128415 37216
rect 128357 37207 128415 37213
rect 128446 37204 128452 37216
rect 128504 37204 128510 37256
rect 128722 37204 128728 37256
rect 128780 37244 128786 37256
rect 129093 37247 129151 37253
rect 129093 37244 129105 37247
rect 128780 37216 129105 37244
rect 128780 37204 128786 37216
rect 129093 37213 129105 37216
rect 129139 37213 129151 37247
rect 129093 37207 129151 37213
rect 129550 37204 129556 37256
rect 129608 37244 129614 37256
rect 130197 37247 130255 37253
rect 130197 37244 130209 37247
rect 129608 37216 130209 37244
rect 129608 37204 129614 37216
rect 130197 37213 130209 37216
rect 130243 37213 130255 37247
rect 130197 37207 130255 37213
rect 131114 37204 131120 37256
rect 131172 37244 131178 37256
rect 131209 37247 131267 37253
rect 131209 37244 131221 37247
rect 131172 37216 131221 37244
rect 131172 37204 131178 37216
rect 131209 37213 131221 37216
rect 131255 37213 131267 37247
rect 131666 37244 131672 37256
rect 131627 37216 131672 37244
rect 131209 37207 131267 37213
rect 131666 37204 131672 37216
rect 131724 37204 131730 37256
rect 132494 37204 132500 37256
rect 132552 37244 132558 37256
rect 133049 37247 133107 37253
rect 133049 37244 133061 37247
rect 132552 37216 133061 37244
rect 132552 37204 132558 37216
rect 133049 37213 133061 37216
rect 133095 37244 133107 37247
rect 133230 37244 133236 37256
rect 133095 37216 133236 37244
rect 133095 37213 133107 37216
rect 133049 37207 133107 37213
rect 133230 37204 133236 37216
rect 133288 37204 133294 37256
rect 133506 37244 133512 37256
rect 133467 37216 133512 37244
rect 133506 37204 133512 37216
rect 133564 37204 133570 37256
rect 134242 37204 134248 37256
rect 134300 37244 134306 37256
rect 134337 37247 134395 37253
rect 134337 37244 134349 37247
rect 134300 37216 134349 37244
rect 134300 37204 134306 37216
rect 134337 37213 134349 37216
rect 134383 37213 134395 37247
rect 134337 37207 134395 37213
rect 134426 37204 134432 37256
rect 134484 37244 134490 37256
rect 135349 37247 135407 37253
rect 135349 37244 135361 37247
rect 134484 37216 135361 37244
rect 134484 37204 134490 37216
rect 135349 37213 135361 37216
rect 135395 37213 135407 37247
rect 135349 37207 135407 37213
rect 135990 37204 135996 37256
rect 136048 37244 136054 37256
rect 137097 37247 137155 37253
rect 137097 37244 137109 37247
rect 136048 37216 137109 37244
rect 136048 37204 136054 37216
rect 137097 37213 137109 37216
rect 137143 37213 137155 37247
rect 137097 37207 137155 37213
rect 138014 37204 138020 37256
rect 138072 37244 138078 37256
rect 138201 37247 138259 37253
rect 138201 37244 138213 37247
rect 138072 37216 138213 37244
rect 138072 37204 138078 37216
rect 138201 37213 138213 37216
rect 138247 37213 138259 37247
rect 138934 37244 138940 37256
rect 138895 37216 138940 37244
rect 138201 37207 138259 37213
rect 138934 37204 138940 37216
rect 138992 37204 138998 37256
rect 121564 37148 136036 37176
rect 111242 37108 111248 37120
rect 110472 37080 110550 37108
rect 111203 37080 111248 37108
rect 110472 37068 110478 37080
rect 111242 37068 111248 37080
rect 111300 37068 111306 37120
rect 111794 37068 111800 37120
rect 111852 37108 111858 37120
rect 112349 37111 112407 37117
rect 112349 37108 112361 37111
rect 111852 37080 112361 37108
rect 111852 37068 111858 37080
rect 112349 37077 112361 37080
rect 112395 37077 112407 37111
rect 112349 37071 112407 37077
rect 112990 37068 112996 37120
rect 113048 37108 113054 37120
rect 113085 37111 113143 37117
rect 113085 37108 113097 37111
rect 113048 37080 113097 37108
rect 113048 37068 113054 37080
rect 113085 37077 113097 37080
rect 113131 37077 113143 37111
rect 113085 37071 113143 37077
rect 113174 37068 113180 37120
rect 113232 37108 113238 37120
rect 113821 37111 113879 37117
rect 113821 37108 113833 37111
rect 113232 37080 113833 37108
rect 113232 37068 113238 37080
rect 113821 37077 113833 37080
rect 113867 37077 113879 37111
rect 113821 37071 113879 37077
rect 114554 37068 114560 37120
rect 114612 37108 114618 37120
rect 114925 37111 114983 37117
rect 114925 37108 114937 37111
rect 114612 37080 114937 37108
rect 114612 37068 114618 37080
rect 114925 37077 114937 37080
rect 114971 37077 114983 37111
rect 114925 37071 114983 37077
rect 115014 37068 115020 37120
rect 115072 37108 115078 37120
rect 115661 37111 115719 37117
rect 115661 37108 115673 37111
rect 115072 37080 115673 37108
rect 115072 37068 115078 37080
rect 115661 37077 115673 37080
rect 115707 37077 115719 37111
rect 115661 37071 115719 37077
rect 117314 37068 117320 37120
rect 117372 37108 117378 37120
rect 117501 37111 117559 37117
rect 117501 37108 117513 37111
rect 117372 37080 117513 37108
rect 117372 37068 117378 37080
rect 117501 37077 117513 37080
rect 117547 37077 117559 37111
rect 117501 37071 117559 37077
rect 118694 37068 118700 37120
rect 118752 37108 118758 37120
rect 118881 37111 118939 37117
rect 118881 37108 118893 37111
rect 118752 37080 118893 37108
rect 118752 37068 118758 37080
rect 118881 37077 118893 37080
rect 118927 37077 118939 37111
rect 118881 37071 118939 37077
rect 122834 37068 122840 37120
rect 122892 37108 122898 37120
rect 123389 37111 123447 37117
rect 123389 37108 123401 37111
rect 122892 37080 123401 37108
rect 122892 37068 122898 37080
rect 123389 37077 123401 37080
rect 123435 37077 123447 37111
rect 124030 37108 124036 37120
rect 123991 37080 124036 37108
rect 123389 37071 123447 37077
rect 124030 37068 124036 37080
rect 124088 37068 124094 37120
rect 124214 37068 124220 37120
rect 124272 37108 124278 37120
rect 125229 37111 125287 37117
rect 125229 37108 125241 37111
rect 124272 37080 125241 37108
rect 124272 37068 124278 37080
rect 125229 37077 125241 37080
rect 125275 37077 125287 37111
rect 125229 37071 125287 37077
rect 126054 37068 126060 37120
rect 126112 37108 126118 37120
rect 126701 37111 126759 37117
rect 126701 37108 126713 37111
rect 126112 37080 126713 37108
rect 126112 37068 126118 37080
rect 126701 37077 126713 37080
rect 126747 37077 126759 37111
rect 127802 37108 127808 37120
rect 127763 37080 127808 37108
rect 126701 37071 126759 37077
rect 127802 37068 127808 37080
rect 127860 37068 127866 37120
rect 128354 37068 128360 37120
rect 128412 37108 128418 37120
rect 128541 37111 128599 37117
rect 128541 37108 128553 37111
rect 128412 37080 128553 37108
rect 128412 37068 128418 37080
rect 128541 37077 128553 37080
rect 128587 37077 128599 37111
rect 129274 37108 129280 37120
rect 129235 37080 129280 37108
rect 128541 37071 128599 37077
rect 129274 37068 129280 37080
rect 129332 37068 129338 37120
rect 129734 37068 129740 37120
rect 129792 37108 129798 37120
rect 130381 37111 130439 37117
rect 130381 37108 130393 37111
rect 129792 37080 130393 37108
rect 129792 37068 129798 37080
rect 130381 37077 130393 37080
rect 130427 37077 130439 37111
rect 130381 37071 130439 37077
rect 130470 37068 130476 37120
rect 130528 37108 130534 37120
rect 131025 37111 131083 37117
rect 131025 37108 131037 37111
rect 130528 37080 131037 37108
rect 130528 37068 130534 37080
rect 131025 37077 131037 37080
rect 131071 37077 131083 37111
rect 131025 37071 131083 37077
rect 131482 37068 131488 37120
rect 131540 37108 131546 37120
rect 131853 37111 131911 37117
rect 131853 37108 131865 37111
rect 131540 37080 131865 37108
rect 131540 37068 131546 37080
rect 131853 37077 131865 37080
rect 131899 37077 131911 37111
rect 132862 37108 132868 37120
rect 132823 37080 132868 37108
rect 131853 37071 131911 37077
rect 132862 37068 132868 37080
rect 132920 37068 132926 37120
rect 133322 37068 133328 37120
rect 133380 37108 133386 37120
rect 133693 37111 133751 37117
rect 133693 37108 133705 37111
rect 133380 37080 133705 37108
rect 133380 37068 133386 37080
rect 133693 37077 133705 37080
rect 133739 37077 133751 37111
rect 134518 37108 134524 37120
rect 134479 37080 134524 37108
rect 133693 37071 133751 37077
rect 134518 37068 134524 37080
rect 134576 37068 134582 37120
rect 135530 37108 135536 37120
rect 135491 37080 135536 37108
rect 135530 37068 135536 37080
rect 135588 37068 135594 37120
rect 136008 37108 136036 37148
rect 136082 37136 136088 37188
rect 136140 37176 136146 37188
rect 136361 37179 136419 37185
rect 136361 37176 136373 37179
rect 136140 37148 136373 37176
rect 136140 37136 136146 37148
rect 136361 37145 136373 37148
rect 136407 37145 136419 37179
rect 139596 37176 139624 37284
rect 139673 37247 139731 37253
rect 139673 37213 139685 37247
rect 139719 37213 139731 37247
rect 139673 37207 139731 37213
rect 136361 37139 136419 37145
rect 136468 37148 139624 37176
rect 136468 37108 136496 37148
rect 136008 37080 136496 37108
rect 137002 37068 137008 37120
rect 137060 37108 137066 37120
rect 137281 37111 137339 37117
rect 137281 37108 137293 37111
rect 137060 37080 137293 37108
rect 137060 37068 137066 37080
rect 137281 37077 137293 37080
rect 137327 37077 137339 37111
rect 137281 37071 137339 37077
rect 138842 37068 138848 37120
rect 138900 37108 138906 37120
rect 139121 37111 139179 37117
rect 139121 37108 139133 37111
rect 138900 37080 139133 37108
rect 138900 37068 138906 37080
rect 139121 37077 139133 37080
rect 139167 37077 139179 37111
rect 139121 37071 139179 37077
rect 139486 37068 139492 37120
rect 139544 37108 139550 37120
rect 139688 37108 139716 37207
rect 139762 37204 139768 37256
rect 139820 37244 139826 37256
rect 140498 37244 140504 37256
rect 139820 37216 140504 37244
rect 139820 37204 139826 37216
rect 140498 37204 140504 37216
rect 140556 37204 140562 37256
rect 140608 37244 140636 37284
rect 141160 37284 141372 37312
rect 141160 37244 141188 37284
rect 140608 37216 141188 37244
rect 141237 37247 141295 37253
rect 141237 37213 141249 37247
rect 141283 37213 141295 37247
rect 141237 37207 141295 37213
rect 141252 37176 141280 37207
rect 139872 37148 141280 37176
rect 141344 37176 141372 37284
rect 141602 37204 141608 37256
rect 141660 37244 141666 37256
rect 142246 37244 142252 37256
rect 141660 37216 142252 37244
rect 141660 37204 141666 37216
rect 142246 37204 142252 37216
rect 142304 37204 142310 37256
rect 143074 37244 143080 37256
rect 143035 37216 143080 37244
rect 143074 37204 143080 37216
rect 143132 37204 143138 37256
rect 143534 37204 143540 37256
rect 143592 37244 143598 37256
rect 143813 37247 143871 37253
rect 143813 37244 143825 37247
rect 143592 37216 143825 37244
rect 143592 37204 143598 37216
rect 143813 37213 143825 37216
rect 143859 37213 143871 37247
rect 144546 37244 144552 37256
rect 144507 37216 144552 37244
rect 143813 37207 143871 37213
rect 144546 37204 144552 37216
rect 144604 37204 144610 37256
rect 145282 37204 145288 37256
rect 145340 37244 145346 37256
rect 145653 37247 145711 37253
rect 145653 37244 145665 37247
rect 145340 37216 145665 37244
rect 145340 37204 145346 37216
rect 145653 37213 145665 37216
rect 145699 37213 145711 37247
rect 145653 37207 145711 37213
rect 146294 37204 146300 37256
rect 146352 37244 146358 37256
rect 146389 37247 146447 37253
rect 146389 37244 146401 37247
rect 146352 37216 146401 37244
rect 146352 37204 146358 37216
rect 146389 37213 146401 37216
rect 146435 37213 146447 37247
rect 146389 37207 146447 37213
rect 147122 37204 147128 37256
rect 147180 37244 147186 37256
rect 147217 37247 147275 37253
rect 147217 37244 147229 37247
rect 147180 37216 147229 37244
rect 147180 37204 147186 37216
rect 147217 37213 147229 37216
rect 147263 37213 147275 37247
rect 147217 37207 147275 37213
rect 141344 37148 142108 37176
rect 139872 37117 139900 37148
rect 139544 37080 139716 37108
rect 139857 37111 139915 37117
rect 139544 37068 139550 37080
rect 139857 37077 139869 37111
rect 139903 37077 139915 37111
rect 140682 37108 140688 37120
rect 140643 37080 140688 37108
rect 139857 37071 139915 37077
rect 140682 37068 140688 37080
rect 140740 37068 140746 37120
rect 140774 37068 140780 37120
rect 140832 37108 140838 37120
rect 142080 37117 142108 37148
rect 142154 37136 142160 37188
rect 142212 37176 142218 37188
rect 142212 37148 145880 37176
rect 142212 37136 142218 37148
rect 141421 37111 141479 37117
rect 141421 37108 141433 37111
rect 140832 37080 141433 37108
rect 140832 37068 140838 37080
rect 141421 37077 141433 37080
rect 141467 37077 141479 37111
rect 141421 37071 141479 37077
rect 142065 37111 142123 37117
rect 142065 37077 142077 37111
rect 142111 37077 142123 37111
rect 142065 37071 142123 37077
rect 142522 37068 142528 37120
rect 142580 37108 142586 37120
rect 143261 37111 143319 37117
rect 143261 37108 143273 37111
rect 142580 37080 143273 37108
rect 142580 37068 142586 37080
rect 143261 37077 143273 37080
rect 143307 37077 143319 37111
rect 143994 37108 144000 37120
rect 143955 37080 144000 37108
rect 143261 37071 143319 37077
rect 143994 37068 144000 37080
rect 144052 37068 144058 37120
rect 144362 37068 144368 37120
rect 144420 37108 144426 37120
rect 145852 37117 145880 37148
rect 144733 37111 144791 37117
rect 144733 37108 144745 37111
rect 144420 37080 144745 37108
rect 144420 37068 144426 37080
rect 144733 37077 144745 37080
rect 144779 37077 144791 37111
rect 144733 37071 144791 37077
rect 145837 37111 145895 37117
rect 145837 37077 145849 37111
rect 145883 37077 145895 37111
rect 145837 37071 145895 37077
rect 146202 37068 146208 37120
rect 146260 37108 146266 37120
rect 146573 37111 146631 37117
rect 146573 37108 146585 37111
rect 146260 37080 146585 37108
rect 146260 37068 146266 37080
rect 146573 37077 146585 37080
rect 146619 37077 146631 37111
rect 147398 37108 147404 37120
rect 147359 37080 147404 37108
rect 146573 37071 146631 37077
rect 147398 37068 147404 37080
rect 147456 37068 147462 37120
rect 1104 37018 148856 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 81014 37018
rect 81066 36966 81078 37018
rect 81130 36966 81142 37018
rect 81194 36966 81206 37018
rect 81258 36966 81270 37018
rect 81322 36966 111734 37018
rect 111786 36966 111798 37018
rect 111850 36966 111862 37018
rect 111914 36966 111926 37018
rect 111978 36966 111990 37018
rect 112042 36966 142454 37018
rect 142506 36966 142518 37018
rect 142570 36966 142582 37018
rect 142634 36966 142646 37018
rect 142698 36966 142710 37018
rect 142762 36966 148856 37018
rect 1104 36944 148856 36966
rect 3602 36864 3608 36916
rect 3660 36904 3666 36916
rect 3789 36907 3847 36913
rect 3789 36904 3801 36907
rect 3660 36876 3801 36904
rect 3660 36864 3666 36876
rect 3789 36873 3801 36876
rect 3835 36873 3847 36907
rect 4522 36904 4528 36916
rect 4483 36876 4528 36904
rect 3789 36867 3847 36873
rect 4522 36864 4528 36876
rect 4580 36864 4586 36916
rect 8202 36904 8208 36916
rect 8163 36876 8208 36904
rect 8202 36864 8208 36876
rect 8260 36864 8266 36916
rect 9766 36904 9772 36916
rect 9727 36876 9772 36904
rect 9766 36864 9772 36876
rect 9824 36864 9830 36916
rect 12250 36864 12256 36916
rect 12308 36904 12314 36916
rect 12437 36907 12495 36913
rect 12437 36904 12449 36907
rect 12308 36876 12449 36904
rect 12308 36864 12314 36876
rect 12437 36873 12449 36876
rect 12483 36904 12495 36907
rect 16574 36904 16580 36916
rect 12483 36876 16580 36904
rect 12483 36873 12495 36876
rect 12437 36867 12495 36873
rect 16574 36864 16580 36876
rect 16632 36864 16638 36916
rect 17310 36904 17316 36916
rect 17271 36876 17316 36904
rect 17310 36864 17316 36876
rect 17368 36864 17374 36916
rect 19058 36904 19064 36916
rect 19019 36876 19064 36904
rect 19058 36864 19064 36876
rect 19116 36864 19122 36916
rect 19150 36864 19156 36916
rect 19208 36904 19214 36916
rect 20438 36904 20444 36916
rect 19208 36876 20444 36904
rect 19208 36864 19214 36876
rect 20438 36864 20444 36876
rect 20496 36864 20502 36916
rect 20622 36904 20628 36916
rect 20583 36876 20628 36904
rect 20622 36864 20628 36876
rect 20680 36864 20686 36916
rect 28350 36904 28356 36916
rect 28311 36876 28356 36904
rect 28350 36864 28356 36876
rect 28408 36864 28414 36916
rect 28442 36864 28448 36916
rect 28500 36904 28506 36916
rect 28905 36907 28963 36913
rect 28905 36904 28917 36907
rect 28500 36876 28917 36904
rect 28500 36864 28506 36876
rect 28905 36873 28917 36876
rect 28951 36873 28963 36907
rect 29641 36907 29699 36913
rect 29641 36904 29653 36907
rect 28905 36867 28963 36873
rect 29012 36876 29653 36904
rect 3973 36771 4031 36777
rect 3973 36737 3985 36771
rect 4019 36768 4031 36771
rect 4540 36768 4568 36864
rect 4890 36796 4896 36848
rect 4948 36836 4954 36848
rect 4948 36808 11744 36836
rect 4948 36796 4954 36808
rect 4019 36740 4568 36768
rect 4019 36737 4031 36740
rect 3973 36731 4031 36737
rect 6362 36728 6368 36780
rect 6420 36768 6426 36780
rect 6549 36771 6607 36777
rect 6549 36768 6561 36771
rect 6420 36740 6561 36768
rect 6420 36728 6426 36740
rect 6549 36737 6561 36740
rect 6595 36768 6607 36771
rect 7193 36771 7251 36777
rect 7193 36768 7205 36771
rect 6595 36740 7205 36768
rect 6595 36737 6607 36740
rect 6549 36731 6607 36737
rect 7193 36737 7205 36740
rect 7239 36737 7251 36771
rect 8386 36768 8392 36780
rect 8347 36740 8392 36768
rect 7193 36731 7251 36737
rect 8386 36728 8392 36740
rect 8444 36728 8450 36780
rect 9953 36771 10011 36777
rect 9953 36737 9965 36771
rect 9999 36768 10011 36771
rect 10502 36768 10508 36780
rect 9999 36740 10508 36768
rect 9999 36737 10011 36740
rect 9953 36731 10011 36737
rect 10502 36728 10508 36740
rect 10560 36728 10566 36780
rect 11716 36700 11744 36808
rect 13170 36796 13176 36848
rect 13228 36836 13234 36848
rect 21542 36836 21548 36848
rect 13228 36808 21548 36836
rect 13228 36796 13234 36808
rect 21542 36796 21548 36808
rect 21600 36796 21606 36848
rect 23934 36836 23940 36848
rect 21652 36808 23940 36836
rect 13814 36768 13820 36780
rect 13775 36740 13820 36768
rect 13814 36728 13820 36740
rect 13872 36768 13878 36780
rect 14461 36771 14519 36777
rect 14461 36768 14473 36771
rect 13872 36740 14473 36768
rect 13872 36728 13878 36740
rect 14461 36737 14473 36740
rect 14507 36737 14519 36771
rect 14461 36731 14519 36737
rect 17497 36771 17555 36777
rect 17497 36737 17509 36771
rect 17543 36768 17555 36771
rect 17954 36768 17960 36780
rect 17543 36740 17960 36768
rect 17543 36737 17555 36740
rect 17497 36731 17555 36737
rect 17954 36728 17960 36740
rect 18012 36728 18018 36780
rect 18046 36728 18052 36780
rect 18104 36768 18110 36780
rect 19150 36768 19156 36780
rect 18104 36740 19156 36768
rect 18104 36728 18110 36740
rect 19150 36728 19156 36740
rect 19208 36728 19214 36780
rect 19245 36771 19303 36777
rect 19245 36737 19257 36771
rect 19291 36768 19303 36771
rect 19889 36771 19947 36777
rect 19291 36740 19840 36768
rect 19291 36737 19303 36740
rect 19245 36731 19303 36737
rect 18509 36703 18567 36709
rect 11716 36672 18276 36700
rect 6733 36635 6791 36641
rect 6733 36601 6745 36635
rect 6779 36632 6791 36635
rect 12894 36632 12900 36644
rect 6779 36604 12900 36632
rect 6779 36601 6791 36604
rect 6733 36595 6791 36601
rect 12894 36592 12900 36604
rect 12952 36592 12958 36644
rect 14001 36635 14059 36641
rect 14001 36601 14013 36635
rect 14047 36632 14059 36635
rect 18046 36632 18052 36644
rect 14047 36604 18052 36632
rect 14047 36601 14059 36604
rect 14001 36595 14059 36601
rect 18046 36592 18052 36604
rect 18104 36592 18110 36644
rect 8386 36524 8392 36576
rect 8444 36564 8450 36576
rect 8941 36567 8999 36573
rect 8941 36564 8953 36567
rect 8444 36536 8953 36564
rect 8444 36524 8450 36536
rect 8941 36533 8953 36536
rect 8987 36564 8999 36567
rect 9582 36564 9588 36576
rect 8987 36536 9588 36564
rect 8987 36533 8999 36536
rect 8941 36527 8999 36533
rect 9582 36524 9588 36536
rect 9640 36524 9646 36576
rect 10502 36564 10508 36576
rect 10463 36536 10508 36564
rect 10502 36524 10508 36536
rect 10560 36524 10566 36576
rect 15930 36524 15936 36576
rect 15988 36564 15994 36576
rect 16117 36567 16175 36573
rect 16117 36564 16129 36567
rect 15988 36536 16129 36564
rect 15988 36524 15994 36536
rect 16117 36533 16129 36536
rect 16163 36564 16175 36567
rect 17678 36564 17684 36576
rect 16163 36536 17684 36564
rect 16163 36533 16175 36536
rect 16117 36527 16175 36533
rect 17678 36524 17684 36536
rect 17736 36524 17742 36576
rect 17954 36564 17960 36576
rect 17915 36536 17960 36564
rect 17954 36524 17960 36536
rect 18012 36524 18018 36576
rect 18248 36564 18276 36672
rect 18509 36669 18521 36703
rect 18555 36700 18567 36703
rect 19260 36700 19288 36731
rect 18555 36672 19288 36700
rect 18555 36669 18567 36672
rect 18509 36663 18567 36669
rect 19518 36660 19524 36712
rect 19576 36700 19582 36712
rect 19576 36672 19748 36700
rect 19576 36660 19582 36672
rect 19720 36641 19748 36672
rect 19705 36635 19763 36641
rect 19705 36601 19717 36635
rect 19751 36601 19763 36635
rect 19812 36632 19840 36740
rect 19889 36737 19901 36771
rect 19935 36768 19947 36771
rect 20714 36768 20720 36780
rect 19935 36740 20720 36768
rect 19935 36737 19947 36740
rect 19889 36731 19947 36737
rect 20714 36728 20720 36740
rect 20772 36728 20778 36780
rect 20809 36771 20867 36777
rect 20809 36737 20821 36771
rect 20855 36737 20867 36771
rect 20809 36731 20867 36737
rect 20162 36660 20168 36712
rect 20220 36700 20226 36712
rect 20824 36700 20852 36731
rect 21266 36728 21272 36780
rect 21324 36768 21330 36780
rect 21453 36771 21511 36777
rect 21453 36768 21465 36771
rect 21324 36740 21465 36768
rect 21324 36728 21330 36740
rect 21453 36737 21465 36740
rect 21499 36737 21511 36771
rect 21453 36731 21511 36737
rect 21652 36700 21680 36808
rect 23934 36796 23940 36808
rect 23992 36796 23998 36848
rect 24486 36836 24492 36848
rect 24447 36808 24492 36836
rect 24486 36796 24492 36808
rect 24544 36796 24550 36848
rect 24670 36796 24676 36848
rect 24728 36836 24734 36848
rect 24728 36808 25820 36836
rect 24728 36796 24734 36808
rect 21818 36728 21824 36780
rect 21876 36768 21882 36780
rect 22005 36771 22063 36777
rect 22005 36768 22017 36771
rect 21876 36740 22017 36768
rect 21876 36728 21882 36740
rect 22005 36737 22017 36740
rect 22051 36737 22063 36771
rect 22738 36768 22744 36780
rect 22699 36740 22744 36768
rect 22005 36731 22063 36737
rect 22738 36728 22744 36740
rect 22796 36728 22802 36780
rect 23293 36771 23351 36777
rect 23293 36737 23305 36771
rect 23339 36768 23351 36771
rect 23474 36768 23480 36780
rect 23339 36740 23480 36768
rect 23339 36737 23351 36740
rect 23293 36731 23351 36737
rect 23474 36728 23480 36740
rect 23532 36768 23538 36780
rect 23842 36768 23848 36780
rect 23532 36740 23848 36768
rect 23532 36728 23538 36740
rect 23842 36728 23848 36740
rect 23900 36728 23906 36780
rect 24118 36728 24124 36780
rect 24176 36768 24182 36780
rect 25314 36768 25320 36780
rect 24176 36740 25176 36768
rect 25275 36740 25320 36768
rect 24176 36728 24182 36740
rect 20220 36672 21680 36700
rect 20220 36660 20226 36672
rect 21726 36660 21732 36712
rect 21784 36700 21790 36712
rect 24397 36703 24455 36709
rect 24397 36700 24409 36703
rect 21784 36672 24409 36700
rect 21784 36660 21790 36672
rect 24397 36669 24409 36672
rect 24443 36669 24455 36703
rect 24397 36663 24455 36669
rect 24581 36703 24639 36709
rect 24581 36669 24593 36703
rect 24627 36700 24639 36703
rect 25038 36700 25044 36712
rect 24627 36672 25044 36700
rect 24627 36669 24639 36672
rect 24581 36663 24639 36669
rect 25038 36660 25044 36672
rect 25096 36660 25102 36712
rect 25148 36700 25176 36740
rect 25314 36728 25320 36740
rect 25372 36728 25378 36780
rect 25792 36777 25820 36808
rect 25866 36796 25872 36848
rect 25924 36836 25930 36848
rect 27246 36836 27252 36848
rect 25924 36808 27252 36836
rect 25924 36796 25930 36808
rect 27246 36796 27252 36808
rect 27304 36796 27310 36848
rect 27338 36796 27344 36848
rect 27396 36836 27402 36848
rect 29012 36836 29040 36876
rect 29641 36873 29653 36876
rect 29687 36904 29699 36907
rect 29822 36904 29828 36916
rect 29687 36876 29828 36904
rect 29687 36873 29699 36876
rect 29641 36867 29699 36873
rect 29822 36864 29828 36876
rect 29880 36864 29886 36916
rect 30374 36864 30380 36916
rect 30432 36904 30438 36916
rect 30469 36907 30527 36913
rect 30469 36904 30481 36907
rect 30432 36876 30481 36904
rect 30432 36864 30438 36876
rect 30469 36873 30481 36876
rect 30515 36873 30527 36907
rect 30469 36867 30527 36873
rect 30558 36864 30564 36916
rect 30616 36904 30622 36916
rect 32309 36907 32367 36913
rect 32309 36904 32321 36907
rect 30616 36876 32321 36904
rect 30616 36864 30622 36876
rect 32309 36873 32321 36876
rect 32355 36873 32367 36907
rect 32309 36867 32367 36873
rect 33134 36864 33140 36916
rect 33192 36904 33198 36916
rect 33229 36907 33287 36913
rect 33229 36904 33241 36907
rect 33192 36876 33241 36904
rect 33192 36864 33198 36876
rect 33229 36873 33241 36876
rect 33275 36873 33287 36907
rect 33229 36867 33287 36873
rect 34241 36907 34299 36913
rect 34241 36873 34253 36907
rect 34287 36904 34299 36907
rect 36446 36904 36452 36916
rect 34287 36876 36452 36904
rect 34287 36873 34299 36876
rect 34241 36867 34299 36873
rect 36446 36864 36452 36876
rect 36504 36864 36510 36916
rect 36722 36904 36728 36916
rect 36683 36876 36728 36904
rect 36722 36864 36728 36876
rect 36780 36864 36786 36916
rect 36814 36864 36820 36916
rect 36872 36904 36878 36916
rect 36872 36876 41414 36904
rect 36872 36864 36878 36876
rect 27396 36808 29040 36836
rect 29288 36808 33916 36836
rect 27396 36796 27402 36808
rect 25777 36771 25835 36777
rect 25777 36737 25789 36771
rect 25823 36737 25835 36771
rect 27985 36771 28043 36777
rect 27985 36768 27997 36771
rect 25777 36731 25835 36737
rect 25884 36740 27997 36768
rect 25884 36700 25912 36740
rect 27985 36737 27997 36740
rect 28031 36737 28043 36771
rect 27985 36731 28043 36737
rect 28626 36728 28632 36780
rect 28684 36768 28690 36780
rect 28810 36768 28816 36780
rect 28684 36740 28816 36768
rect 28684 36728 28690 36740
rect 28810 36728 28816 36740
rect 28868 36728 28874 36780
rect 29086 36728 29092 36780
rect 29144 36768 29150 36780
rect 29144 36740 29189 36768
rect 29144 36728 29150 36740
rect 25148 36672 25912 36700
rect 25958 36660 25964 36712
rect 26016 36700 26022 36712
rect 27801 36703 27859 36709
rect 27801 36700 27813 36703
rect 26016 36672 27813 36700
rect 26016 36660 26022 36672
rect 27801 36669 27813 36672
rect 27847 36669 27859 36703
rect 27801 36663 27859 36669
rect 27893 36703 27951 36709
rect 27893 36669 27905 36703
rect 27939 36700 27951 36703
rect 28534 36700 28540 36712
rect 27939 36672 28540 36700
rect 27939 36669 27951 36672
rect 27893 36663 27951 36669
rect 27154 36632 27160 36644
rect 19812 36604 27160 36632
rect 19705 36595 19763 36601
rect 27154 36592 27160 36604
rect 27212 36592 27218 36644
rect 27246 36592 27252 36644
rect 27304 36632 27310 36644
rect 27816 36632 27844 36663
rect 28534 36660 28540 36672
rect 28592 36700 28598 36712
rect 29288 36700 29316 36808
rect 30650 36768 30656 36780
rect 30611 36740 30656 36768
rect 30650 36728 30656 36740
rect 30708 36728 30714 36780
rect 31110 36768 31116 36780
rect 31071 36740 31116 36768
rect 31110 36728 31116 36740
rect 31168 36768 31174 36780
rect 31478 36768 31484 36780
rect 31168 36740 31484 36768
rect 31168 36728 31174 36740
rect 31478 36728 31484 36740
rect 31536 36728 31542 36780
rect 31757 36771 31815 36777
rect 31757 36737 31769 36771
rect 31803 36768 31815 36771
rect 32493 36771 32551 36777
rect 32493 36768 32505 36771
rect 31803 36740 32505 36768
rect 31803 36737 31815 36740
rect 31757 36731 31815 36737
rect 32493 36737 32505 36740
rect 32539 36768 32551 36771
rect 33042 36768 33048 36780
rect 32539 36740 33048 36768
rect 32539 36737 32551 36740
rect 32493 36731 32551 36737
rect 33042 36728 33048 36740
rect 33100 36728 33106 36780
rect 33134 36728 33140 36780
rect 33192 36768 33198 36780
rect 33410 36768 33416 36780
rect 33192 36740 33416 36768
rect 33192 36728 33198 36740
rect 33410 36728 33416 36740
rect 33468 36728 33474 36780
rect 33888 36700 33916 36808
rect 37274 36796 37280 36848
rect 37332 36836 37338 36848
rect 37719 36839 37777 36845
rect 37719 36836 37731 36839
rect 37332 36808 37731 36836
rect 37332 36796 37338 36808
rect 37719 36805 37731 36808
rect 37765 36805 37777 36839
rect 37719 36799 37777 36805
rect 38102 36796 38108 36848
rect 38160 36836 38166 36848
rect 38657 36839 38715 36845
rect 38657 36836 38669 36839
rect 38160 36808 38669 36836
rect 38160 36796 38166 36808
rect 38657 36805 38669 36808
rect 38703 36805 38715 36839
rect 40126 36836 40132 36848
rect 38657 36799 38715 36805
rect 38764 36808 40132 36836
rect 33962 36728 33968 36780
rect 34020 36768 34026 36780
rect 34057 36771 34115 36777
rect 34057 36768 34069 36771
rect 34020 36740 34069 36768
rect 34020 36728 34026 36740
rect 34057 36737 34069 36740
rect 34103 36737 34115 36771
rect 34057 36731 34115 36737
rect 34238 36728 34244 36780
rect 34296 36768 34302 36780
rect 35253 36771 35311 36777
rect 35253 36768 35265 36771
rect 34296 36740 35265 36768
rect 34296 36728 34302 36740
rect 35253 36737 35265 36740
rect 35299 36737 35311 36771
rect 35986 36768 35992 36780
rect 35947 36740 35992 36768
rect 35253 36731 35311 36737
rect 35986 36728 35992 36740
rect 36044 36728 36050 36780
rect 36906 36777 36912 36780
rect 36902 36731 36912 36777
rect 36964 36768 36970 36780
rect 36964 36740 37002 36768
rect 36906 36728 36912 36731
rect 36964 36728 36970 36740
rect 37090 36728 37096 36780
rect 37148 36768 37154 36780
rect 38764 36768 38792 36808
rect 40126 36796 40132 36808
rect 40184 36796 40190 36848
rect 41141 36839 41199 36845
rect 41141 36836 41153 36839
rect 40236 36808 41153 36836
rect 40236 36780 40264 36808
rect 41141 36805 41153 36808
rect 41187 36805 41199 36839
rect 41386 36836 41414 36876
rect 41598 36864 41604 36916
rect 41656 36904 41662 36916
rect 42613 36907 42671 36913
rect 42613 36904 42625 36907
rect 41656 36876 42625 36904
rect 41656 36864 41662 36876
rect 42613 36873 42625 36876
rect 42659 36873 42671 36907
rect 42613 36867 42671 36873
rect 42702 36864 42708 36916
rect 42760 36904 42766 36916
rect 42981 36907 43039 36913
rect 42981 36904 42993 36907
rect 42760 36876 42993 36904
rect 42760 36864 42766 36876
rect 42981 36873 42993 36876
rect 43027 36873 43039 36907
rect 42981 36867 43039 36873
rect 43901 36907 43959 36913
rect 43901 36873 43913 36907
rect 43947 36904 43959 36907
rect 44082 36904 44088 36916
rect 43947 36876 44088 36904
rect 43947 36873 43959 36876
rect 43901 36867 43959 36873
rect 44082 36864 44088 36876
rect 44140 36864 44146 36916
rect 44174 36864 44180 36916
rect 44232 36904 44238 36916
rect 53006 36904 53012 36916
rect 44232 36876 53012 36904
rect 44232 36864 44238 36876
rect 53006 36864 53012 36876
rect 53064 36864 53070 36916
rect 53098 36864 53104 36916
rect 53156 36904 53162 36916
rect 58437 36907 58495 36913
rect 58437 36904 58449 36907
rect 53156 36876 58449 36904
rect 53156 36864 53162 36876
rect 58437 36873 58449 36876
rect 58483 36873 58495 36907
rect 58437 36867 58495 36873
rect 60277 36907 60335 36913
rect 60277 36873 60289 36907
rect 60323 36904 60335 36907
rect 60642 36904 60648 36916
rect 60323 36876 60648 36904
rect 60323 36873 60335 36876
rect 60277 36867 60335 36873
rect 60642 36864 60648 36876
rect 60700 36864 60706 36916
rect 62669 36907 62727 36913
rect 62669 36873 62681 36907
rect 62715 36904 62727 36907
rect 64782 36904 64788 36916
rect 62715 36876 64788 36904
rect 62715 36873 62727 36876
rect 62669 36867 62727 36873
rect 64782 36864 64788 36876
rect 64840 36864 64846 36916
rect 65429 36907 65487 36913
rect 65429 36904 65441 36907
rect 65168 36876 65441 36904
rect 64874 36836 64880 36848
rect 41386 36808 64880 36836
rect 41141 36799 41199 36805
rect 64874 36796 64880 36808
rect 64932 36796 64938 36848
rect 37148 36740 38792 36768
rect 37148 36728 37154 36740
rect 38838 36728 38844 36780
rect 38896 36768 38902 36780
rect 39853 36771 39911 36777
rect 38896 36740 38941 36768
rect 38896 36728 38902 36740
rect 39853 36737 39865 36771
rect 39899 36768 39911 36771
rect 40218 36768 40224 36780
rect 39899 36740 40224 36768
rect 39899 36737 39911 36740
rect 39853 36731 39911 36737
rect 40218 36728 40224 36740
rect 40276 36728 40282 36780
rect 40589 36771 40647 36777
rect 40589 36737 40601 36771
rect 40635 36768 40647 36771
rect 40954 36768 40960 36780
rect 40635 36740 40960 36768
rect 40635 36737 40647 36740
rect 40589 36731 40647 36737
rect 40954 36728 40960 36740
rect 41012 36768 41018 36780
rect 41877 36771 41935 36777
rect 41877 36768 41889 36771
rect 41012 36740 41889 36768
rect 41012 36728 41018 36740
rect 41877 36737 41889 36740
rect 41923 36737 41935 36771
rect 41877 36731 41935 36737
rect 42794 36728 42800 36780
rect 42852 36768 42858 36780
rect 42852 36740 43208 36768
rect 42852 36728 42858 36740
rect 43070 36700 43076 36712
rect 28592 36672 29316 36700
rect 29380 36672 33456 36700
rect 33888 36672 42932 36700
rect 43031 36672 43076 36700
rect 28592 36660 28598 36672
rect 27982 36632 27988 36644
rect 27304 36604 27752 36632
rect 27816 36604 27988 36632
rect 27304 36592 27310 36604
rect 20254 36564 20260 36576
rect 18248 36536 20260 36564
rect 20254 36524 20260 36536
rect 20312 36524 20318 36576
rect 20806 36524 20812 36576
rect 20864 36564 20870 36576
rect 21269 36567 21327 36573
rect 21269 36564 21281 36567
rect 20864 36536 21281 36564
rect 20864 36524 20870 36536
rect 21269 36533 21281 36536
rect 21315 36533 21327 36567
rect 22186 36564 22192 36576
rect 22147 36536 22192 36564
rect 21269 36527 21327 36533
rect 22186 36524 22192 36536
rect 22244 36524 22250 36576
rect 23477 36567 23535 36573
rect 23477 36533 23489 36567
rect 23523 36564 23535 36567
rect 23934 36564 23940 36576
rect 23523 36536 23940 36564
rect 23523 36533 23535 36536
rect 23477 36527 23535 36533
rect 23934 36524 23940 36536
rect 23992 36524 23998 36576
rect 24029 36567 24087 36573
rect 24029 36533 24041 36567
rect 24075 36564 24087 36567
rect 24670 36564 24676 36576
rect 24075 36536 24676 36564
rect 24075 36533 24087 36536
rect 24029 36527 24087 36533
rect 24670 36524 24676 36536
rect 24728 36524 24734 36576
rect 24854 36524 24860 36576
rect 24912 36564 24918 36576
rect 25133 36567 25191 36573
rect 25133 36564 25145 36567
rect 24912 36536 25145 36564
rect 24912 36524 24918 36536
rect 25133 36533 25145 36536
rect 25179 36533 25191 36567
rect 25958 36564 25964 36576
rect 25919 36536 25964 36564
rect 25133 36527 25191 36533
rect 25958 36524 25964 36536
rect 26016 36524 26022 36576
rect 26605 36567 26663 36573
rect 26605 36533 26617 36567
rect 26651 36564 26663 36567
rect 26694 36564 26700 36576
rect 26651 36536 26700 36564
rect 26651 36533 26663 36536
rect 26605 36527 26663 36533
rect 26694 36524 26700 36536
rect 26752 36564 26758 36576
rect 27338 36564 27344 36576
rect 26752 36536 27344 36564
rect 26752 36524 26758 36536
rect 27338 36524 27344 36536
rect 27396 36524 27402 36576
rect 27724 36564 27752 36604
rect 27982 36592 27988 36604
rect 28040 36632 28046 36644
rect 28626 36632 28632 36644
rect 28040 36604 28632 36632
rect 28040 36592 28046 36604
rect 28626 36592 28632 36604
rect 28684 36592 28690 36644
rect 28902 36592 28908 36644
rect 28960 36632 28966 36644
rect 29380 36632 29408 36672
rect 28960 36604 29408 36632
rect 28960 36592 28966 36604
rect 29638 36592 29644 36644
rect 29696 36632 29702 36644
rect 33428 36632 33456 36672
rect 33594 36632 33600 36644
rect 29696 36604 33364 36632
rect 33428 36604 33600 36632
rect 29696 36592 29702 36604
rect 33226 36564 33232 36576
rect 27724 36536 33232 36564
rect 33226 36524 33232 36536
rect 33284 36524 33290 36576
rect 33336 36564 33364 36604
rect 33594 36592 33600 36604
rect 33652 36592 33658 36644
rect 35618 36632 35624 36644
rect 33704 36604 35624 36632
rect 33704 36564 33732 36604
rect 35618 36592 35624 36604
rect 35676 36592 35682 36644
rect 35710 36592 35716 36644
rect 35768 36632 35774 36644
rect 39669 36635 39727 36641
rect 39669 36632 39681 36635
rect 35768 36604 39681 36632
rect 35768 36592 35774 36604
rect 39669 36601 39681 36604
rect 39715 36601 39727 36635
rect 39669 36595 39727 36601
rect 40310 36592 40316 36644
rect 40368 36632 40374 36644
rect 40405 36635 40463 36641
rect 40405 36632 40417 36635
rect 40368 36604 40417 36632
rect 40368 36592 40374 36604
rect 40405 36601 40417 36604
rect 40451 36601 40463 36635
rect 41046 36632 41052 36644
rect 40405 36595 40463 36601
rect 40880 36604 41052 36632
rect 33336 36536 33732 36564
rect 33778 36524 33784 36576
rect 33836 36564 33842 36576
rect 34606 36564 34612 36576
rect 33836 36536 34612 36564
rect 33836 36524 33842 36536
rect 34606 36524 34612 36536
rect 34664 36524 34670 36576
rect 35342 36564 35348 36576
rect 35303 36536 35348 36564
rect 35342 36524 35348 36536
rect 35400 36524 35406 36576
rect 36081 36567 36139 36573
rect 36081 36533 36093 36567
rect 36127 36564 36139 36567
rect 37182 36564 37188 36576
rect 36127 36536 37188 36564
rect 36127 36533 36139 36536
rect 36081 36527 36139 36533
rect 37182 36524 37188 36536
rect 37240 36524 37246 36576
rect 37550 36524 37556 36576
rect 37608 36564 37614 36576
rect 37829 36567 37887 36573
rect 37829 36564 37841 36567
rect 37608 36536 37841 36564
rect 37608 36524 37614 36536
rect 37829 36533 37841 36536
rect 37875 36533 37887 36567
rect 37829 36527 37887 36533
rect 39298 36524 39304 36576
rect 39356 36564 39362 36576
rect 40880 36564 40908 36604
rect 41046 36592 41052 36604
rect 41104 36592 41110 36644
rect 41322 36632 41328 36644
rect 41283 36604 41328 36632
rect 41322 36592 41328 36604
rect 41380 36592 41386 36644
rect 42904 36632 42932 36672
rect 43070 36660 43076 36672
rect 43128 36660 43134 36712
rect 43180 36709 43208 36740
rect 43990 36728 43996 36780
rect 44048 36768 44054 36780
rect 44085 36771 44143 36777
rect 44085 36768 44097 36771
rect 44048 36740 44097 36768
rect 44048 36728 44054 36740
rect 44085 36737 44097 36740
rect 44131 36737 44143 36771
rect 44634 36768 44640 36780
rect 44595 36740 44640 36768
rect 44085 36731 44143 36737
rect 44634 36728 44640 36740
rect 44692 36728 44698 36780
rect 45002 36728 45008 36780
rect 45060 36768 45066 36780
rect 45281 36771 45339 36777
rect 45281 36768 45293 36771
rect 45060 36740 45293 36768
rect 45060 36728 45066 36740
rect 45281 36737 45293 36740
rect 45327 36737 45339 36771
rect 46290 36768 46296 36780
rect 46251 36740 46296 36768
rect 45281 36731 45339 36737
rect 46290 36728 46296 36740
rect 46348 36728 46354 36780
rect 47210 36768 47216 36780
rect 47171 36740 47216 36768
rect 47210 36728 47216 36740
rect 47268 36728 47274 36780
rect 47302 36728 47308 36780
rect 47360 36768 47366 36780
rect 48133 36771 48191 36777
rect 48133 36768 48145 36771
rect 47360 36740 48145 36768
rect 47360 36728 47366 36740
rect 48133 36737 48145 36740
rect 48179 36737 48191 36771
rect 48133 36731 48191 36737
rect 48590 36728 48596 36780
rect 48648 36768 48654 36780
rect 49053 36771 49111 36777
rect 49053 36768 49065 36771
rect 48648 36740 49065 36768
rect 48648 36728 48654 36740
rect 49053 36737 49065 36740
rect 49099 36737 49111 36771
rect 50246 36768 50252 36780
rect 50207 36740 50252 36768
rect 49053 36731 49111 36737
rect 50246 36728 50252 36740
rect 50304 36728 50310 36780
rect 50433 36771 50491 36777
rect 50433 36737 50445 36771
rect 50479 36768 50491 36771
rect 50890 36768 50896 36780
rect 50479 36740 50896 36768
rect 50479 36737 50491 36740
rect 50433 36731 50491 36737
rect 50890 36728 50896 36740
rect 50948 36728 50954 36780
rect 51626 36768 51632 36780
rect 51587 36740 51632 36768
rect 51626 36728 51632 36740
rect 51684 36728 51690 36780
rect 52086 36768 52092 36780
rect 52047 36740 52092 36768
rect 52086 36728 52092 36740
rect 52144 36728 52150 36780
rect 52273 36771 52331 36777
rect 52273 36737 52285 36771
rect 52319 36737 52331 36771
rect 52273 36731 52331 36737
rect 43165 36703 43223 36709
rect 43165 36669 43177 36703
rect 43211 36669 43223 36703
rect 43165 36663 43223 36669
rect 43456 36672 46244 36700
rect 43456 36632 43484 36672
rect 44818 36632 44824 36644
rect 42904 36604 43484 36632
rect 44779 36604 44824 36632
rect 44818 36592 44824 36604
rect 44876 36592 44882 36644
rect 45830 36632 45836 36644
rect 44928 36604 45836 36632
rect 41966 36564 41972 36576
rect 39356 36536 40908 36564
rect 41927 36536 41972 36564
rect 39356 36524 39362 36536
rect 41966 36524 41972 36536
rect 42024 36524 42030 36576
rect 42058 36524 42064 36576
rect 42116 36564 42122 36576
rect 44928 36564 44956 36604
rect 45830 36592 45836 36604
rect 45888 36592 45894 36644
rect 45922 36592 45928 36644
rect 45980 36632 45986 36644
rect 46109 36635 46167 36641
rect 46109 36632 46121 36635
rect 45980 36604 46121 36632
rect 45980 36592 45986 36604
rect 46109 36601 46121 36604
rect 46155 36601 46167 36635
rect 46216 36632 46244 36672
rect 47854 36660 47860 36712
rect 47912 36700 47918 36712
rect 48038 36700 48044 36712
rect 47912 36672 47957 36700
rect 47999 36672 48044 36700
rect 47912 36660 47918 36672
rect 48038 36660 48044 36672
rect 48096 36660 48102 36712
rect 51810 36700 51816 36712
rect 48286 36672 51816 36700
rect 48286 36632 48314 36672
rect 51810 36660 51816 36672
rect 51868 36660 51874 36712
rect 52288 36700 52316 36731
rect 53006 36728 53012 36780
rect 53064 36768 53070 36780
rect 53561 36771 53619 36777
rect 53561 36768 53573 36771
rect 53064 36740 53573 36768
rect 53064 36728 53070 36740
rect 53561 36737 53573 36740
rect 53607 36737 53619 36771
rect 53561 36731 53619 36737
rect 53926 36728 53932 36780
rect 53984 36768 53990 36780
rect 54297 36771 54355 36777
rect 54297 36768 54309 36771
rect 53984 36740 54309 36768
rect 53984 36728 53990 36740
rect 54297 36737 54309 36740
rect 54343 36737 54355 36771
rect 54297 36731 54355 36737
rect 54941 36771 54999 36777
rect 54941 36737 54953 36771
rect 54987 36737 54999 36771
rect 55582 36768 55588 36780
rect 55543 36740 55588 36768
rect 54941 36731 54999 36737
rect 53944 36700 53972 36728
rect 52012 36672 53972 36700
rect 46216 36604 48314 36632
rect 48501 36635 48559 36641
rect 46109 36595 46167 36601
rect 48501 36601 48513 36635
rect 48547 36632 48559 36635
rect 49510 36632 49516 36644
rect 48547 36604 49516 36632
rect 48547 36601 48559 36604
rect 48501 36595 48559 36601
rect 49510 36592 49516 36604
rect 49568 36592 49574 36644
rect 50985 36635 51043 36641
rect 50985 36601 50997 36635
rect 51031 36632 51043 36635
rect 52012 36632 52040 36672
rect 54202 36660 54208 36712
rect 54260 36700 54266 36712
rect 54754 36700 54760 36712
rect 54260 36672 54760 36700
rect 54260 36660 54266 36672
rect 54754 36660 54760 36672
rect 54812 36700 54818 36712
rect 54956 36700 54984 36731
rect 55582 36728 55588 36740
rect 55640 36728 55646 36780
rect 55769 36771 55827 36777
rect 55769 36737 55781 36771
rect 55815 36737 55827 36771
rect 55769 36731 55827 36737
rect 54812 36672 54984 36700
rect 55784 36700 55812 36731
rect 56042 36728 56048 36780
rect 56100 36768 56106 36780
rect 56321 36771 56379 36777
rect 56321 36768 56333 36771
rect 56100 36740 56333 36768
rect 56100 36728 56106 36740
rect 56321 36737 56333 36740
rect 56367 36737 56379 36771
rect 56321 36731 56379 36737
rect 57149 36771 57207 36777
rect 57149 36737 57161 36771
rect 57195 36768 57207 36771
rect 57330 36768 57336 36780
rect 57195 36740 57336 36768
rect 57195 36737 57207 36740
rect 57149 36731 57207 36737
rect 57330 36728 57336 36740
rect 57388 36728 57394 36780
rect 57422 36728 57428 36780
rect 57480 36768 57486 36780
rect 59357 36771 59415 36777
rect 59357 36768 59369 36771
rect 57480 36740 59369 36768
rect 57480 36728 57486 36740
rect 59357 36737 59369 36740
rect 59403 36737 59415 36771
rect 59357 36731 59415 36737
rect 59541 36771 59599 36777
rect 59541 36737 59553 36771
rect 59587 36737 59599 36771
rect 60090 36768 60096 36780
rect 60051 36740 60096 36768
rect 59541 36731 59599 36737
rect 56594 36700 56600 36712
rect 55784 36672 56600 36700
rect 54812 36660 54818 36672
rect 56594 36660 56600 36672
rect 56652 36660 56658 36712
rect 58250 36700 58256 36712
rect 58211 36672 58256 36700
rect 58250 36660 58256 36672
rect 58308 36660 58314 36712
rect 58345 36703 58403 36709
rect 58345 36669 58357 36703
rect 58391 36700 58403 36703
rect 58526 36700 58532 36712
rect 58391 36672 58532 36700
rect 58391 36669 58403 36672
rect 58345 36663 58403 36669
rect 58526 36660 58532 36672
rect 58584 36660 58590 36712
rect 59556 36700 59584 36731
rect 60090 36728 60096 36740
rect 60148 36728 60154 36780
rect 60734 36768 60740 36780
rect 60568 36740 60740 36768
rect 60568 36700 60596 36740
rect 60734 36728 60740 36740
rect 60792 36768 60798 36780
rect 60921 36771 60979 36777
rect 60921 36768 60933 36771
rect 60792 36740 60933 36768
rect 60792 36728 60798 36740
rect 60921 36737 60933 36740
rect 60967 36737 60979 36771
rect 61654 36768 61660 36780
rect 61615 36740 61660 36768
rect 60921 36731 60979 36737
rect 61654 36728 61660 36740
rect 61712 36728 61718 36780
rect 62114 36728 62120 36780
rect 62172 36768 62178 36780
rect 62485 36771 62543 36777
rect 62485 36768 62497 36771
rect 62172 36740 62497 36768
rect 62172 36728 62178 36740
rect 62485 36737 62497 36740
rect 62531 36737 62543 36771
rect 62485 36731 62543 36737
rect 63221 36771 63279 36777
rect 63221 36737 63233 36771
rect 63267 36768 63279 36771
rect 63402 36768 63408 36780
rect 63267 36740 63408 36768
rect 63267 36737 63279 36740
rect 63221 36731 63279 36737
rect 63402 36728 63408 36740
rect 63460 36728 63466 36780
rect 64230 36768 64236 36780
rect 64191 36740 64236 36768
rect 64230 36728 64236 36740
rect 64288 36728 64294 36780
rect 64325 36771 64383 36777
rect 64325 36737 64337 36771
rect 64371 36768 64383 36771
rect 64414 36768 64420 36780
rect 64371 36740 64420 36768
rect 64371 36737 64383 36740
rect 64325 36731 64383 36737
rect 64414 36728 64420 36740
rect 64472 36728 64478 36780
rect 64598 36728 64604 36780
rect 64656 36768 64662 36780
rect 65168 36768 65196 36876
rect 65429 36873 65441 36876
rect 65475 36873 65487 36907
rect 65429 36867 65487 36873
rect 66254 36864 66260 36916
rect 66312 36904 66318 36916
rect 66349 36907 66407 36913
rect 66349 36904 66361 36907
rect 66312 36876 66361 36904
rect 66312 36864 66318 36876
rect 66349 36873 66361 36876
rect 66395 36873 66407 36907
rect 66349 36867 66407 36873
rect 67361 36907 67419 36913
rect 67361 36873 67373 36907
rect 67407 36904 67419 36907
rect 72786 36904 72792 36916
rect 67407 36876 72792 36904
rect 67407 36873 67419 36876
rect 67361 36867 67419 36873
rect 72786 36864 72792 36876
rect 72844 36864 72850 36916
rect 72881 36907 72939 36913
rect 72881 36873 72893 36907
rect 72927 36904 72939 36907
rect 74718 36904 74724 36916
rect 72927 36876 74724 36904
rect 72927 36873 72939 36876
rect 72881 36867 72939 36873
rect 74718 36864 74724 36876
rect 74776 36864 74782 36916
rect 76282 36864 76288 36916
rect 76340 36904 76346 36916
rect 76561 36907 76619 36913
rect 76561 36904 76573 36907
rect 76340 36876 76573 36904
rect 76340 36864 76346 36876
rect 76561 36873 76573 36876
rect 76607 36873 76619 36907
rect 76561 36867 76619 36873
rect 77018 36864 77024 36916
rect 77076 36904 77082 36916
rect 77113 36907 77171 36913
rect 77113 36904 77125 36907
rect 77076 36876 77125 36904
rect 77076 36864 77082 36876
rect 77113 36873 77125 36876
rect 77159 36873 77171 36907
rect 77113 36867 77171 36873
rect 78674 36864 78680 36916
rect 78732 36904 78738 36916
rect 78769 36907 78827 36913
rect 78769 36904 78781 36907
rect 78732 36876 78781 36904
rect 78732 36864 78738 36876
rect 78769 36873 78781 36876
rect 78815 36873 78827 36907
rect 78769 36867 78827 36873
rect 80149 36907 80207 36913
rect 80149 36873 80161 36907
rect 80195 36904 80207 36907
rect 80238 36904 80244 36916
rect 80195 36876 80244 36904
rect 80195 36873 80207 36876
rect 80149 36867 80207 36873
rect 80238 36864 80244 36876
rect 80296 36864 80302 36916
rect 80330 36864 80336 36916
rect 80388 36904 80394 36916
rect 119706 36904 119712 36916
rect 80388 36876 119712 36904
rect 80388 36864 80394 36876
rect 119706 36864 119712 36876
rect 119764 36864 119770 36916
rect 119890 36904 119896 36916
rect 119851 36876 119896 36904
rect 119890 36864 119896 36876
rect 119948 36864 119954 36916
rect 119982 36864 119988 36916
rect 120040 36904 120046 36916
rect 123570 36904 123576 36916
rect 120040 36876 123576 36904
rect 120040 36864 120046 36876
rect 123570 36864 123576 36876
rect 123628 36864 123634 36916
rect 124398 36904 124404 36916
rect 124359 36876 124404 36904
rect 124398 36864 124404 36876
rect 124456 36864 124462 36916
rect 124950 36864 124956 36916
rect 125008 36904 125014 36916
rect 125045 36907 125103 36913
rect 125045 36904 125057 36907
rect 125008 36876 125057 36904
rect 125008 36864 125014 36876
rect 125045 36873 125057 36876
rect 125091 36873 125103 36907
rect 125594 36904 125600 36916
rect 125555 36876 125600 36904
rect 125045 36867 125103 36873
rect 125594 36864 125600 36876
rect 125652 36864 125658 36916
rect 126514 36904 126520 36916
rect 126475 36876 126520 36904
rect 126514 36864 126520 36876
rect 126572 36864 126578 36916
rect 127710 36904 127716 36916
rect 127671 36876 127716 36904
rect 127710 36864 127716 36876
rect 127768 36864 127774 36916
rect 128354 36904 128360 36916
rect 128315 36876 128360 36904
rect 128354 36864 128360 36876
rect 128412 36864 128418 36916
rect 128722 36864 128728 36916
rect 128780 36904 128786 36916
rect 128909 36907 128967 36913
rect 128909 36904 128921 36907
rect 128780 36876 128921 36904
rect 128780 36864 128786 36876
rect 128909 36873 128921 36876
rect 128955 36873 128967 36907
rect 128909 36867 128967 36873
rect 131114 36864 131120 36916
rect 131172 36904 131178 36916
rect 131485 36907 131543 36913
rect 131485 36904 131497 36907
rect 131172 36876 131497 36904
rect 131172 36864 131178 36876
rect 131485 36873 131497 36876
rect 131531 36873 131543 36907
rect 131485 36867 131543 36873
rect 132221 36907 132279 36913
rect 132221 36873 132233 36907
rect 132267 36904 132279 36907
rect 133230 36904 133236 36916
rect 132267 36876 132494 36904
rect 133191 36876 133236 36904
rect 132267 36873 132279 36876
rect 132221 36867 132279 36873
rect 65334 36796 65340 36848
rect 65392 36836 65398 36848
rect 65392 36808 65437 36836
rect 65392 36796 65398 36808
rect 65518 36796 65524 36848
rect 65576 36836 65582 36848
rect 87230 36836 87236 36848
rect 65576 36808 87236 36836
rect 65576 36796 65582 36808
rect 87230 36796 87236 36808
rect 87288 36796 87294 36848
rect 87506 36836 87512 36848
rect 87467 36808 87512 36836
rect 87506 36796 87512 36808
rect 87564 36796 87570 36848
rect 87598 36796 87604 36848
rect 87656 36836 87662 36848
rect 87656 36808 96108 36836
rect 87656 36796 87662 36808
rect 66530 36768 66536 36780
rect 64656 36740 65196 36768
rect 66491 36740 66536 36768
rect 64656 36728 64662 36740
rect 66530 36728 66536 36740
rect 66588 36728 66594 36780
rect 67082 36728 67088 36780
rect 67140 36768 67146 36780
rect 67177 36771 67235 36777
rect 67177 36768 67189 36771
rect 67140 36740 67189 36768
rect 67140 36728 67146 36740
rect 67177 36737 67189 36740
rect 67223 36737 67235 36771
rect 68646 36768 68652 36780
rect 68607 36740 68652 36768
rect 67177 36731 67235 36737
rect 68646 36728 68652 36740
rect 68704 36728 68710 36780
rect 68833 36771 68891 36777
rect 68833 36737 68845 36771
rect 68879 36768 68891 36771
rect 69198 36768 69204 36780
rect 68879 36740 69204 36768
rect 68879 36737 68891 36740
rect 68833 36731 68891 36737
rect 69198 36728 69204 36740
rect 69256 36768 69262 36780
rect 69477 36771 69535 36777
rect 69477 36768 69489 36771
rect 69256 36740 69489 36768
rect 69256 36728 69262 36740
rect 69477 36737 69489 36740
rect 69523 36737 69535 36771
rect 69658 36768 69664 36780
rect 69619 36740 69664 36768
rect 69477 36731 69535 36737
rect 69658 36728 69664 36740
rect 69716 36728 69722 36780
rect 70397 36771 70455 36777
rect 70397 36737 70409 36771
rect 70443 36768 70455 36771
rect 70762 36768 70768 36780
rect 70443 36740 70768 36768
rect 70443 36737 70455 36740
rect 70397 36731 70455 36737
rect 70762 36728 70768 36740
rect 70820 36768 70826 36780
rect 70857 36771 70915 36777
rect 70857 36768 70869 36771
rect 70820 36740 70869 36768
rect 70820 36728 70826 36740
rect 70857 36737 70869 36740
rect 70903 36737 70915 36771
rect 70857 36731 70915 36737
rect 72237 36771 72295 36777
rect 72237 36737 72249 36771
rect 72283 36768 72295 36771
rect 72602 36768 72608 36780
rect 72283 36740 72608 36768
rect 72283 36737 72295 36740
rect 72237 36731 72295 36737
rect 72602 36728 72608 36740
rect 72660 36768 72666 36780
rect 72697 36771 72755 36777
rect 72697 36768 72709 36771
rect 72660 36740 72709 36768
rect 72660 36728 72666 36740
rect 72697 36737 72709 36740
rect 72743 36737 72755 36771
rect 72697 36731 72755 36737
rect 74534 36728 74540 36780
rect 74592 36768 74598 36780
rect 75178 36768 75184 36780
rect 74592 36740 75184 36768
rect 74592 36728 74598 36740
rect 75178 36728 75184 36740
rect 75236 36768 75242 36780
rect 75273 36771 75331 36777
rect 75273 36768 75285 36771
rect 75236 36740 75285 36768
rect 75236 36728 75242 36740
rect 75273 36737 75285 36740
rect 75319 36768 75331 36771
rect 76190 36768 76196 36780
rect 75319 36740 76196 36768
rect 75319 36737 75331 36740
rect 75273 36731 75331 36737
rect 76190 36728 76196 36740
rect 76248 36728 76254 36780
rect 76282 36728 76288 36780
rect 76340 36768 76346 36780
rect 76377 36771 76435 36777
rect 76377 36768 76389 36771
rect 76340 36740 76389 36768
rect 76340 36728 76346 36740
rect 76377 36737 76389 36740
rect 76423 36737 76435 36771
rect 78950 36768 78956 36780
rect 78911 36740 78956 36768
rect 76377 36731 76435 36737
rect 78950 36728 78956 36740
rect 79008 36728 79014 36780
rect 79134 36728 79140 36780
rect 79192 36768 79198 36780
rect 80057 36771 80115 36777
rect 79192 36766 80008 36768
rect 80057 36766 80069 36771
rect 79192 36740 80069 36766
rect 79192 36728 79198 36740
rect 79980 36738 80069 36740
rect 80057 36737 80069 36738
rect 80103 36737 80115 36771
rect 80514 36768 80520 36780
rect 80057 36731 80115 36737
rect 80256 36740 80520 36768
rect 59556 36672 60596 36700
rect 61933 36703 61991 36709
rect 61933 36669 61945 36703
rect 61979 36700 61991 36703
rect 62390 36700 62396 36712
rect 61979 36672 62396 36700
rect 61979 36669 61991 36672
rect 61933 36663 61991 36669
rect 62390 36660 62396 36672
rect 62448 36700 62454 36712
rect 63954 36700 63960 36712
rect 62448 36672 63960 36700
rect 62448 36660 62454 36672
rect 63954 36660 63960 36672
rect 64012 36660 64018 36712
rect 64509 36703 64567 36709
rect 64509 36669 64521 36703
rect 64555 36700 64567 36703
rect 65058 36700 65064 36712
rect 64555 36672 65064 36700
rect 64555 36669 64567 36672
rect 64509 36663 64567 36669
rect 65058 36660 65064 36672
rect 65116 36700 65122 36712
rect 65153 36703 65211 36709
rect 65153 36700 65165 36703
rect 65116 36672 65165 36700
rect 65116 36660 65122 36672
rect 65153 36669 65165 36672
rect 65199 36669 65211 36703
rect 65153 36663 65211 36669
rect 65536 36672 65748 36700
rect 53006 36632 53012 36644
rect 51031 36604 52040 36632
rect 52967 36604 53012 36632
rect 51031 36601 51043 36604
rect 50985 36595 51043 36601
rect 53006 36592 53012 36604
rect 53064 36592 53070 36644
rect 64966 36632 64972 36644
rect 53116 36604 64972 36632
rect 42116 36536 44956 36564
rect 45465 36567 45523 36573
rect 42116 36524 42122 36536
rect 45465 36533 45477 36567
rect 45511 36564 45523 36567
rect 46750 36564 46756 36576
rect 45511 36536 46756 36564
rect 45511 36533 45523 36536
rect 45465 36527 45523 36533
rect 46750 36524 46756 36536
rect 46808 36524 46814 36576
rect 47026 36564 47032 36576
rect 46987 36536 47032 36564
rect 47026 36524 47032 36536
rect 47084 36524 47090 36576
rect 47118 36524 47124 36576
rect 47176 36564 47182 36576
rect 47854 36564 47860 36576
rect 47176 36536 47860 36564
rect 47176 36524 47182 36536
rect 47854 36524 47860 36536
rect 47912 36524 47918 36576
rect 48038 36524 48044 36576
rect 48096 36564 48102 36576
rect 48222 36564 48228 36576
rect 48096 36536 48228 36564
rect 48096 36524 48102 36536
rect 48222 36524 48228 36536
rect 48280 36524 48286 36576
rect 49142 36564 49148 36576
rect 49103 36536 49148 36564
rect 49142 36524 49148 36536
rect 49200 36524 49206 36576
rect 51442 36564 51448 36576
rect 51403 36536 51448 36564
rect 51442 36524 51448 36536
rect 51500 36524 51506 36576
rect 51810 36524 51816 36576
rect 51868 36564 51874 36576
rect 53116 36564 53144 36604
rect 64966 36592 64972 36604
rect 65024 36592 65030 36644
rect 65536 36632 65564 36672
rect 65352 36604 65564 36632
rect 65720 36632 65748 36672
rect 65794 36660 65800 36712
rect 65852 36700 65858 36712
rect 75454 36700 75460 36712
rect 65852 36672 75460 36700
rect 65852 36660 65858 36672
rect 75454 36660 75460 36672
rect 75512 36660 75518 36712
rect 76650 36660 76656 36712
rect 76708 36700 76714 36712
rect 80256 36700 80284 36740
rect 80514 36728 80520 36740
rect 80572 36728 80578 36780
rect 80606 36728 80612 36780
rect 80664 36768 80670 36780
rect 81253 36771 81311 36777
rect 81253 36768 81265 36771
rect 80664 36740 81265 36768
rect 80664 36728 80670 36740
rect 81253 36737 81265 36740
rect 81299 36737 81311 36771
rect 82078 36768 82084 36780
rect 82039 36740 82084 36768
rect 81253 36731 81311 36737
rect 82078 36728 82084 36740
rect 82136 36728 82142 36780
rect 82262 36768 82268 36780
rect 82223 36740 82268 36768
rect 82262 36728 82268 36740
rect 82320 36728 82326 36780
rect 83093 36771 83151 36777
rect 83093 36737 83105 36771
rect 83139 36768 83151 36771
rect 83182 36768 83188 36780
rect 83139 36740 83188 36768
rect 83139 36737 83151 36740
rect 83093 36731 83151 36737
rect 83182 36728 83188 36740
rect 83240 36768 83246 36780
rect 83734 36768 83740 36780
rect 83240 36740 83740 36768
rect 83240 36728 83246 36740
rect 83734 36728 83740 36740
rect 83792 36728 83798 36780
rect 83826 36728 83832 36780
rect 83884 36768 83890 36780
rect 84930 36768 84936 36780
rect 83884 36740 83929 36768
rect 84891 36740 84936 36768
rect 83884 36728 83890 36740
rect 84930 36728 84936 36740
rect 84988 36728 84994 36780
rect 85117 36771 85175 36777
rect 85117 36737 85129 36771
rect 85163 36768 85175 36771
rect 85482 36768 85488 36780
rect 85163 36740 85488 36768
rect 85163 36737 85175 36740
rect 85117 36731 85175 36737
rect 85482 36728 85488 36740
rect 85540 36768 85546 36780
rect 86313 36771 86371 36777
rect 86313 36768 86325 36771
rect 85540 36740 86325 36768
rect 85540 36728 85546 36740
rect 86313 36737 86325 36740
rect 86359 36737 86371 36771
rect 86313 36731 86371 36737
rect 89070 36728 89076 36780
rect 89128 36768 89134 36780
rect 89257 36771 89315 36777
rect 89257 36768 89269 36771
rect 89128 36740 89269 36768
rect 89128 36728 89134 36740
rect 89257 36737 89269 36740
rect 89303 36737 89315 36771
rect 90358 36768 90364 36780
rect 90319 36740 90364 36768
rect 89257 36731 89315 36737
rect 90358 36728 90364 36740
rect 90416 36768 90422 36780
rect 91005 36771 91063 36777
rect 91005 36768 91017 36771
rect 90416 36740 91017 36768
rect 90416 36728 90422 36740
rect 91005 36737 91017 36740
rect 91051 36737 91063 36771
rect 93026 36768 93032 36780
rect 92987 36740 93032 36768
rect 91005 36731 91063 36737
rect 93026 36728 93032 36740
rect 93084 36728 93090 36780
rect 93213 36771 93271 36777
rect 93213 36737 93225 36771
rect 93259 36768 93271 36771
rect 94314 36768 94320 36780
rect 93259 36740 94320 36768
rect 93259 36737 93271 36740
rect 93213 36731 93271 36737
rect 94314 36728 94320 36740
rect 94372 36728 94378 36780
rect 95234 36768 95240 36780
rect 95195 36740 95240 36768
rect 95234 36728 95240 36740
rect 95292 36728 95298 36780
rect 95878 36728 95884 36780
rect 95936 36768 95942 36780
rect 95973 36771 96031 36777
rect 95973 36768 95985 36771
rect 95936 36740 95985 36768
rect 95936 36728 95942 36740
rect 95973 36737 95985 36740
rect 96019 36737 96031 36771
rect 96080 36768 96108 36808
rect 96706 36796 96712 36848
rect 96764 36836 96770 36848
rect 96985 36839 97043 36845
rect 96985 36836 96997 36839
rect 96764 36808 96997 36836
rect 96764 36796 96770 36808
rect 96985 36805 96997 36808
rect 97031 36805 97043 36839
rect 98546 36836 98552 36848
rect 96985 36799 97043 36805
rect 97092 36808 98552 36836
rect 97092 36768 97120 36808
rect 98546 36796 98552 36808
rect 98604 36796 98610 36848
rect 98730 36796 98736 36848
rect 98788 36836 98794 36848
rect 99374 36836 99380 36848
rect 98788 36808 99380 36836
rect 98788 36796 98794 36808
rect 99374 36796 99380 36808
rect 99432 36796 99438 36848
rect 99834 36836 99840 36848
rect 99795 36808 99840 36836
rect 99834 36796 99840 36808
rect 99892 36796 99898 36848
rect 102870 36796 102876 36848
rect 102928 36836 102934 36848
rect 103793 36839 103851 36845
rect 103793 36836 103805 36839
rect 102928 36808 103805 36836
rect 102928 36796 102934 36808
rect 103793 36805 103805 36808
rect 103839 36805 103851 36839
rect 103793 36799 103851 36805
rect 105262 36796 105268 36848
rect 105320 36836 105326 36848
rect 105357 36839 105415 36845
rect 105357 36836 105369 36839
rect 105320 36808 105369 36836
rect 105320 36796 105326 36808
rect 105357 36805 105369 36808
rect 105403 36805 105415 36839
rect 105357 36799 105415 36805
rect 105541 36839 105599 36845
rect 105541 36805 105553 36839
rect 105587 36836 105599 36839
rect 106458 36836 106464 36848
rect 105587 36808 106464 36836
rect 105587 36805 105599 36808
rect 105541 36799 105599 36805
rect 106458 36796 106464 36808
rect 106516 36836 106522 36848
rect 106516 36808 106872 36836
rect 106516 36796 106522 36808
rect 96080 36740 97120 36768
rect 95973 36731 96031 36737
rect 97994 36728 98000 36780
rect 98052 36768 98058 36780
rect 98457 36772 98515 36777
rect 98288 36771 98515 36772
rect 98288 36768 98469 36771
rect 98052 36744 98469 36768
rect 98052 36740 98316 36744
rect 98052 36728 98058 36740
rect 98457 36737 98469 36744
rect 98503 36737 98515 36771
rect 98457 36731 98515 36737
rect 100754 36728 100760 36780
rect 100812 36768 100818 36780
rect 101217 36771 101275 36777
rect 101217 36768 101229 36771
rect 100812 36740 101229 36768
rect 100812 36728 100818 36740
rect 101217 36737 101229 36740
rect 101263 36737 101275 36771
rect 103054 36768 103060 36780
rect 103015 36740 103060 36768
rect 101217 36731 101275 36737
rect 103054 36728 103060 36740
rect 103112 36728 103118 36780
rect 106366 36768 106372 36780
rect 106327 36740 106372 36768
rect 106366 36728 106372 36740
rect 106424 36728 106430 36780
rect 106844 36777 106872 36808
rect 107286 36796 107292 36848
rect 107344 36836 107350 36848
rect 108025 36839 108083 36845
rect 108025 36836 108037 36839
rect 107344 36808 108037 36836
rect 107344 36796 107350 36808
rect 108025 36805 108037 36808
rect 108071 36805 108083 36839
rect 108025 36799 108083 36805
rect 108482 36796 108488 36848
rect 108540 36836 108546 36848
rect 108577 36839 108635 36845
rect 108577 36836 108589 36839
rect 108540 36808 108589 36836
rect 108540 36796 108546 36808
rect 108577 36805 108589 36808
rect 108623 36805 108635 36839
rect 112530 36836 112536 36848
rect 108577 36799 108635 36805
rect 108776 36808 112536 36836
rect 106829 36771 106887 36777
rect 106829 36737 106841 36771
rect 106875 36768 106887 36771
rect 107473 36771 107531 36777
rect 107473 36768 107485 36771
rect 106875 36740 107485 36768
rect 106875 36737 106887 36740
rect 106829 36731 106887 36737
rect 107473 36737 107485 36740
rect 107519 36737 107531 36771
rect 107473 36731 107531 36737
rect 107562 36728 107568 36780
rect 107620 36768 107626 36780
rect 108776 36768 108804 36808
rect 112530 36796 112536 36808
rect 112588 36796 112594 36848
rect 112625 36839 112683 36845
rect 112625 36805 112637 36839
rect 112671 36836 112683 36839
rect 113269 36839 113327 36845
rect 113269 36836 113281 36839
rect 112671 36808 113281 36836
rect 112671 36805 112683 36808
rect 112625 36799 112683 36805
rect 113269 36805 113281 36808
rect 113315 36836 113327 36839
rect 113315 36808 115980 36836
rect 113315 36805 113327 36808
rect 113269 36799 113327 36805
rect 107620 36740 108804 36768
rect 107620 36728 107626 36740
rect 110506 36728 110512 36780
rect 110564 36768 110570 36780
rect 110785 36771 110843 36777
rect 110785 36768 110797 36771
rect 110564 36740 110797 36768
rect 110564 36728 110570 36740
rect 110785 36737 110797 36740
rect 110831 36768 110843 36771
rect 111429 36771 111487 36777
rect 111429 36768 111441 36771
rect 110831 36740 111441 36768
rect 110831 36737 110843 36740
rect 110785 36731 110843 36737
rect 111429 36737 111441 36740
rect 111475 36737 111487 36771
rect 111429 36731 111487 36737
rect 112070 36728 112076 36780
rect 112128 36768 112134 36780
rect 112441 36771 112499 36777
rect 112441 36768 112453 36771
rect 112128 36740 112453 36768
rect 112128 36728 112134 36740
rect 112441 36737 112453 36740
rect 112487 36737 112499 36771
rect 113726 36768 113732 36780
rect 113687 36740 113732 36768
rect 112441 36731 112499 36737
rect 113726 36728 113732 36740
rect 113784 36728 113790 36780
rect 113913 36771 113971 36777
rect 113913 36737 113925 36771
rect 113959 36768 113971 36771
rect 114646 36768 114652 36780
rect 113959 36740 114652 36768
rect 113959 36737 113971 36740
rect 113913 36731 113971 36737
rect 114646 36728 114652 36740
rect 114704 36768 114710 36780
rect 115017 36771 115075 36777
rect 115017 36768 115029 36771
rect 114704 36740 115029 36768
rect 114704 36728 114710 36740
rect 115017 36737 115029 36740
rect 115063 36768 115075 36771
rect 115661 36771 115719 36777
rect 115661 36768 115673 36771
rect 115063 36740 115673 36768
rect 115063 36737 115075 36740
rect 115017 36731 115075 36737
rect 115661 36737 115673 36740
rect 115707 36737 115719 36771
rect 115661 36731 115719 36737
rect 76708 36672 80284 36700
rect 80333 36703 80391 36709
rect 76708 36660 76714 36672
rect 80333 36669 80345 36703
rect 80379 36700 80391 36703
rect 80790 36700 80796 36712
rect 80379 36672 80796 36700
rect 80379 36669 80391 36672
rect 80333 36663 80391 36669
rect 80790 36660 80796 36672
rect 80848 36700 80854 36712
rect 80977 36703 81035 36709
rect 80977 36700 80989 36703
rect 80848 36672 80989 36700
rect 80848 36660 80854 36672
rect 80977 36669 80989 36672
rect 81023 36669 81035 36703
rect 80977 36663 81035 36669
rect 81161 36703 81219 36709
rect 81161 36669 81173 36703
rect 81207 36700 81219 36703
rect 81894 36700 81900 36712
rect 81207 36672 81900 36700
rect 81207 36669 81219 36672
rect 81161 36663 81219 36669
rect 81894 36660 81900 36672
rect 81952 36660 81958 36712
rect 84838 36660 84844 36712
rect 84896 36700 84902 36712
rect 85669 36703 85727 36709
rect 85669 36700 85681 36703
rect 84896 36672 85681 36700
rect 84896 36660 84902 36672
rect 85669 36669 85681 36672
rect 85715 36669 85727 36703
rect 85669 36663 85727 36669
rect 85758 36660 85764 36712
rect 85816 36700 85822 36712
rect 108298 36700 108304 36712
rect 85816 36672 108304 36700
rect 85816 36660 85822 36672
rect 108298 36660 108304 36672
rect 108356 36660 108362 36712
rect 115952 36700 115980 36808
rect 116118 36796 116124 36848
rect 116176 36836 116182 36848
rect 116213 36839 116271 36845
rect 116213 36836 116225 36839
rect 116176 36808 116225 36836
rect 116176 36796 116182 36808
rect 116213 36805 116225 36808
rect 116259 36805 116271 36839
rect 116213 36799 116271 36805
rect 116302 36796 116308 36848
rect 116360 36836 116366 36848
rect 132126 36836 132132 36848
rect 116360 36808 128354 36836
rect 116360 36796 116366 36808
rect 116026 36728 116032 36780
rect 116084 36768 116090 36780
rect 117130 36768 117136 36780
rect 116084 36740 117136 36768
rect 116084 36728 116090 36740
rect 117130 36728 117136 36740
rect 117188 36728 117194 36780
rect 117866 36768 117872 36780
rect 117827 36740 117872 36768
rect 117866 36728 117872 36740
rect 117924 36728 117930 36780
rect 118053 36771 118111 36777
rect 118053 36737 118065 36771
rect 118099 36768 118111 36771
rect 118694 36768 118700 36780
rect 118099 36740 118700 36768
rect 118099 36737 118111 36740
rect 118053 36731 118111 36737
rect 118694 36728 118700 36740
rect 118752 36768 118758 36780
rect 119982 36768 119988 36780
rect 118752 36740 119988 36768
rect 118752 36728 118758 36740
rect 119982 36728 119988 36740
rect 120040 36728 120046 36780
rect 120997 36771 121055 36777
rect 120997 36737 121009 36771
rect 121043 36768 121055 36771
rect 121362 36768 121368 36780
rect 121043 36740 121368 36768
rect 121043 36737 121055 36740
rect 120997 36731 121055 36737
rect 121362 36728 121368 36740
rect 121420 36768 121426 36780
rect 121457 36771 121515 36777
rect 121457 36768 121469 36771
rect 121420 36740 121469 36768
rect 121420 36728 121426 36740
rect 121457 36737 121469 36740
rect 121503 36737 121515 36771
rect 121457 36731 121515 36737
rect 122834 36728 122840 36780
rect 122892 36768 122898 36780
rect 123205 36771 123263 36777
rect 123205 36768 123217 36771
rect 122892 36740 123217 36768
rect 122892 36728 122898 36740
rect 123205 36737 123217 36740
rect 123251 36768 123263 36771
rect 123849 36771 123907 36777
rect 123849 36768 123861 36771
rect 123251 36740 123861 36768
rect 123251 36737 123263 36740
rect 123205 36731 123263 36737
rect 123849 36737 123861 36740
rect 123895 36737 123907 36771
rect 123849 36731 123907 36737
rect 126701 36771 126759 36777
rect 126701 36737 126713 36771
rect 126747 36768 126759 36771
rect 126974 36768 126980 36780
rect 126747 36740 126980 36768
rect 126747 36737 126759 36740
rect 126701 36731 126759 36737
rect 126974 36728 126980 36740
rect 127032 36728 127038 36780
rect 128326 36768 128354 36808
rect 129200 36808 131068 36836
rect 129200 36768 129228 36808
rect 129550 36768 129556 36780
rect 128326 36740 129228 36768
rect 129511 36740 129556 36768
rect 129550 36728 129556 36740
rect 129608 36728 129614 36780
rect 130473 36771 130531 36777
rect 130473 36737 130485 36771
rect 130519 36768 130531 36771
rect 130930 36768 130936 36780
rect 130519 36740 130936 36768
rect 130519 36737 130531 36740
rect 130473 36731 130531 36737
rect 130930 36728 130936 36740
rect 130988 36728 130994 36780
rect 131040 36768 131068 36808
rect 131132 36808 132132 36836
rect 131132 36768 131160 36808
rect 132126 36796 132132 36808
rect 132184 36796 132190 36848
rect 132466 36836 132494 36876
rect 133230 36864 133236 36876
rect 133288 36864 133294 36916
rect 134242 36904 134248 36916
rect 134203 36876 134248 36904
rect 134242 36864 134248 36876
rect 134300 36864 134306 36916
rect 135990 36904 135996 36916
rect 135951 36876 135996 36904
rect 135990 36864 135996 36876
rect 136048 36864 136054 36916
rect 137833 36907 137891 36913
rect 137833 36873 137845 36907
rect 137879 36904 137891 36907
rect 138934 36904 138940 36916
rect 137879 36876 138940 36904
rect 137879 36873 137891 36876
rect 137833 36867 137891 36873
rect 138934 36864 138940 36876
rect 138992 36864 138998 36916
rect 140498 36904 140504 36916
rect 140459 36876 140504 36904
rect 140498 36864 140504 36876
rect 140556 36864 140562 36916
rect 141605 36907 141663 36913
rect 141605 36873 141617 36907
rect 141651 36904 141663 36907
rect 143074 36904 143080 36916
rect 141651 36876 143080 36904
rect 141651 36873 141663 36876
rect 141605 36867 141663 36873
rect 143074 36864 143080 36876
rect 143132 36864 143138 36916
rect 143813 36907 143871 36913
rect 143813 36873 143825 36907
rect 143859 36904 143871 36907
rect 144546 36904 144552 36916
rect 143859 36876 144552 36904
rect 143859 36873 143871 36876
rect 143813 36867 143871 36873
rect 144546 36864 144552 36876
rect 144604 36864 144610 36916
rect 145101 36907 145159 36913
rect 145101 36873 145113 36907
rect 145147 36904 145159 36907
rect 145282 36904 145288 36916
rect 145147 36876 145288 36904
rect 145147 36873 145159 36876
rect 145101 36867 145159 36873
rect 145282 36864 145288 36876
rect 145340 36864 145346 36916
rect 146294 36904 146300 36916
rect 146255 36876 146300 36904
rect 146294 36864 146300 36876
rect 146352 36864 146358 36916
rect 147122 36864 147128 36916
rect 147180 36904 147186 36916
rect 147309 36907 147367 36913
rect 147309 36904 147321 36907
rect 147180 36876 147321 36904
rect 147180 36864 147186 36876
rect 147309 36873 147321 36876
rect 147355 36873 147367 36907
rect 147309 36867 147367 36873
rect 133506 36836 133512 36848
rect 132466 36808 133512 36836
rect 133506 36796 133512 36808
rect 133564 36796 133570 36848
rect 137278 36796 137284 36848
rect 137336 36836 137342 36848
rect 142154 36836 142160 36848
rect 137336 36808 142160 36836
rect 137336 36796 137342 36808
rect 142154 36796 142160 36808
rect 142212 36796 142218 36848
rect 142246 36796 142252 36848
rect 142304 36836 142310 36848
rect 142617 36839 142675 36845
rect 142617 36836 142629 36839
rect 142304 36808 142629 36836
rect 142304 36796 142310 36808
rect 142617 36805 142629 36808
rect 142663 36805 142675 36839
rect 142617 36799 142675 36805
rect 132034 36768 132040 36780
rect 131040 36740 131160 36768
rect 131995 36740 132040 36768
rect 132034 36728 132040 36740
rect 132092 36768 132098 36780
rect 132681 36771 132739 36777
rect 132681 36768 132693 36771
rect 132092 36740 132693 36768
rect 132092 36728 132098 36740
rect 132681 36737 132693 36740
rect 132727 36737 132739 36771
rect 135809 36771 135867 36777
rect 135809 36768 135821 36771
rect 132681 36731 132739 36737
rect 134904 36740 135821 36768
rect 123294 36700 123300 36712
rect 111076 36672 112576 36700
rect 115952 36672 123300 36700
rect 71314 36632 71320 36644
rect 65720 36604 71320 36632
rect 51868 36536 53144 36564
rect 53653 36567 53711 36573
rect 51868 36524 51874 36536
rect 53653 36533 53665 36567
rect 53699 36564 53711 36567
rect 53742 36564 53748 36576
rect 53699 36536 53748 36564
rect 53699 36533 53711 36536
rect 53653 36527 53711 36533
rect 53742 36524 53748 36536
rect 53800 36524 53806 36576
rect 54386 36564 54392 36576
rect 54347 36536 54392 36564
rect 54386 36524 54392 36536
rect 54444 36524 54450 36576
rect 55122 36564 55128 36576
rect 55083 36536 55128 36564
rect 55122 36524 55128 36536
rect 55180 36524 55186 36576
rect 56505 36567 56563 36573
rect 56505 36533 56517 36567
rect 56551 36564 56563 36567
rect 56686 36564 56692 36576
rect 56551 36536 56692 36564
rect 56551 36533 56563 36536
rect 56505 36527 56563 36533
rect 56686 36524 56692 36536
rect 56744 36524 56750 36576
rect 57054 36564 57060 36576
rect 57015 36536 57060 36564
rect 57054 36524 57060 36536
rect 57112 36524 57118 36576
rect 58805 36567 58863 36573
rect 58805 36533 58817 36567
rect 58851 36564 58863 36567
rect 59078 36564 59084 36576
rect 58851 36536 59084 36564
rect 58851 36533 58863 36536
rect 58805 36527 58863 36533
rect 59078 36524 59084 36536
rect 59136 36524 59142 36576
rect 61010 36564 61016 36576
rect 60971 36536 61016 36564
rect 61010 36524 61016 36536
rect 61068 36524 61074 36576
rect 63310 36524 63316 36576
rect 63368 36564 63374 36576
rect 63405 36567 63463 36573
rect 63405 36564 63417 36567
rect 63368 36536 63417 36564
rect 63368 36524 63374 36536
rect 63405 36533 63417 36536
rect 63451 36533 63463 36567
rect 63405 36527 63463 36533
rect 63494 36524 63500 36576
rect 63552 36564 63558 36576
rect 63865 36567 63923 36573
rect 63865 36564 63877 36567
rect 63552 36536 63877 36564
rect 63552 36524 63558 36536
rect 63865 36533 63877 36536
rect 63911 36533 63923 36567
rect 63865 36527 63923 36533
rect 63954 36524 63960 36576
rect 64012 36564 64018 36576
rect 64782 36564 64788 36576
rect 64012 36536 64788 36564
rect 64012 36524 64018 36536
rect 64782 36524 64788 36536
rect 64840 36524 64846 36576
rect 64874 36524 64880 36576
rect 64932 36564 64938 36576
rect 65352 36564 65380 36604
rect 71314 36592 71320 36604
rect 71372 36592 71378 36644
rect 73617 36635 73675 36641
rect 73617 36601 73629 36635
rect 73663 36632 73675 36635
rect 73798 36632 73804 36644
rect 73663 36604 73804 36632
rect 73663 36601 73675 36604
rect 73617 36595 73675 36601
rect 73798 36592 73804 36604
rect 73856 36632 73862 36644
rect 74626 36632 74632 36644
rect 73856 36604 74632 36632
rect 73856 36592 73862 36604
rect 74626 36592 74632 36604
rect 74684 36592 74690 36644
rect 74813 36635 74871 36641
rect 74813 36601 74825 36635
rect 74859 36632 74871 36635
rect 75270 36632 75276 36644
rect 74859 36604 75276 36632
rect 74859 36601 74871 36604
rect 74813 36595 74871 36601
rect 75270 36592 75276 36604
rect 75328 36592 75334 36644
rect 76558 36592 76564 36644
rect 76616 36632 76622 36644
rect 111076 36632 111104 36672
rect 76616 36604 80100 36632
rect 76616 36592 76622 36604
rect 64932 36536 65380 36564
rect 64932 36524 64938 36536
rect 65702 36524 65708 36576
rect 65760 36564 65766 36576
rect 65797 36567 65855 36573
rect 65797 36564 65809 36567
rect 65760 36536 65809 36564
rect 65760 36524 65766 36536
rect 65797 36533 65809 36536
rect 65843 36533 65855 36567
rect 65797 36527 65855 36533
rect 66254 36524 66260 36576
rect 66312 36564 66318 36576
rect 70854 36564 70860 36576
rect 66312 36536 70860 36564
rect 66312 36524 66318 36536
rect 70854 36524 70860 36536
rect 70912 36524 70918 36576
rect 71038 36564 71044 36576
rect 70999 36536 71044 36564
rect 71038 36524 71044 36536
rect 71096 36524 71102 36576
rect 71682 36564 71688 36576
rect 71643 36536 71688 36564
rect 71682 36524 71688 36536
rect 71740 36524 71746 36576
rect 73982 36524 73988 36576
rect 74040 36564 74046 36576
rect 74077 36567 74135 36573
rect 74077 36564 74089 36567
rect 74040 36536 74089 36564
rect 74040 36524 74046 36536
rect 74077 36533 74089 36536
rect 74123 36564 74135 36567
rect 75365 36567 75423 36573
rect 75365 36564 75377 36567
rect 74123 36536 75377 36564
rect 74123 36533 74135 36536
rect 74077 36527 74135 36533
rect 75365 36533 75377 36536
rect 75411 36533 75423 36567
rect 75365 36527 75423 36533
rect 75733 36567 75791 36573
rect 75733 36533 75745 36567
rect 75779 36564 75791 36567
rect 76098 36564 76104 36576
rect 75779 36536 76104 36564
rect 75779 36533 75791 36536
rect 75733 36527 75791 36533
rect 76098 36524 76104 36536
rect 76156 36524 76162 36576
rect 77294 36524 77300 36576
rect 77352 36564 77358 36576
rect 77754 36564 77760 36576
rect 77352 36536 77760 36564
rect 77352 36524 77358 36536
rect 77754 36524 77760 36536
rect 77812 36524 77818 36576
rect 79689 36567 79747 36573
rect 79689 36533 79701 36567
rect 79735 36564 79747 36567
rect 79778 36564 79784 36576
rect 79735 36536 79784 36564
rect 79735 36533 79747 36536
rect 79689 36527 79747 36533
rect 79778 36524 79784 36536
rect 79836 36524 79842 36576
rect 80072 36564 80100 36604
rect 80256 36604 111104 36632
rect 112548 36632 112576 36672
rect 123294 36660 123300 36672
rect 123352 36660 123358 36712
rect 134426 36700 134432 36712
rect 123404 36672 134432 36700
rect 123404 36641 123432 36672
rect 134426 36660 134432 36672
rect 134484 36660 134490 36712
rect 123389 36635 123447 36641
rect 112548 36604 123248 36632
rect 80256 36564 80284 36604
rect 80072 36536 80284 36564
rect 81621 36567 81679 36573
rect 81621 36533 81633 36567
rect 81667 36564 81679 36567
rect 82078 36564 82084 36576
rect 81667 36536 82084 36564
rect 81667 36533 81679 36536
rect 81621 36527 81679 36533
rect 82078 36524 82084 36536
rect 82136 36524 82142 36576
rect 82262 36524 82268 36576
rect 82320 36564 82326 36576
rect 82909 36567 82967 36573
rect 82909 36564 82921 36567
rect 82320 36536 82921 36564
rect 82320 36524 82326 36536
rect 82909 36533 82921 36536
rect 82955 36533 82967 36567
rect 82909 36527 82967 36533
rect 83642 36524 83648 36576
rect 83700 36564 83706 36576
rect 84013 36567 84071 36573
rect 84013 36564 84025 36567
rect 83700 36536 84025 36564
rect 83700 36524 83706 36536
rect 84013 36533 84025 36536
rect 84059 36533 84071 36567
rect 86402 36564 86408 36576
rect 86363 36536 86408 36564
rect 84013 36527 84071 36533
rect 86402 36524 86408 36536
rect 86460 36524 86466 36576
rect 86862 36524 86868 36576
rect 86920 36564 86926 36576
rect 86957 36567 87015 36573
rect 86957 36564 86969 36567
rect 86920 36536 86969 36564
rect 86920 36524 86926 36536
rect 86957 36533 86969 36536
rect 87003 36533 87015 36567
rect 88058 36564 88064 36576
rect 88019 36536 88064 36564
rect 86957 36527 87015 36533
rect 88058 36524 88064 36536
rect 88116 36524 88122 36576
rect 89162 36524 89168 36576
rect 89220 36564 89226 36576
rect 89441 36567 89499 36573
rect 89441 36564 89453 36567
rect 89220 36536 89453 36564
rect 89220 36524 89226 36536
rect 89441 36533 89453 36536
rect 89487 36533 89499 36567
rect 90450 36564 90456 36576
rect 90411 36536 90456 36564
rect 89441 36527 89499 36533
rect 90450 36524 90456 36536
rect 90508 36524 90514 36576
rect 91554 36564 91560 36576
rect 91515 36536 91560 36564
rect 91554 36524 91560 36536
rect 91612 36524 91618 36576
rect 92106 36564 92112 36576
rect 92067 36536 92112 36564
rect 92106 36524 92112 36536
rect 92164 36524 92170 36576
rect 94225 36567 94283 36573
rect 94225 36533 94237 36567
rect 94271 36564 94283 36567
rect 94314 36564 94320 36576
rect 94271 36536 94320 36564
rect 94271 36533 94283 36536
rect 94225 36527 94283 36533
rect 94314 36524 94320 36536
rect 94372 36524 94378 36576
rect 95050 36564 95056 36576
rect 95011 36536 95056 36564
rect 95050 36524 95056 36536
rect 95108 36524 95114 36576
rect 95602 36524 95608 36576
rect 95660 36564 95666 36576
rect 95789 36567 95847 36573
rect 95789 36564 95801 36567
rect 95660 36536 95801 36564
rect 95660 36524 95666 36536
rect 95789 36533 95801 36536
rect 95835 36533 95847 36567
rect 95789 36527 95847 36533
rect 96154 36524 96160 36576
rect 96212 36564 96218 36576
rect 96433 36567 96491 36573
rect 96433 36564 96445 36567
rect 96212 36536 96445 36564
rect 96212 36524 96218 36536
rect 96433 36533 96445 36536
rect 96479 36533 96491 36567
rect 97994 36564 98000 36576
rect 97955 36536 98000 36564
rect 96433 36527 96491 36533
rect 97994 36524 98000 36536
rect 98052 36524 98058 36576
rect 98638 36564 98644 36576
rect 98599 36536 98644 36564
rect 98638 36524 98644 36536
rect 98696 36524 98702 36576
rect 100754 36564 100760 36576
rect 100715 36536 100760 36564
rect 100754 36524 100760 36536
rect 100812 36524 100818 36576
rect 101122 36524 101128 36576
rect 101180 36564 101186 36576
rect 101401 36567 101459 36573
rect 101401 36564 101413 36567
rect 101180 36536 101413 36564
rect 101180 36524 101186 36536
rect 101401 36533 101413 36536
rect 101447 36533 101459 36567
rect 101401 36527 101459 36533
rect 102134 36524 102140 36576
rect 102192 36564 102198 36576
rect 102229 36567 102287 36573
rect 102229 36564 102241 36567
rect 102192 36536 102241 36564
rect 102192 36524 102198 36536
rect 102229 36533 102241 36536
rect 102275 36533 102287 36567
rect 102229 36527 102287 36533
rect 102962 36524 102968 36576
rect 103020 36564 103026 36576
rect 103241 36567 103299 36573
rect 103241 36564 103253 36567
rect 103020 36536 103253 36564
rect 103020 36524 103026 36536
rect 103241 36533 103253 36536
rect 103287 36533 103299 36567
rect 104434 36564 104440 36576
rect 104395 36536 104440 36564
rect 103241 36527 103299 36533
rect 104434 36524 104440 36536
rect 104492 36524 104498 36576
rect 105722 36524 105728 36576
rect 105780 36564 105786 36576
rect 106185 36567 106243 36573
rect 106185 36564 106197 36567
rect 105780 36536 106197 36564
rect 105780 36524 105786 36536
rect 106185 36533 106197 36536
rect 106231 36533 106243 36567
rect 106185 36527 106243 36533
rect 107013 36567 107071 36573
rect 107013 36533 107025 36567
rect 107059 36564 107071 36567
rect 109402 36564 109408 36576
rect 107059 36536 109408 36564
rect 107059 36533 107071 36536
rect 107013 36527 107071 36533
rect 109402 36524 109408 36536
rect 109460 36524 109466 36576
rect 109586 36564 109592 36576
rect 109547 36536 109592 36564
rect 109586 36524 109592 36536
rect 109644 36524 109650 36576
rect 110325 36567 110383 36573
rect 110325 36533 110337 36567
rect 110371 36564 110383 36567
rect 110506 36564 110512 36576
rect 110371 36536 110512 36564
rect 110371 36533 110383 36536
rect 110325 36527 110383 36533
rect 110506 36524 110512 36536
rect 110564 36524 110570 36576
rect 110969 36567 111027 36573
rect 110969 36533 110981 36567
rect 111015 36564 111027 36567
rect 111886 36564 111892 36576
rect 111015 36536 111892 36564
rect 111015 36533 111027 36536
rect 110969 36527 111027 36533
rect 111886 36524 111892 36536
rect 111944 36524 111950 36576
rect 115201 36567 115259 36573
rect 115201 36533 115213 36567
rect 115247 36564 115259 36567
rect 116946 36564 116952 36576
rect 115247 36536 116952 36564
rect 115247 36533 115259 36536
rect 115201 36527 115259 36533
rect 116946 36524 116952 36536
rect 117004 36524 117010 36576
rect 119154 36564 119160 36576
rect 119115 36536 119160 36564
rect 119154 36524 119160 36536
rect 119212 36524 119218 36576
rect 121454 36524 121460 36576
rect 121512 36564 121518 36576
rect 121641 36567 121699 36573
rect 121641 36564 121653 36567
rect 121512 36536 121653 36564
rect 121512 36524 121518 36536
rect 121641 36533 121653 36536
rect 121687 36533 121699 36567
rect 121641 36527 121699 36533
rect 122745 36567 122803 36573
rect 122745 36533 122757 36567
rect 122791 36564 122803 36567
rect 122834 36564 122840 36576
rect 122791 36536 122840 36564
rect 122791 36533 122803 36536
rect 122745 36527 122803 36533
rect 122834 36524 122840 36536
rect 122892 36524 122898 36576
rect 123220 36564 123248 36604
rect 123389 36601 123401 36635
rect 123435 36601 123447 36635
rect 127802 36632 127808 36644
rect 123389 36595 123447 36601
rect 123496 36604 127808 36632
rect 123496 36564 123524 36604
rect 127802 36592 127808 36604
rect 127860 36592 127866 36644
rect 134904 36632 134932 36740
rect 135809 36737 135821 36740
rect 135855 36768 135867 36771
rect 136453 36771 136511 36777
rect 136453 36768 136465 36771
rect 135855 36740 136465 36768
rect 135855 36737 135867 36740
rect 135809 36731 135867 36737
rect 136453 36737 136465 36740
rect 136499 36737 136511 36771
rect 137646 36768 137652 36780
rect 137607 36740 137652 36768
rect 136453 36731 136511 36737
rect 137646 36728 137652 36740
rect 137704 36768 137710 36780
rect 138293 36771 138351 36777
rect 138293 36768 138305 36771
rect 137704 36740 138305 36768
rect 137704 36728 137710 36740
rect 138293 36737 138305 36740
rect 138339 36737 138351 36771
rect 138293 36731 138351 36737
rect 141421 36771 141479 36777
rect 141421 36737 141433 36771
rect 141467 36737 141479 36771
rect 143626 36768 143632 36780
rect 143539 36740 143632 36768
rect 141421 36731 141479 36737
rect 135898 36660 135904 36712
rect 135956 36700 135962 36712
rect 141326 36700 141332 36712
rect 135956 36672 141332 36700
rect 135956 36660 135962 36672
rect 141326 36660 141332 36672
rect 141384 36700 141390 36712
rect 141436 36700 141464 36731
rect 143626 36728 143632 36740
rect 143684 36768 143690 36780
rect 144273 36771 144331 36777
rect 144273 36768 144285 36771
rect 143684 36740 144285 36768
rect 143684 36728 143690 36740
rect 144273 36737 144285 36740
rect 144319 36737 144331 36771
rect 144273 36731 144331 36737
rect 146113 36771 146171 36777
rect 146113 36737 146125 36771
rect 146159 36768 146171 36771
rect 146294 36768 146300 36780
rect 146159 36740 146300 36768
rect 146159 36737 146171 36740
rect 146113 36731 146171 36737
rect 146294 36728 146300 36740
rect 146352 36768 146358 36780
rect 146757 36771 146815 36777
rect 146757 36768 146769 36771
rect 146352 36740 146769 36768
rect 146352 36728 146358 36740
rect 146757 36737 146769 36740
rect 146803 36737 146815 36771
rect 146757 36731 146815 36737
rect 142065 36703 142123 36709
rect 142065 36700 142077 36703
rect 141384 36672 142077 36700
rect 141384 36660 141390 36672
rect 142065 36669 142077 36672
rect 142111 36669 142123 36703
rect 142065 36663 142123 36669
rect 128326 36604 134932 36632
rect 123220 36536 123524 36564
rect 123570 36524 123576 36576
rect 123628 36564 123634 36576
rect 126514 36564 126520 36576
rect 123628 36536 126520 36564
rect 123628 36524 123634 36536
rect 126514 36524 126520 36536
rect 126572 36524 126578 36576
rect 126974 36524 126980 36576
rect 127032 36564 127038 36576
rect 127161 36567 127219 36573
rect 127161 36564 127173 36567
rect 127032 36536 127173 36564
rect 127032 36524 127038 36536
rect 127161 36533 127173 36536
rect 127207 36564 127219 36567
rect 128326 36564 128354 36604
rect 130286 36564 130292 36576
rect 127207 36536 128354 36564
rect 130247 36536 130292 36564
rect 127207 36533 127219 36536
rect 127161 36527 127219 36533
rect 130286 36524 130292 36536
rect 130344 36524 130350 36576
rect 130930 36564 130936 36576
rect 130891 36536 130936 36564
rect 130930 36524 130936 36536
rect 130988 36524 130994 36576
rect 139486 36564 139492 36576
rect 139447 36536 139492 36564
rect 139486 36524 139492 36536
rect 139544 36524 139550 36576
rect 1104 36474 148856 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 65654 36474
rect 65706 36422 65718 36474
rect 65770 36422 65782 36474
rect 65834 36422 65846 36474
rect 65898 36422 65910 36474
rect 65962 36422 96374 36474
rect 96426 36422 96438 36474
rect 96490 36422 96502 36474
rect 96554 36422 96566 36474
rect 96618 36422 96630 36474
rect 96682 36422 127094 36474
rect 127146 36422 127158 36474
rect 127210 36422 127222 36474
rect 127274 36422 127286 36474
rect 127338 36422 127350 36474
rect 127402 36422 148856 36474
rect 1104 36400 148856 36422
rect 10042 36360 10048 36372
rect 10003 36332 10048 36360
rect 10042 36320 10048 36332
rect 10100 36320 10106 36372
rect 17402 36360 17408 36372
rect 17363 36332 17408 36360
rect 17402 36320 17408 36332
rect 17460 36320 17466 36372
rect 17770 36320 17776 36372
rect 17828 36360 17834 36372
rect 22462 36360 22468 36372
rect 17828 36332 22094 36360
rect 22423 36332 22468 36360
rect 17828 36320 17834 36332
rect 21726 36292 21732 36304
rect 14936 36264 21732 36292
rect 10502 36184 10508 36236
rect 10560 36224 10566 36236
rect 14826 36224 14832 36236
rect 10560 36196 14832 36224
rect 10560 36184 10566 36196
rect 14826 36184 14832 36196
rect 14884 36184 14890 36236
rect 10318 36116 10324 36168
rect 10376 36156 10382 36168
rect 14936 36156 14964 36264
rect 21726 36252 21732 36264
rect 21784 36252 21790 36304
rect 22066 36292 22094 36332
rect 22462 36320 22468 36332
rect 22520 36320 22526 36372
rect 23474 36360 23480 36372
rect 23435 36332 23480 36360
rect 23474 36320 23480 36332
rect 23532 36320 23538 36372
rect 24118 36360 24124 36372
rect 23952 36332 24124 36360
rect 23952 36292 23980 36332
rect 24118 36320 24124 36332
rect 24176 36320 24182 36372
rect 24854 36320 24860 36372
rect 24912 36360 24918 36372
rect 24949 36363 25007 36369
rect 24949 36360 24961 36363
rect 24912 36332 24961 36360
rect 24912 36320 24918 36332
rect 24949 36329 24961 36332
rect 24995 36329 25007 36363
rect 24949 36323 25007 36329
rect 25682 36320 25688 36372
rect 25740 36360 25746 36372
rect 25869 36363 25927 36369
rect 25869 36360 25881 36363
rect 25740 36332 25881 36360
rect 25740 36320 25746 36332
rect 25869 36329 25881 36332
rect 25915 36329 25927 36363
rect 25869 36323 25927 36329
rect 27614 36320 27620 36372
rect 27672 36360 27678 36372
rect 27709 36363 27767 36369
rect 27709 36360 27721 36363
rect 27672 36332 27721 36360
rect 27672 36320 27678 36332
rect 27709 36329 27721 36332
rect 27755 36329 27767 36363
rect 27709 36323 27767 36329
rect 29362 36320 29368 36372
rect 29420 36360 29426 36372
rect 29733 36363 29791 36369
rect 29733 36360 29745 36363
rect 29420 36332 29745 36360
rect 29420 36320 29426 36332
rect 29733 36329 29745 36332
rect 29779 36329 29791 36363
rect 29733 36323 29791 36329
rect 30650 36320 30656 36372
rect 30708 36360 30714 36372
rect 30745 36363 30803 36369
rect 30745 36360 30757 36363
rect 30708 36332 30757 36360
rect 30708 36320 30714 36332
rect 30745 36329 30757 36332
rect 30791 36329 30803 36363
rect 30745 36323 30803 36329
rect 32306 36320 32312 36372
rect 32364 36360 32370 36372
rect 33686 36360 33692 36372
rect 32364 36332 33692 36360
rect 32364 36320 32370 36332
rect 33686 36320 33692 36332
rect 33744 36320 33750 36372
rect 33781 36363 33839 36369
rect 33781 36329 33793 36363
rect 33827 36360 33839 36363
rect 33962 36360 33968 36372
rect 33827 36332 33968 36360
rect 33827 36329 33839 36332
rect 33781 36323 33839 36329
rect 33962 36320 33968 36332
rect 34020 36320 34026 36372
rect 36538 36360 36544 36372
rect 34164 36332 36544 36360
rect 22066 36264 23980 36292
rect 24029 36295 24087 36301
rect 24029 36261 24041 36295
rect 24075 36292 24087 36295
rect 25130 36292 25136 36304
rect 24075 36264 25136 36292
rect 24075 36261 24087 36264
rect 24029 36255 24087 36261
rect 25130 36252 25136 36264
rect 25188 36252 25194 36304
rect 25406 36252 25412 36304
rect 25464 36292 25470 36304
rect 26326 36292 26332 36304
rect 25464 36264 26332 36292
rect 25464 36252 25470 36264
rect 26326 36252 26332 36264
rect 26384 36252 26390 36304
rect 34164 36292 34192 36332
rect 36538 36320 36544 36332
rect 36596 36320 36602 36372
rect 39298 36360 39304 36372
rect 37292 36332 39304 36360
rect 37292 36304 37320 36332
rect 39298 36320 39304 36332
rect 39356 36320 39362 36372
rect 39482 36360 39488 36372
rect 39443 36332 39488 36360
rect 39482 36320 39488 36332
rect 39540 36320 39546 36372
rect 39684 36332 41736 36360
rect 26436 36264 34192 36292
rect 17954 36184 17960 36236
rect 18012 36224 18018 36236
rect 18012 36196 22094 36224
rect 18012 36184 18018 36196
rect 10376 36128 14964 36156
rect 10376 36116 10382 36128
rect 15010 36116 15016 36168
rect 15068 36156 15074 36168
rect 15068 36128 15240 36156
rect 15068 36116 15074 36128
rect 6914 36048 6920 36100
rect 6972 36088 6978 36100
rect 14458 36088 14464 36100
rect 6972 36060 14464 36088
rect 6972 36048 6978 36060
rect 14458 36048 14464 36060
rect 14516 36088 14522 36100
rect 15102 36088 15108 36100
rect 14516 36060 15108 36088
rect 14516 36048 14522 36060
rect 15102 36048 15108 36060
rect 15160 36048 15166 36100
rect 15212 36088 15240 36128
rect 15470 36116 15476 36168
rect 15528 36156 15534 36168
rect 19518 36156 19524 36168
rect 15528 36128 19524 36156
rect 15528 36116 15534 36128
rect 19518 36116 19524 36128
rect 19576 36116 19582 36168
rect 20162 36156 20168 36168
rect 20123 36128 20168 36156
rect 20162 36116 20168 36128
rect 20220 36116 20226 36168
rect 21082 36116 21088 36168
rect 21140 36156 21146 36168
rect 21177 36159 21235 36165
rect 21177 36156 21189 36159
rect 21140 36128 21189 36156
rect 21140 36116 21146 36128
rect 21177 36125 21189 36128
rect 21223 36125 21235 36159
rect 21818 36156 21824 36168
rect 21177 36119 21235 36125
rect 21284 36128 21824 36156
rect 19426 36088 19432 36100
rect 15212 36060 19432 36088
rect 19426 36048 19432 36060
rect 19484 36048 19490 36100
rect 19613 36091 19671 36097
rect 19613 36057 19625 36091
rect 19659 36088 19671 36091
rect 20714 36088 20720 36100
rect 19659 36060 20720 36088
rect 19659 36057 19671 36060
rect 19613 36051 19671 36057
rect 20714 36048 20720 36060
rect 20772 36088 20778 36100
rect 21284 36088 21312 36128
rect 21818 36116 21824 36128
rect 21876 36116 21882 36168
rect 22066 36156 22094 36196
rect 23934 36184 23940 36236
rect 23992 36224 23998 36236
rect 26436 36224 26464 36264
rect 34238 36252 34244 36304
rect 34296 36292 34302 36304
rect 36081 36295 36139 36301
rect 34296 36264 34341 36292
rect 34296 36252 34302 36264
rect 36081 36261 36093 36295
rect 36127 36292 36139 36295
rect 36354 36292 36360 36304
rect 36127 36264 36360 36292
rect 36127 36261 36139 36264
rect 36081 36255 36139 36261
rect 36354 36252 36360 36264
rect 36412 36252 36418 36304
rect 37274 36292 37280 36304
rect 36464 36264 37280 36292
rect 34422 36224 34428 36236
rect 23992 36196 26464 36224
rect 26528 36196 34428 36224
rect 23992 36184 23998 36196
rect 25130 36156 25136 36168
rect 22066 36128 24164 36156
rect 25091 36128 25136 36156
rect 24136 36088 24164 36128
rect 25130 36116 25136 36128
rect 25188 36116 25194 36168
rect 26053 36159 26111 36165
rect 26053 36125 26065 36159
rect 26099 36156 26111 36159
rect 26528 36156 26556 36196
rect 34422 36184 34428 36196
rect 34480 36184 34486 36236
rect 34606 36184 34612 36236
rect 34664 36224 34670 36236
rect 36464 36224 36492 36264
rect 37274 36252 37280 36264
rect 37332 36252 37338 36304
rect 37921 36295 37979 36301
rect 37921 36261 37933 36295
rect 37967 36292 37979 36295
rect 39684 36292 39712 36332
rect 37967 36264 39712 36292
rect 41601 36295 41659 36301
rect 37967 36261 37979 36264
rect 37921 36255 37979 36261
rect 41601 36261 41613 36295
rect 41647 36261 41659 36295
rect 41708 36292 41736 36332
rect 42242 36320 42248 36372
rect 42300 36360 42306 36372
rect 42429 36363 42487 36369
rect 42429 36360 42441 36363
rect 42300 36332 42441 36360
rect 42300 36320 42306 36332
rect 42429 36329 42441 36332
rect 42475 36329 42487 36363
rect 42429 36323 42487 36329
rect 42886 36320 42892 36372
rect 42944 36360 42950 36372
rect 43441 36363 43499 36369
rect 43441 36360 43453 36363
rect 42944 36332 43453 36360
rect 42944 36320 42950 36332
rect 43441 36329 43453 36332
rect 43487 36329 43499 36363
rect 43441 36323 43499 36329
rect 44269 36363 44327 36369
rect 44269 36329 44281 36363
rect 44315 36360 44327 36363
rect 44315 36332 53328 36360
rect 44315 36329 44327 36332
rect 44269 36323 44327 36329
rect 47302 36292 47308 36304
rect 41708 36264 47308 36292
rect 41601 36255 41659 36261
rect 34664 36196 36492 36224
rect 34664 36184 34670 36196
rect 36538 36184 36544 36236
rect 36596 36224 36602 36236
rect 39942 36224 39948 36236
rect 36596 36196 39948 36224
rect 36596 36184 36602 36196
rect 39942 36184 39948 36196
rect 40000 36184 40006 36236
rect 41506 36224 41512 36236
rect 40144 36196 41512 36224
rect 26099 36128 26556 36156
rect 26099 36125 26111 36128
rect 26053 36119 26111 36125
rect 26602 36116 26608 36168
rect 26660 36156 26666 36168
rect 26697 36159 26755 36165
rect 26697 36156 26709 36159
rect 26660 36128 26709 36156
rect 26660 36116 26666 36128
rect 26697 36125 26709 36128
rect 26743 36125 26755 36159
rect 27890 36156 27896 36168
rect 27851 36128 27896 36156
rect 26697 36119 26755 36125
rect 27890 36116 27896 36128
rect 27948 36116 27954 36168
rect 30834 36156 30840 36168
rect 28368 36128 30840 36156
rect 25406 36088 25412 36100
rect 20772 36060 21312 36088
rect 21376 36060 24072 36088
rect 24136 36060 25412 36088
rect 20772 36048 20778 36060
rect 8570 35980 8576 36032
rect 8628 36020 8634 36032
rect 9217 36023 9275 36029
rect 9217 36020 9229 36023
rect 8628 35992 9229 36020
rect 8628 35980 8634 35992
rect 9217 35989 9229 35992
rect 9263 36020 9275 36023
rect 14734 36020 14740 36032
rect 9263 35992 14740 36020
rect 9263 35989 9275 35992
rect 9217 35983 9275 35989
rect 14734 35980 14740 35992
rect 14792 35980 14798 36032
rect 14826 35980 14832 36032
rect 14884 36020 14890 36032
rect 20530 36020 20536 36032
rect 14884 35992 20536 36020
rect 14884 35980 14890 35992
rect 20530 35980 20536 35992
rect 20588 35980 20594 36032
rect 20625 36023 20683 36029
rect 20625 35989 20637 36023
rect 20671 36020 20683 36023
rect 21266 36020 21272 36032
rect 20671 35992 21272 36020
rect 20671 35989 20683 35992
rect 20625 35983 20683 35989
rect 21266 35980 21272 35992
rect 21324 35980 21330 36032
rect 21376 36029 21404 36060
rect 21361 36023 21419 36029
rect 21361 35989 21373 36023
rect 21407 35989 21419 36023
rect 24044 36020 24072 36060
rect 25406 36048 25412 36060
rect 25464 36048 25470 36100
rect 26326 36048 26332 36100
rect 26384 36088 26390 36100
rect 28368 36088 28396 36128
rect 30834 36116 30840 36128
rect 30892 36116 30898 36168
rect 31757 36159 31815 36165
rect 31757 36125 31769 36159
rect 31803 36156 31815 36159
rect 32122 36156 32128 36168
rect 31803 36128 32128 36156
rect 31803 36125 31815 36128
rect 31757 36119 31815 36125
rect 32122 36116 32128 36128
rect 32180 36156 32186 36168
rect 32217 36159 32275 36165
rect 32217 36156 32229 36159
rect 32180 36128 32229 36156
rect 32180 36116 32186 36128
rect 32217 36125 32229 36128
rect 32263 36125 32275 36159
rect 34698 36156 34704 36168
rect 32217 36119 32275 36125
rect 32324 36128 34704 36156
rect 32324 36088 32352 36128
rect 34698 36116 34704 36128
rect 34756 36116 34762 36168
rect 35894 36156 35900 36168
rect 35855 36128 35900 36156
rect 35894 36116 35900 36128
rect 35952 36116 35958 36168
rect 36725 36159 36783 36165
rect 36372 36128 36676 36156
rect 36372 36088 36400 36128
rect 26384 36060 28396 36088
rect 28460 36060 32352 36088
rect 32416 36060 36400 36088
rect 36648 36088 36676 36128
rect 36725 36125 36737 36159
rect 36771 36156 36783 36159
rect 37274 36156 37280 36168
rect 36771 36128 37280 36156
rect 36771 36125 36783 36128
rect 36725 36119 36783 36125
rect 37274 36116 37280 36128
rect 37332 36116 37338 36168
rect 37642 36116 37648 36168
rect 37700 36156 37706 36168
rect 37737 36159 37795 36165
rect 37737 36156 37749 36159
rect 37700 36128 37749 36156
rect 37700 36116 37706 36128
rect 37737 36125 37749 36128
rect 37783 36125 37795 36159
rect 37737 36119 37795 36125
rect 39482 36116 39488 36168
rect 39540 36156 39546 36168
rect 40037 36159 40095 36165
rect 40037 36156 40049 36159
rect 39540 36128 40049 36156
rect 39540 36116 39546 36128
rect 40037 36125 40049 36128
rect 40083 36125 40095 36159
rect 40037 36119 40095 36125
rect 40144 36088 40172 36196
rect 41506 36184 41512 36196
rect 41564 36184 41570 36236
rect 41616 36224 41644 36255
rect 47302 36252 47308 36264
rect 47360 36252 47366 36304
rect 48590 36292 48596 36304
rect 48056 36264 48596 36292
rect 46477 36227 46535 36233
rect 41616 36196 45554 36224
rect 40957 36159 41015 36165
rect 40957 36125 40969 36159
rect 41003 36156 41015 36159
rect 41138 36156 41144 36168
rect 41003 36128 41144 36156
rect 41003 36125 41015 36128
rect 40957 36119 41015 36125
rect 41138 36116 41144 36128
rect 41196 36156 41202 36168
rect 41417 36159 41475 36165
rect 41417 36156 41429 36159
rect 41196 36128 41429 36156
rect 41196 36116 41202 36128
rect 41417 36125 41429 36128
rect 41463 36125 41475 36159
rect 42610 36156 42616 36168
rect 42571 36128 42616 36156
rect 41417 36119 41475 36125
rect 42610 36116 42616 36128
rect 42668 36116 42674 36168
rect 43625 36159 43683 36165
rect 43625 36125 43637 36159
rect 43671 36125 43683 36159
rect 44082 36156 44088 36168
rect 44043 36128 44088 36156
rect 43625 36119 43683 36125
rect 36648 36060 40172 36088
rect 40236 36060 41000 36088
rect 26384 36048 26390 36060
rect 26786 36020 26792 36032
rect 24044 35992 26792 36020
rect 21361 35983 21419 35989
rect 26786 35980 26792 35992
rect 26844 35980 26850 36032
rect 26881 36023 26939 36029
rect 26881 35989 26893 36023
rect 26927 36020 26939 36023
rect 28460 36020 28488 36060
rect 28626 36020 28632 36032
rect 26927 35992 28488 36020
rect 28587 35992 28632 36020
rect 26927 35989 26939 35992
rect 26881 35983 26939 35989
rect 28626 35980 28632 35992
rect 28684 35980 28690 36032
rect 29270 35980 29276 36032
rect 29328 36020 29334 36032
rect 32306 36020 32312 36032
rect 29328 35992 32312 36020
rect 29328 35980 29334 35992
rect 32306 35980 32312 35992
rect 32364 35980 32370 36032
rect 32416 36029 32444 36060
rect 32401 36023 32459 36029
rect 32401 35989 32413 36023
rect 32447 35989 32459 36023
rect 33134 36020 33140 36032
rect 33095 35992 33140 36020
rect 32401 35983 32459 35989
rect 33134 35980 33140 35992
rect 33192 35980 33198 36032
rect 33226 35980 33232 36032
rect 33284 36020 33290 36032
rect 35437 36023 35495 36029
rect 35437 36020 35449 36023
rect 33284 35992 35449 36020
rect 33284 35980 33290 35992
rect 35437 35989 35449 35992
rect 35483 36020 35495 36023
rect 35986 36020 35992 36032
rect 35483 35992 35992 36020
rect 35483 35989 35495 35992
rect 35437 35983 35495 35989
rect 35986 35980 35992 35992
rect 36044 35980 36050 36032
rect 36538 36020 36544 36032
rect 36499 35992 36544 36020
rect 36538 35980 36544 35992
rect 36596 35980 36602 36032
rect 38933 36023 38991 36029
rect 38933 35989 38945 36023
rect 38979 36020 38991 36023
rect 40034 36020 40040 36032
rect 38979 35992 40040 36020
rect 38979 35989 38991 35992
rect 38933 35983 38991 35989
rect 40034 35980 40040 35992
rect 40092 35980 40098 36032
rect 40236 36029 40264 36060
rect 40221 36023 40279 36029
rect 40221 35989 40233 36023
rect 40267 35989 40279 36023
rect 40972 36020 41000 36060
rect 41046 36048 41052 36100
rect 41104 36088 41110 36100
rect 43640 36088 43668 36119
rect 44082 36116 44088 36128
rect 44140 36116 44146 36168
rect 44358 36088 44364 36100
rect 41104 36060 43576 36088
rect 43640 36060 44364 36088
rect 41104 36048 41110 36060
rect 42058 36020 42064 36032
rect 40972 35992 42064 36020
rect 40221 35983 40279 35989
rect 42058 35980 42064 35992
rect 42116 35980 42122 36032
rect 43548 36020 43576 36060
rect 44358 36048 44364 36060
rect 44416 36088 44422 36100
rect 44634 36088 44640 36100
rect 44416 36060 44640 36088
rect 44416 36048 44422 36060
rect 44634 36048 44640 36060
rect 44692 36048 44698 36100
rect 45526 36088 45554 36196
rect 46477 36193 46489 36227
rect 46523 36224 46535 36227
rect 47210 36224 47216 36236
rect 46523 36196 47216 36224
rect 46523 36193 46535 36196
rect 46477 36187 46535 36193
rect 47210 36184 47216 36196
rect 47268 36224 47274 36236
rect 48056 36224 48084 36264
rect 48590 36252 48596 36264
rect 48648 36252 48654 36304
rect 49513 36295 49571 36301
rect 49513 36261 49525 36295
rect 49559 36261 49571 36295
rect 49513 36255 49571 36261
rect 50801 36295 50859 36301
rect 50801 36261 50813 36295
rect 50847 36292 50859 36295
rect 51258 36292 51264 36304
rect 50847 36264 51264 36292
rect 50847 36261 50859 36264
rect 50801 36255 50859 36261
rect 47268 36196 48084 36224
rect 48133 36227 48191 36233
rect 47268 36184 47274 36196
rect 48133 36193 48145 36227
rect 48179 36224 48191 36227
rect 49528 36224 49556 36255
rect 51258 36252 51264 36264
rect 51316 36252 51322 36304
rect 52181 36295 52239 36301
rect 52181 36261 52193 36295
rect 52227 36292 52239 36295
rect 53006 36292 53012 36304
rect 52227 36264 53012 36292
rect 52227 36261 52239 36264
rect 52181 36255 52239 36261
rect 53006 36252 53012 36264
rect 53064 36252 53070 36304
rect 53300 36224 53328 36332
rect 53374 36320 53380 36372
rect 53432 36360 53438 36372
rect 53469 36363 53527 36369
rect 53469 36360 53481 36363
rect 53432 36332 53481 36360
rect 53432 36320 53438 36332
rect 53469 36329 53481 36332
rect 53515 36329 53527 36363
rect 53469 36323 53527 36329
rect 54205 36363 54263 36369
rect 54205 36329 54217 36363
rect 54251 36360 54263 36363
rect 54294 36360 54300 36372
rect 54251 36332 54300 36360
rect 54251 36329 54263 36332
rect 54205 36323 54263 36329
rect 54294 36320 54300 36332
rect 54352 36320 54358 36372
rect 54754 36360 54760 36372
rect 54715 36332 54760 36360
rect 54754 36320 54760 36332
rect 54812 36320 54818 36372
rect 55861 36363 55919 36369
rect 55861 36329 55873 36363
rect 55907 36360 55919 36363
rect 56042 36360 56048 36372
rect 55907 36332 56048 36360
rect 55907 36329 55919 36332
rect 55861 36323 55919 36329
rect 56042 36320 56048 36332
rect 56100 36320 56106 36372
rect 56134 36320 56140 36372
rect 56192 36360 56198 36372
rect 58710 36360 58716 36372
rect 56192 36332 58716 36360
rect 56192 36320 56198 36332
rect 58710 36320 58716 36332
rect 58768 36320 58774 36372
rect 58802 36320 58808 36372
rect 58860 36360 58866 36372
rect 59633 36363 59691 36369
rect 59633 36360 59645 36363
rect 58860 36332 59645 36360
rect 58860 36320 58866 36332
rect 59633 36329 59645 36332
rect 59679 36329 59691 36363
rect 59633 36323 59691 36329
rect 59814 36320 59820 36372
rect 59872 36360 59878 36372
rect 61654 36360 61660 36372
rect 59872 36332 61660 36360
rect 59872 36320 59878 36332
rect 61654 36320 61660 36332
rect 61712 36320 61718 36372
rect 62482 36320 62488 36372
rect 62540 36360 62546 36372
rect 62669 36363 62727 36369
rect 62669 36360 62681 36363
rect 62540 36332 62681 36360
rect 62540 36320 62546 36332
rect 62669 36329 62681 36332
rect 62715 36329 62727 36363
rect 62669 36323 62727 36329
rect 64322 36320 64328 36372
rect 64380 36360 64386 36372
rect 64509 36363 64567 36369
rect 64509 36360 64521 36363
rect 64380 36332 64521 36360
rect 64380 36320 64386 36332
rect 64509 36329 64521 36332
rect 64555 36329 64567 36363
rect 64509 36323 64567 36329
rect 64782 36320 64788 36372
rect 64840 36360 64846 36372
rect 66254 36360 66260 36372
rect 64840 36332 66260 36360
rect 64840 36320 64846 36332
rect 66254 36320 66260 36332
rect 66312 36320 66318 36372
rect 67082 36360 67088 36372
rect 67043 36332 67088 36360
rect 67082 36320 67088 36332
rect 67140 36320 67146 36372
rect 68002 36320 68008 36372
rect 68060 36360 68066 36372
rect 68189 36363 68247 36369
rect 68189 36360 68201 36363
rect 68060 36332 68201 36360
rect 68060 36320 68066 36332
rect 68189 36329 68201 36332
rect 68235 36329 68247 36363
rect 68189 36323 68247 36329
rect 70394 36320 70400 36372
rect 70452 36360 70458 36372
rect 72326 36360 72332 36372
rect 70452 36332 70497 36360
rect 70780 36332 72332 36360
rect 70452 36320 70458 36332
rect 55122 36252 55128 36304
rect 55180 36292 55186 36304
rect 60829 36295 60887 36301
rect 55180 36264 60780 36292
rect 55180 36252 55186 36264
rect 48179 36196 49464 36224
rect 49528 36196 53052 36224
rect 53300 36196 59676 36224
rect 48179 36193 48191 36196
rect 48133 36187 48191 36193
rect 45925 36159 45983 36165
rect 45925 36125 45937 36159
rect 45971 36156 45983 36159
rect 46842 36156 46848 36168
rect 45971 36128 46848 36156
rect 45971 36125 45983 36128
rect 45925 36119 45983 36125
rect 46842 36116 46848 36128
rect 46900 36156 46906 36168
rect 46937 36159 46995 36165
rect 46937 36156 46949 36159
rect 46900 36128 46949 36156
rect 46900 36116 46906 36128
rect 46937 36125 46949 36128
rect 46983 36125 46995 36159
rect 48498 36156 48504 36168
rect 46937 36119 46995 36125
rect 47044 36128 48504 36156
rect 47044 36088 47072 36128
rect 48498 36116 48504 36128
rect 48556 36116 48562 36168
rect 48682 36116 48688 36168
rect 48740 36156 48746 36168
rect 49329 36159 49387 36165
rect 49329 36156 49341 36159
rect 48740 36128 49341 36156
rect 48740 36116 48746 36128
rect 49329 36125 49341 36128
rect 49375 36125 49387 36159
rect 49329 36119 49387 36125
rect 45526 36060 47072 36088
rect 48406 36048 48412 36100
rect 48464 36088 48470 36100
rect 48593 36091 48651 36097
rect 48593 36088 48605 36091
rect 48464 36060 48605 36088
rect 48464 36048 48470 36060
rect 48593 36057 48605 36060
rect 48639 36057 48651 36091
rect 48593 36051 48651 36057
rect 48777 36091 48835 36097
rect 48777 36057 48789 36091
rect 48823 36088 48835 36091
rect 49436 36088 49464 36196
rect 50614 36156 50620 36168
rect 50575 36128 50620 36156
rect 50614 36116 50620 36128
rect 50672 36116 50678 36168
rect 51997 36159 52055 36165
rect 51997 36125 52009 36159
rect 52043 36156 52055 36159
rect 52270 36156 52276 36168
rect 52043 36128 52276 36156
rect 52043 36125 52055 36128
rect 51997 36119 52055 36125
rect 52270 36116 52276 36128
rect 52328 36116 52334 36168
rect 53024 36152 53052 36196
rect 53098 36152 53104 36168
rect 53024 36124 53104 36152
rect 53098 36116 53104 36124
rect 53156 36116 53162 36168
rect 53653 36159 53711 36165
rect 53653 36125 53665 36159
rect 53699 36156 53711 36159
rect 54294 36156 54300 36168
rect 53699 36128 54300 36156
rect 53699 36125 53711 36128
rect 53653 36119 53711 36125
rect 54294 36116 54300 36128
rect 54352 36116 54358 36168
rect 57974 36156 57980 36168
rect 56244 36128 57284 36156
rect 57935 36128 57980 36156
rect 49694 36088 49700 36100
rect 48823 36060 49700 36088
rect 48823 36057 48835 36060
rect 48777 36051 48835 36057
rect 49694 36048 49700 36060
rect 49752 36088 49758 36100
rect 50246 36088 50252 36100
rect 49752 36060 50252 36088
rect 49752 36048 49758 36060
rect 50246 36048 50252 36060
rect 50304 36048 50310 36100
rect 52730 36088 52736 36100
rect 52691 36060 52736 36088
rect 52730 36048 52736 36060
rect 52788 36048 52794 36100
rect 52914 36088 52920 36100
rect 52875 36060 52920 36088
rect 52914 36048 52920 36060
rect 52972 36048 52978 36100
rect 44174 36020 44180 36032
rect 43548 35992 44180 36020
rect 44174 35980 44180 35992
rect 44232 35980 44238 36032
rect 45278 36020 45284 36032
rect 45239 35992 45284 36020
rect 45278 35980 45284 35992
rect 45336 35980 45342 36032
rect 47121 36023 47179 36029
rect 47121 35989 47133 36023
rect 47167 36020 47179 36023
rect 50706 36020 50712 36032
rect 47167 35992 50712 36020
rect 47167 35989 47179 35992
rect 47121 35983 47179 35989
rect 50706 35980 50712 35992
rect 50764 35980 50770 36032
rect 51534 36020 51540 36032
rect 51495 35992 51540 36020
rect 51534 35980 51540 35992
rect 51592 35980 51598 36032
rect 53006 35980 53012 36032
rect 53064 36020 53070 36032
rect 56244 36020 56272 36128
rect 56965 36091 57023 36097
rect 56965 36088 56977 36091
rect 56612 36060 56977 36088
rect 56612 36032 56640 36060
rect 56965 36057 56977 36060
rect 57011 36057 57023 36091
rect 57146 36088 57152 36100
rect 57107 36060 57152 36088
rect 56965 36051 57023 36057
rect 57146 36048 57152 36060
rect 57204 36048 57210 36100
rect 57256 36088 57284 36128
rect 57974 36116 57980 36128
rect 58032 36116 58038 36168
rect 58066 36088 58072 36100
rect 57256 36060 58072 36088
rect 58066 36048 58072 36060
rect 58124 36048 58130 36100
rect 58894 36088 58900 36100
rect 58855 36060 58900 36088
rect 58894 36048 58900 36060
rect 58952 36048 58958 36100
rect 59081 36091 59139 36097
rect 59081 36057 59093 36091
rect 59127 36088 59139 36091
rect 59262 36088 59268 36100
rect 59127 36060 59268 36088
rect 59127 36057 59139 36060
rect 59081 36051 59139 36057
rect 59262 36048 59268 36060
rect 59320 36048 59326 36100
rect 59648 36088 59676 36196
rect 59722 36184 59728 36236
rect 59780 36224 59786 36236
rect 60752 36224 60780 36264
rect 60829 36261 60841 36295
rect 60875 36292 60887 36295
rect 62574 36292 62580 36304
rect 60875 36264 62580 36292
rect 60875 36261 60887 36264
rect 60829 36255 60887 36261
rect 62574 36252 62580 36264
rect 62632 36252 62638 36304
rect 63310 36252 63316 36304
rect 63368 36292 63374 36304
rect 67818 36292 67824 36304
rect 63368 36264 67824 36292
rect 63368 36252 63374 36264
rect 67818 36252 67824 36264
rect 67876 36252 67882 36304
rect 69201 36295 69259 36301
rect 69201 36261 69213 36295
rect 69247 36292 69259 36295
rect 70780 36292 70808 36332
rect 72326 36320 72332 36332
rect 72384 36320 72390 36372
rect 72602 36360 72608 36372
rect 72563 36332 72608 36360
rect 72602 36320 72608 36332
rect 72660 36320 72666 36372
rect 74077 36363 74135 36369
rect 74077 36329 74089 36363
rect 74123 36360 74135 36363
rect 74442 36360 74448 36372
rect 74123 36332 74448 36360
rect 74123 36329 74135 36332
rect 74077 36323 74135 36329
rect 74442 36320 74448 36332
rect 74500 36320 74506 36372
rect 74721 36363 74779 36369
rect 74721 36329 74733 36363
rect 74767 36360 74779 36363
rect 75546 36360 75552 36372
rect 74767 36332 75552 36360
rect 74767 36329 74779 36332
rect 74721 36323 74779 36329
rect 75546 36320 75552 36332
rect 75604 36320 75610 36372
rect 76282 36360 76288 36372
rect 76243 36332 76288 36360
rect 76282 36320 76288 36332
rect 76340 36320 76346 36372
rect 79962 36360 79968 36372
rect 76392 36332 79968 36360
rect 69247 36264 70808 36292
rect 69247 36261 69259 36264
rect 69201 36255 69259 36261
rect 70854 36252 70860 36304
rect 70912 36292 70918 36304
rect 70949 36295 71007 36301
rect 70949 36292 70961 36295
rect 70912 36264 70961 36292
rect 70912 36252 70918 36264
rect 70949 36261 70961 36264
rect 70995 36261 71007 36295
rect 70949 36255 71007 36261
rect 71130 36252 71136 36304
rect 71188 36292 71194 36304
rect 76392 36292 76420 36332
rect 79962 36320 79968 36332
rect 80020 36320 80026 36372
rect 80146 36320 80152 36372
rect 80204 36360 80210 36372
rect 80241 36363 80299 36369
rect 80241 36360 80253 36363
rect 80204 36332 80253 36360
rect 80204 36320 80210 36332
rect 80241 36329 80253 36332
rect 80287 36329 80299 36363
rect 80241 36323 80299 36329
rect 80514 36320 80520 36372
rect 80572 36360 80578 36372
rect 89254 36360 89260 36372
rect 80572 36332 89260 36360
rect 80572 36320 80578 36332
rect 89254 36320 89260 36332
rect 89312 36320 89318 36372
rect 90726 36360 90732 36372
rect 90687 36332 90732 36360
rect 90726 36320 90732 36332
rect 90784 36320 90790 36372
rect 93854 36320 93860 36372
rect 93912 36360 93918 36372
rect 93949 36363 94007 36369
rect 93949 36360 93961 36363
rect 93912 36332 93961 36360
rect 93912 36320 93918 36332
rect 93949 36329 93961 36332
rect 93995 36329 94007 36363
rect 93949 36323 94007 36329
rect 102870 36320 102876 36372
rect 102928 36360 102934 36372
rect 102965 36363 103023 36369
rect 102965 36360 102977 36363
rect 102928 36332 102977 36360
rect 102928 36320 102934 36332
rect 102965 36329 102977 36332
rect 103011 36360 103023 36363
rect 103054 36360 103060 36372
rect 103011 36332 103060 36360
rect 103011 36329 103023 36332
rect 102965 36323 103023 36329
rect 103054 36320 103060 36332
rect 103112 36320 103118 36372
rect 103422 36360 103428 36372
rect 103383 36332 103428 36360
rect 103422 36320 103428 36332
rect 103480 36320 103486 36372
rect 104894 36320 104900 36372
rect 104952 36360 104958 36372
rect 104989 36363 105047 36369
rect 104989 36360 105001 36363
rect 104952 36332 105001 36360
rect 104952 36320 104958 36332
rect 104989 36329 105001 36332
rect 105035 36329 105047 36363
rect 106366 36360 106372 36372
rect 106327 36332 106372 36360
rect 104989 36323 105047 36329
rect 106366 36320 106372 36332
rect 106424 36320 106430 36372
rect 106550 36320 106556 36372
rect 106608 36360 106614 36372
rect 107105 36363 107163 36369
rect 107105 36360 107117 36363
rect 106608 36332 107117 36360
rect 106608 36320 106614 36332
rect 107105 36329 107117 36332
rect 107151 36360 107163 36363
rect 107562 36360 107568 36372
rect 107151 36332 107568 36360
rect 107151 36329 107163 36332
rect 107105 36323 107163 36329
rect 107562 36320 107568 36332
rect 107620 36320 107626 36372
rect 107657 36363 107715 36369
rect 107657 36329 107669 36363
rect 107703 36360 107715 36363
rect 107746 36360 107752 36372
rect 107703 36332 107752 36360
rect 107703 36329 107715 36332
rect 107657 36323 107715 36329
rect 107746 36320 107752 36332
rect 107804 36320 107810 36372
rect 110690 36320 110696 36372
rect 110748 36360 110754 36372
rect 110877 36363 110935 36369
rect 110877 36360 110889 36363
rect 110748 36332 110889 36360
rect 110748 36320 110754 36332
rect 110877 36329 110889 36332
rect 110923 36329 110935 36363
rect 110877 36323 110935 36329
rect 112346 36320 112352 36372
rect 112404 36360 112410 36372
rect 115293 36363 115351 36369
rect 115293 36360 115305 36363
rect 112404 36332 115305 36360
rect 112404 36320 112410 36332
rect 115293 36329 115305 36332
rect 115339 36360 115351 36363
rect 115474 36360 115480 36372
rect 115339 36332 115480 36360
rect 115339 36329 115351 36332
rect 115293 36323 115351 36329
rect 115474 36320 115480 36332
rect 115532 36320 115538 36372
rect 117682 36320 117688 36372
rect 117740 36360 117746 36372
rect 117869 36363 117927 36369
rect 117869 36360 117881 36363
rect 117740 36332 117881 36360
rect 117740 36320 117746 36332
rect 117869 36329 117881 36332
rect 117915 36329 117927 36363
rect 117869 36323 117927 36329
rect 119706 36320 119712 36372
rect 119764 36360 119770 36372
rect 123202 36360 123208 36372
rect 119764 36332 123208 36360
rect 119764 36320 119770 36332
rect 123202 36320 123208 36332
rect 123260 36320 123266 36372
rect 123294 36320 123300 36372
rect 123352 36360 123358 36372
rect 135898 36360 135904 36372
rect 123352 36332 135904 36360
rect 123352 36320 123358 36332
rect 135898 36320 135904 36332
rect 135956 36320 135962 36372
rect 136082 36360 136088 36372
rect 136043 36332 136088 36360
rect 136082 36320 136088 36332
rect 136140 36320 136146 36372
rect 138014 36360 138020 36372
rect 137975 36332 138020 36360
rect 138014 36320 138020 36332
rect 138072 36320 138078 36372
rect 143534 36320 143540 36372
rect 143592 36360 143598 36372
rect 143629 36363 143687 36369
rect 143629 36360 143641 36363
rect 143592 36332 143641 36360
rect 143592 36320 143598 36332
rect 143629 36329 143641 36332
rect 143675 36329 143687 36363
rect 143629 36323 143687 36329
rect 71188 36264 76420 36292
rect 78677 36295 78735 36301
rect 71188 36252 71194 36264
rect 78677 36261 78689 36295
rect 78723 36292 78735 36295
rect 78723 36264 83964 36292
rect 78723 36261 78735 36264
rect 78677 36255 78735 36261
rect 64598 36224 64604 36236
rect 59780 36196 60320 36224
rect 60752 36196 64604 36224
rect 59780 36184 59786 36196
rect 59817 36159 59875 36165
rect 59817 36125 59829 36159
rect 59863 36156 59875 36159
rect 59906 36156 59912 36168
rect 59863 36128 59912 36156
rect 59863 36125 59875 36128
rect 59817 36119 59875 36125
rect 59906 36116 59912 36128
rect 59964 36116 59970 36168
rect 60292 36156 60320 36196
rect 64598 36184 64604 36196
rect 64656 36184 64662 36236
rect 67637 36227 67695 36233
rect 67637 36193 67649 36227
rect 67683 36224 67695 36227
rect 67726 36224 67732 36236
rect 67683 36196 67732 36224
rect 67683 36193 67695 36196
rect 67637 36187 67695 36193
rect 67726 36184 67732 36196
rect 67784 36224 67790 36236
rect 67784 36196 70256 36224
rect 67784 36184 67790 36196
rect 60366 36156 60372 36168
rect 60279 36128 60372 36156
rect 60366 36116 60372 36128
rect 60424 36156 60430 36168
rect 60645 36159 60703 36165
rect 60645 36156 60657 36159
rect 60424 36152 60504 36156
rect 60568 36152 60657 36156
rect 60424 36128 60657 36152
rect 60424 36116 60430 36128
rect 60476 36124 60596 36128
rect 60645 36125 60657 36128
rect 60691 36125 60703 36159
rect 61378 36156 61384 36168
rect 61339 36128 61384 36156
rect 60645 36119 60703 36125
rect 61378 36116 61384 36128
rect 61436 36116 61442 36168
rect 62574 36156 62580 36168
rect 61580 36128 62580 36156
rect 61580 36088 61608 36128
rect 62574 36116 62580 36128
rect 62632 36116 62638 36168
rect 62850 36156 62856 36168
rect 62811 36128 62856 36156
rect 62850 36116 62856 36128
rect 62908 36116 62914 36168
rect 64690 36156 64696 36168
rect 64651 36128 64696 36156
rect 64690 36116 64696 36128
rect 64748 36116 64754 36168
rect 65334 36116 65340 36168
rect 65392 36156 65398 36168
rect 68186 36156 68192 36168
rect 65392 36128 68192 36156
rect 65392 36116 65398 36128
rect 68186 36116 68192 36128
rect 68244 36116 68250 36168
rect 68370 36156 68376 36168
rect 68331 36128 68376 36156
rect 68370 36116 68376 36128
rect 68428 36116 68434 36168
rect 68922 36116 68928 36168
rect 68980 36156 68986 36168
rect 69017 36159 69075 36165
rect 69017 36156 69029 36159
rect 68980 36128 69029 36156
rect 68980 36116 68986 36128
rect 69017 36125 69029 36128
rect 69063 36156 69075 36159
rect 69661 36159 69719 36165
rect 69661 36156 69673 36159
rect 69063 36128 69673 36156
rect 69063 36125 69075 36128
rect 69017 36119 69075 36125
rect 69661 36125 69673 36128
rect 69707 36125 69719 36159
rect 70228 36156 70256 36196
rect 71038 36184 71044 36236
rect 71096 36224 71102 36236
rect 80606 36224 80612 36236
rect 71096 36196 80612 36224
rect 71096 36184 71102 36196
rect 80606 36184 80612 36196
rect 80664 36184 80670 36236
rect 81342 36224 81348 36236
rect 81303 36196 81348 36224
rect 81342 36184 81348 36196
rect 81400 36184 81406 36236
rect 82449 36227 82507 36233
rect 82449 36224 82461 36227
rect 81452 36196 82461 36224
rect 70228 36128 74120 36156
rect 69661 36119 69719 36125
rect 59648 36060 61608 36088
rect 61654 36048 61660 36100
rect 61712 36088 61718 36100
rect 61749 36091 61807 36097
rect 61749 36088 61761 36091
rect 61712 36060 61761 36088
rect 61712 36048 61718 36060
rect 61749 36057 61761 36060
rect 61795 36088 61807 36091
rect 62022 36088 62028 36100
rect 61795 36060 62028 36088
rect 61795 36057 61807 36060
rect 61749 36051 61807 36057
rect 62022 36048 62028 36060
rect 62080 36048 62086 36100
rect 63678 36088 63684 36100
rect 63639 36060 63684 36088
rect 63678 36048 63684 36060
rect 63736 36048 63742 36100
rect 63862 36088 63868 36100
rect 63823 36060 63868 36088
rect 63862 36048 63868 36060
rect 63920 36048 63926 36100
rect 65426 36088 65432 36100
rect 63972 36060 65432 36088
rect 53064 35992 56272 36020
rect 56413 36023 56471 36029
rect 53064 35980 53070 35992
rect 56413 35989 56425 36023
rect 56459 36020 56471 36023
rect 56594 36020 56600 36032
rect 56459 35992 56600 36020
rect 56459 35989 56471 35992
rect 56413 35983 56471 35989
rect 56594 35980 56600 35992
rect 56652 35980 56658 36032
rect 58161 36023 58219 36029
rect 58161 35989 58173 36023
rect 58207 36020 58219 36023
rect 63972 36020 64000 36060
rect 65426 36048 65432 36060
rect 65484 36048 65490 36100
rect 65889 36091 65947 36097
rect 65889 36057 65901 36091
rect 65935 36057 65947 36091
rect 66070 36088 66076 36100
rect 66031 36060 66076 36088
rect 65889 36051 65947 36057
rect 58207 35992 64000 36020
rect 58207 35989 58219 35992
rect 58161 35983 58219 35989
rect 64782 35980 64788 36032
rect 64840 36020 64846 36032
rect 65153 36023 65211 36029
rect 65153 36020 65165 36023
rect 64840 35992 65165 36020
rect 64840 35980 64846 35992
rect 65153 35989 65165 35992
rect 65199 36020 65211 36023
rect 65904 36020 65932 36051
rect 66070 36048 66076 36060
rect 66128 36048 66134 36100
rect 73982 36088 73988 36100
rect 70366 36060 73988 36088
rect 65199 35992 65932 36020
rect 65199 35989 65211 35992
rect 65153 35983 65211 35989
rect 66438 35980 66444 36032
rect 66496 36020 66502 36032
rect 70366 36020 70394 36060
rect 73982 36048 73988 36060
rect 74040 36048 74046 36100
rect 74092 36088 74120 36128
rect 74442 36116 74448 36168
rect 74500 36156 74506 36168
rect 74537 36159 74595 36165
rect 74537 36156 74549 36159
rect 74500 36128 74549 36156
rect 74500 36116 74506 36128
rect 74537 36125 74549 36128
rect 74583 36125 74595 36159
rect 74537 36119 74595 36125
rect 74626 36116 74632 36168
rect 74684 36156 74690 36168
rect 76098 36156 76104 36168
rect 74684 36128 75592 36156
rect 76059 36128 76104 36156
rect 74684 36116 74690 36128
rect 75086 36088 75092 36100
rect 74092 36060 75092 36088
rect 75086 36048 75092 36060
rect 75144 36048 75150 36100
rect 75564 36088 75592 36128
rect 76098 36116 76104 36128
rect 76156 36116 76162 36168
rect 77294 36156 77300 36168
rect 77255 36128 77300 36156
rect 77294 36116 77300 36128
rect 77352 36116 77358 36168
rect 80054 36116 80060 36168
rect 80112 36156 80118 36168
rect 80112 36128 80157 36156
rect 80112 36116 80118 36128
rect 80422 36116 80428 36168
rect 80480 36156 80486 36168
rect 81452 36156 81480 36196
rect 82449 36193 82461 36196
rect 82495 36193 82507 36227
rect 82449 36187 82507 36193
rect 82814 36184 82820 36236
rect 82872 36224 82878 36236
rect 83642 36224 83648 36236
rect 82872 36196 83648 36224
rect 82872 36184 82878 36196
rect 83642 36184 83648 36196
rect 83700 36184 83706 36236
rect 83936 36224 83964 36264
rect 86402 36252 86408 36304
rect 86460 36292 86466 36304
rect 119154 36292 119160 36304
rect 86460 36264 119160 36292
rect 86460 36252 86466 36264
rect 119154 36252 119160 36264
rect 119212 36252 119218 36304
rect 120810 36252 120816 36304
rect 120868 36292 120874 36304
rect 121089 36295 121147 36301
rect 121089 36292 121101 36295
rect 120868 36264 121101 36292
rect 120868 36252 120874 36264
rect 121089 36261 121101 36264
rect 121135 36292 121147 36295
rect 126422 36292 126428 36304
rect 121135 36264 124352 36292
rect 126383 36264 126428 36292
rect 121135 36261 121147 36264
rect 121089 36255 121147 36261
rect 105817 36227 105875 36233
rect 83936 36196 105768 36224
rect 81618 36156 81624 36168
rect 80480 36128 81480 36156
rect 81579 36128 81624 36156
rect 80480 36116 80486 36128
rect 81618 36116 81624 36128
rect 81676 36116 81682 36168
rect 81710 36116 81716 36168
rect 81768 36156 81774 36168
rect 82354 36156 82360 36168
rect 81768 36128 82360 36156
rect 81768 36116 81774 36128
rect 82354 36116 82360 36128
rect 82412 36156 82418 36168
rect 87598 36156 87604 36168
rect 82412 36128 87604 36156
rect 82412 36116 82418 36128
rect 87598 36116 87604 36128
rect 87656 36116 87662 36168
rect 95050 36156 95056 36168
rect 89686 36128 95056 36156
rect 77941 36091 77999 36097
rect 77941 36088 77953 36091
rect 75564 36060 77953 36088
rect 77941 36057 77953 36060
rect 77987 36088 77999 36091
rect 78490 36088 78496 36100
rect 77987 36060 78496 36088
rect 77987 36057 77999 36060
rect 77941 36051 77999 36057
rect 78490 36048 78496 36060
rect 78548 36048 78554 36100
rect 89686 36088 89714 36128
rect 95050 36116 95056 36128
rect 95108 36116 95114 36168
rect 99374 36156 99380 36168
rect 95160 36128 99380 36156
rect 78600 36060 89714 36088
rect 66496 35992 70394 36020
rect 66496 35980 66502 35992
rect 75178 35980 75184 36032
rect 75236 36020 75242 36032
rect 75236 35992 75281 36020
rect 75236 35980 75242 35992
rect 75730 35980 75736 36032
rect 75788 36020 75794 36032
rect 78600 36020 78628 36060
rect 92382 36048 92388 36100
rect 92440 36088 92446 36100
rect 95160 36088 95188 36128
rect 99374 36116 99380 36128
rect 99432 36116 99438 36168
rect 99466 36116 99472 36168
rect 99524 36156 99530 36168
rect 105630 36156 105636 36168
rect 99524 36128 105636 36156
rect 99524 36116 99530 36128
rect 105630 36116 105636 36128
rect 105688 36116 105694 36168
rect 105740 36156 105768 36196
rect 105817 36193 105829 36227
rect 105863 36224 105875 36227
rect 106458 36224 106464 36236
rect 105863 36196 106464 36224
rect 105863 36193 105875 36196
rect 105817 36187 105875 36193
rect 106458 36184 106464 36196
rect 106516 36184 106522 36236
rect 108298 36184 108304 36236
rect 108356 36224 108362 36236
rect 116302 36224 116308 36236
rect 108356 36196 116308 36224
rect 108356 36184 108362 36196
rect 116302 36184 116308 36196
rect 116360 36184 116366 36236
rect 120902 36184 120908 36236
rect 120960 36224 120966 36236
rect 124214 36224 124220 36236
rect 120960 36196 124220 36224
rect 120960 36184 120966 36196
rect 124214 36184 124220 36196
rect 124272 36184 124278 36236
rect 124324 36224 124352 36264
rect 126422 36252 126428 36264
rect 126480 36252 126486 36304
rect 126514 36252 126520 36304
rect 126572 36292 126578 36304
rect 132034 36292 132040 36304
rect 126572 36264 132040 36292
rect 126572 36252 126578 36264
rect 132034 36252 132040 36264
rect 132092 36252 132098 36304
rect 132126 36252 132132 36304
rect 132184 36292 132190 36304
rect 137278 36292 137284 36304
rect 132184 36264 137284 36292
rect 132184 36252 132190 36264
rect 137278 36252 137284 36264
rect 137336 36252 137342 36304
rect 139486 36224 139492 36236
rect 124324 36196 139492 36224
rect 139486 36184 139492 36196
rect 139544 36184 139550 36236
rect 112346 36156 112352 36168
rect 105740 36128 112352 36156
rect 112346 36116 112352 36128
rect 112404 36116 112410 36168
rect 112530 36116 112536 36168
rect 112588 36156 112594 36168
rect 143626 36156 143632 36168
rect 112588 36128 143632 36156
rect 112588 36116 112594 36128
rect 143626 36116 143632 36128
rect 143684 36116 143690 36168
rect 92440 36060 95188 36088
rect 92440 36048 92446 36060
rect 95234 36048 95240 36100
rect 95292 36088 95298 36100
rect 95421 36091 95479 36097
rect 95421 36088 95433 36091
rect 95292 36060 95433 36088
rect 95292 36048 95298 36060
rect 95421 36057 95433 36060
rect 95467 36088 95479 36091
rect 98454 36088 98460 36100
rect 95467 36060 98460 36088
rect 95467 36057 95479 36060
rect 95421 36051 95479 36057
rect 98454 36048 98460 36060
rect 98512 36048 98518 36100
rect 98638 36048 98644 36100
rect 98696 36088 98702 36100
rect 146294 36088 146300 36100
rect 98696 36060 146300 36088
rect 98696 36048 98702 36060
rect 146294 36048 146300 36060
rect 146352 36088 146358 36100
rect 147306 36088 147312 36100
rect 146352 36060 147312 36088
rect 146352 36048 146358 36060
rect 147306 36048 147312 36060
rect 147364 36048 147370 36100
rect 75788 35992 78628 36020
rect 75788 35980 75794 35992
rect 78950 35980 78956 36032
rect 79008 36020 79014 36032
rect 79134 36020 79140 36032
rect 79008 35992 79140 36020
rect 79008 35980 79014 35992
rect 79134 35980 79140 35992
rect 79192 35980 79198 36032
rect 81529 36023 81587 36029
rect 81529 35989 81541 36023
rect 81575 36020 81587 36023
rect 81710 36020 81716 36032
rect 81575 35992 81716 36020
rect 81575 35989 81587 35992
rect 81529 35983 81587 35989
rect 81710 35980 81716 35992
rect 81768 35980 81774 36032
rect 81986 36020 81992 36032
rect 81947 35992 81992 36020
rect 81986 35980 81992 35992
rect 82044 35980 82050 36032
rect 83090 36020 83096 36032
rect 83051 35992 83096 36020
rect 83090 35980 83096 35992
rect 83148 35980 83154 36032
rect 83642 36020 83648 36032
rect 83603 35992 83648 36020
rect 83642 35980 83648 35992
rect 83700 35980 83706 36032
rect 83734 35980 83740 36032
rect 83792 36020 83798 36032
rect 84105 36023 84163 36029
rect 84105 36020 84117 36023
rect 83792 35992 84117 36020
rect 83792 35980 83798 35992
rect 84105 35989 84117 35992
rect 84151 35989 84163 36023
rect 84105 35983 84163 35989
rect 84194 35980 84200 36032
rect 84252 36020 84258 36032
rect 84746 36020 84752 36032
rect 84252 35992 84752 36020
rect 84252 35980 84258 35992
rect 84746 35980 84752 35992
rect 84804 35980 84810 36032
rect 85393 36023 85451 36029
rect 85393 35989 85405 36023
rect 85439 36020 85451 36023
rect 85482 36020 85488 36032
rect 85439 35992 85488 36020
rect 85439 35989 85451 35992
rect 85393 35983 85451 35989
rect 85482 35980 85488 35992
rect 85540 36020 85546 36032
rect 86405 36023 86463 36029
rect 86405 36020 86417 36023
rect 85540 35992 86417 36020
rect 85540 35980 85546 35992
rect 86405 35989 86417 35992
rect 86451 35989 86463 36023
rect 89070 36020 89076 36032
rect 89031 35992 89076 36020
rect 86405 35983 86463 35989
rect 89070 35980 89076 35992
rect 89128 35980 89134 36032
rect 89622 36020 89628 36032
rect 89583 35992 89628 36020
rect 89622 35980 89628 35992
rect 89680 35980 89686 36032
rect 89714 35980 89720 36032
rect 89772 36020 89778 36032
rect 90177 36023 90235 36029
rect 90177 36020 90189 36023
rect 89772 35992 90189 36020
rect 89772 35980 89778 35992
rect 90177 35989 90189 35992
rect 90223 36020 90235 36023
rect 90358 36020 90364 36032
rect 90223 35992 90364 36020
rect 90223 35989 90235 35992
rect 90177 35983 90235 35989
rect 90358 35980 90364 35992
rect 90416 35980 90422 36032
rect 92842 36020 92848 36032
rect 92803 35992 92848 36020
rect 92842 35980 92848 35992
rect 92900 35980 92906 36032
rect 94314 35980 94320 36032
rect 94372 36020 94378 36032
rect 94685 36023 94743 36029
rect 94685 36020 94697 36023
rect 94372 35992 94697 36020
rect 94372 35980 94378 35992
rect 94685 35989 94697 35992
rect 94731 35989 94743 36023
rect 95878 36020 95884 36032
rect 95839 35992 95884 36020
rect 94685 35983 94743 35989
rect 95878 35980 95884 35992
rect 95936 35980 95942 36032
rect 97810 36020 97816 36032
rect 97771 35992 97816 36020
rect 97810 35980 97816 35992
rect 97868 35980 97874 36032
rect 98362 36020 98368 36032
rect 98323 35992 98368 36020
rect 98362 35980 98368 35992
rect 98420 35980 98426 36032
rect 99374 35980 99380 36032
rect 99432 36020 99438 36032
rect 100570 36020 100576 36032
rect 99432 35992 100576 36020
rect 99432 35980 99438 35992
rect 100570 35980 100576 35992
rect 100628 35980 100634 36032
rect 105814 35980 105820 36032
rect 105872 36020 105878 36032
rect 110230 36020 110236 36032
rect 105872 35992 110236 36020
rect 105872 35980 105878 35992
rect 110230 35980 110236 35992
rect 110288 35980 110294 36032
rect 112162 36020 112168 36032
rect 112123 35992 112168 36020
rect 112162 35980 112168 35992
rect 112220 35980 112226 36032
rect 112714 36020 112720 36032
rect 112675 35992 112720 36020
rect 112714 35980 112720 35992
rect 112772 35980 112778 36032
rect 113450 36020 113456 36032
rect 113411 35992 113456 36020
rect 113450 35980 113456 35992
rect 113508 35980 113514 36032
rect 114189 36023 114247 36029
rect 114189 35989 114201 36023
rect 114235 36020 114247 36023
rect 114646 36020 114652 36032
rect 114235 35992 114652 36020
rect 114235 35989 114247 35992
rect 114189 35983 114247 35989
rect 114646 35980 114652 35992
rect 114704 35980 114710 36032
rect 114741 36023 114799 36029
rect 114741 35989 114753 36023
rect 114787 36020 114799 36023
rect 114922 36020 114928 36032
rect 114787 35992 114928 36020
rect 114787 35989 114799 35992
rect 114741 35983 114799 35989
rect 114922 35980 114928 35992
rect 114980 35980 114986 36032
rect 116946 35980 116952 36032
rect 117004 36020 117010 36032
rect 120902 36020 120908 36032
rect 117004 35992 120908 36020
rect 117004 35980 117010 35992
rect 120902 35980 120908 35992
rect 120960 35980 120966 36032
rect 121546 36020 121552 36032
rect 121507 35992 121552 36020
rect 121546 35980 121552 35992
rect 121604 35980 121610 36032
rect 123110 36020 123116 36032
rect 123071 35992 123116 36020
rect 123110 35980 123116 35992
rect 123168 35980 123174 36032
rect 123202 35980 123208 36032
rect 123260 36020 123266 36032
rect 130470 36020 130476 36032
rect 123260 35992 130476 36020
rect 123260 35980 123266 35992
rect 130470 35980 130476 35992
rect 130528 35980 130534 36032
rect 130930 35980 130936 36032
rect 130988 36020 130994 36032
rect 137646 36020 137652 36032
rect 130988 35992 137652 36020
rect 130988 35980 130994 35992
rect 137646 35980 137652 35992
rect 137704 35980 137710 36032
rect 1104 35930 148856 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 81014 35930
rect 81066 35878 81078 35930
rect 81130 35878 81142 35930
rect 81194 35878 81206 35930
rect 81258 35878 81270 35930
rect 81322 35878 111734 35930
rect 111786 35878 111798 35930
rect 111850 35878 111862 35930
rect 111914 35878 111926 35930
rect 111978 35878 111990 35930
rect 112042 35878 142454 35930
rect 142506 35878 142518 35930
rect 142570 35878 142582 35930
rect 142634 35878 142646 35930
rect 142698 35878 142710 35930
rect 142762 35878 148856 35930
rect 1104 35856 148856 35878
rect 19889 35819 19947 35825
rect 19889 35785 19901 35819
rect 19935 35816 19947 35819
rect 19978 35816 19984 35828
rect 19935 35788 19984 35816
rect 19935 35785 19947 35788
rect 19889 35779 19947 35785
rect 19978 35776 19984 35788
rect 20036 35776 20042 35828
rect 21082 35816 21088 35828
rect 21043 35788 21088 35816
rect 21082 35776 21088 35788
rect 21140 35776 21146 35828
rect 25130 35776 25136 35828
rect 25188 35816 25194 35828
rect 25225 35819 25283 35825
rect 25225 35816 25237 35819
rect 25188 35788 25237 35816
rect 25188 35776 25194 35788
rect 25225 35785 25237 35788
rect 25271 35785 25283 35819
rect 26602 35816 26608 35828
rect 26563 35788 26608 35816
rect 25225 35779 25283 35785
rect 26602 35776 26608 35788
rect 26660 35776 26666 35828
rect 28534 35816 28540 35828
rect 28495 35788 28540 35816
rect 28534 35776 28540 35788
rect 28592 35776 28598 35828
rect 28626 35776 28632 35828
rect 28684 35816 28690 35828
rect 29181 35819 29239 35825
rect 29181 35816 29193 35819
rect 28684 35788 29193 35816
rect 28684 35776 28690 35788
rect 29181 35785 29193 35788
rect 29227 35816 29239 35819
rect 29270 35816 29276 35828
rect 29227 35788 29276 35816
rect 29227 35785 29239 35788
rect 29181 35779 29239 35785
rect 29270 35776 29276 35788
rect 29328 35776 29334 35828
rect 31757 35819 31815 35825
rect 31757 35785 31769 35819
rect 31803 35816 31815 35819
rect 31938 35816 31944 35828
rect 31803 35788 31944 35816
rect 31803 35785 31815 35788
rect 31757 35779 31815 35785
rect 31938 35776 31944 35788
rect 31996 35776 32002 35828
rect 35253 35819 35311 35825
rect 35253 35785 35265 35819
rect 35299 35816 35311 35819
rect 36357 35819 36415 35825
rect 36357 35816 36369 35819
rect 35299 35788 36369 35816
rect 35299 35785 35311 35788
rect 35253 35779 35311 35785
rect 36357 35785 36369 35788
rect 36403 35816 36415 35819
rect 37458 35816 37464 35828
rect 36403 35788 37464 35816
rect 36403 35785 36415 35788
rect 36357 35779 36415 35785
rect 37458 35776 37464 35788
rect 37516 35776 37522 35828
rect 37642 35816 37648 35828
rect 37603 35788 37648 35816
rect 37642 35776 37648 35788
rect 37700 35776 37706 35828
rect 38654 35816 38660 35828
rect 38615 35788 38660 35816
rect 38654 35776 38660 35788
rect 38712 35776 38718 35828
rect 39301 35819 39359 35825
rect 39301 35785 39313 35819
rect 39347 35816 39359 35819
rect 39390 35816 39396 35828
rect 39347 35788 39396 35816
rect 39347 35785 39359 35788
rect 39301 35779 39359 35785
rect 39390 35776 39396 35788
rect 39448 35776 39454 35828
rect 41230 35776 41236 35828
rect 41288 35816 41294 35828
rect 42518 35816 42524 35828
rect 41288 35788 42524 35816
rect 41288 35776 41294 35788
rect 42518 35776 42524 35788
rect 42576 35776 42582 35828
rect 42610 35776 42616 35828
rect 42668 35816 42674 35828
rect 42705 35819 42763 35825
rect 42705 35816 42717 35819
rect 42668 35788 42717 35816
rect 42668 35776 42674 35788
rect 42705 35785 42717 35788
rect 42751 35785 42763 35819
rect 42705 35779 42763 35785
rect 43162 35776 43168 35828
rect 43220 35816 43226 35828
rect 43993 35819 44051 35825
rect 43993 35816 44005 35819
rect 43220 35788 44005 35816
rect 43220 35776 43226 35788
rect 43993 35785 44005 35788
rect 44039 35816 44051 35819
rect 44082 35816 44088 35828
rect 44039 35788 44088 35816
rect 44039 35785 44051 35788
rect 43993 35779 44051 35785
rect 44082 35776 44088 35788
rect 44140 35776 44146 35828
rect 45002 35776 45008 35828
rect 45060 35816 45066 35828
rect 45097 35819 45155 35825
rect 45097 35816 45109 35819
rect 45060 35788 45109 35816
rect 45060 35776 45066 35788
rect 45097 35785 45109 35788
rect 45143 35785 45155 35819
rect 45097 35779 45155 35785
rect 46109 35819 46167 35825
rect 46109 35785 46121 35819
rect 46155 35816 46167 35819
rect 46290 35816 46296 35828
rect 46155 35788 46296 35816
rect 46155 35785 46167 35788
rect 46109 35779 46167 35785
rect 46290 35776 46296 35788
rect 46348 35776 46354 35828
rect 46661 35819 46719 35825
rect 46661 35785 46673 35819
rect 46707 35816 46719 35819
rect 46934 35816 46940 35828
rect 46707 35788 46940 35816
rect 46707 35785 46719 35788
rect 46661 35779 46719 35785
rect 46934 35776 46940 35788
rect 46992 35776 46998 35828
rect 48682 35776 48688 35828
rect 48740 35816 48746 35828
rect 49145 35819 49203 35825
rect 49145 35816 49157 35819
rect 48740 35788 49157 35816
rect 48740 35776 48746 35788
rect 49145 35785 49157 35788
rect 49191 35785 49203 35819
rect 49145 35779 49203 35785
rect 50525 35819 50583 35825
rect 50525 35785 50537 35819
rect 50571 35816 50583 35819
rect 50614 35816 50620 35828
rect 50571 35788 50620 35816
rect 50571 35785 50583 35788
rect 50525 35779 50583 35785
rect 50614 35776 50620 35788
rect 50672 35776 50678 35828
rect 51261 35819 51319 35825
rect 51261 35785 51273 35819
rect 51307 35816 51319 35819
rect 51718 35816 51724 35828
rect 51307 35788 51724 35816
rect 51307 35785 51319 35788
rect 51261 35779 51319 35785
rect 51718 35776 51724 35788
rect 51776 35776 51782 35828
rect 52270 35816 52276 35828
rect 52231 35788 52276 35816
rect 52270 35776 52276 35788
rect 52328 35776 52334 35828
rect 54938 35776 54944 35828
rect 54996 35816 55002 35828
rect 55033 35819 55091 35825
rect 55033 35816 55045 35819
rect 54996 35788 55045 35816
rect 54996 35776 55002 35788
rect 55033 35785 55045 35788
rect 55079 35785 55091 35819
rect 55033 35779 55091 35785
rect 57517 35819 57575 35825
rect 57517 35785 57529 35819
rect 57563 35816 57575 35819
rect 57974 35816 57980 35828
rect 57563 35788 57980 35816
rect 57563 35785 57575 35788
rect 57517 35779 57575 35785
rect 57974 35776 57980 35788
rect 58032 35776 58038 35828
rect 58161 35819 58219 35825
rect 58161 35785 58173 35819
rect 58207 35816 58219 35819
rect 58618 35816 58624 35828
rect 58207 35788 58624 35816
rect 58207 35785 58219 35788
rect 58161 35779 58219 35785
rect 58618 35776 58624 35788
rect 58676 35776 58682 35828
rect 59909 35819 59967 35825
rect 59909 35785 59921 35819
rect 59955 35816 59967 35819
rect 60090 35816 60096 35828
rect 59955 35788 60096 35816
rect 59955 35785 59967 35788
rect 59909 35779 59967 35785
rect 60090 35776 60096 35788
rect 60148 35776 60154 35828
rect 60366 35816 60372 35828
rect 60327 35788 60372 35816
rect 60366 35776 60372 35788
rect 60424 35776 60430 35828
rect 61013 35819 61071 35825
rect 61013 35785 61025 35819
rect 61059 35816 61071 35819
rect 61286 35816 61292 35828
rect 61059 35788 61292 35816
rect 61059 35785 61071 35788
rect 61013 35779 61071 35785
rect 61286 35776 61292 35788
rect 61344 35776 61350 35828
rect 62669 35819 62727 35825
rect 62669 35785 62681 35819
rect 62715 35816 62727 35819
rect 63402 35816 63408 35828
rect 62715 35788 63408 35816
rect 62715 35785 62727 35788
rect 62669 35779 62727 35785
rect 63402 35776 63408 35788
rect 63460 35776 63466 35828
rect 64325 35819 64383 35825
rect 64325 35785 64337 35819
rect 64371 35816 64383 35819
rect 64414 35816 64420 35828
rect 64371 35788 64420 35816
rect 64371 35785 64383 35788
rect 64325 35779 64383 35785
rect 64414 35776 64420 35788
rect 64472 35776 64478 35828
rect 64690 35776 64696 35828
rect 64748 35816 64754 35828
rect 64877 35819 64935 35825
rect 64877 35816 64889 35819
rect 64748 35788 64889 35816
rect 64748 35776 64754 35788
rect 64877 35785 64889 35788
rect 64923 35785 64935 35819
rect 64877 35779 64935 35785
rect 66530 35776 66536 35828
rect 66588 35816 66594 35828
rect 66625 35819 66683 35825
rect 66625 35816 66637 35819
rect 66588 35788 66637 35816
rect 66588 35776 66594 35788
rect 66625 35785 66637 35788
rect 66671 35785 66683 35819
rect 67266 35816 67272 35828
rect 67227 35788 67272 35816
rect 66625 35779 66683 35785
rect 67266 35776 67272 35788
rect 67324 35776 67330 35828
rect 68370 35776 68376 35828
rect 68428 35816 68434 35828
rect 68465 35819 68523 35825
rect 68465 35816 68477 35819
rect 68428 35788 68477 35816
rect 68428 35776 68434 35788
rect 68465 35785 68477 35788
rect 68511 35785 68523 35819
rect 68465 35779 68523 35785
rect 80882 35776 80888 35828
rect 80940 35816 80946 35828
rect 81161 35819 81219 35825
rect 81161 35816 81173 35819
rect 80940 35788 81173 35816
rect 80940 35776 80946 35788
rect 81161 35785 81173 35788
rect 81207 35785 81219 35819
rect 81161 35779 81219 35785
rect 81342 35776 81348 35828
rect 81400 35816 81406 35828
rect 81713 35819 81771 35825
rect 81713 35816 81725 35819
rect 81400 35788 81725 35816
rect 81400 35776 81406 35788
rect 81713 35785 81725 35788
rect 81759 35785 81771 35819
rect 82354 35816 82360 35828
rect 82315 35788 82360 35816
rect 81713 35779 81771 35785
rect 82354 35776 82360 35788
rect 82412 35776 82418 35828
rect 83826 35816 83832 35828
rect 83787 35788 83832 35816
rect 83826 35776 83832 35788
rect 83884 35776 83890 35828
rect 85209 35819 85267 35825
rect 85209 35785 85221 35819
rect 85255 35816 85267 35819
rect 85298 35816 85304 35828
rect 85255 35788 85304 35816
rect 85255 35785 85267 35788
rect 85209 35779 85267 35785
rect 85298 35776 85304 35788
rect 85356 35776 85362 35828
rect 26786 35708 26792 35760
rect 26844 35748 26850 35760
rect 28902 35748 28908 35760
rect 26844 35720 28908 35748
rect 26844 35708 26850 35720
rect 28902 35708 28908 35720
rect 28960 35708 28966 35760
rect 34238 35748 34244 35760
rect 31726 35720 34244 35748
rect 9582 35640 9588 35692
rect 9640 35680 9646 35692
rect 31726 35680 31754 35720
rect 34238 35708 34244 35720
rect 34296 35708 34302 35760
rect 34330 35708 34336 35760
rect 34388 35748 34394 35760
rect 34517 35751 34575 35757
rect 34517 35748 34529 35751
rect 34388 35720 34529 35748
rect 34388 35708 34394 35720
rect 34517 35717 34529 35720
rect 34563 35748 34575 35751
rect 34563 35720 41414 35748
rect 34563 35717 34575 35720
rect 34517 35711 34575 35717
rect 9640 35652 31754 35680
rect 9640 35640 9646 35652
rect 32950 35640 32956 35692
rect 33008 35680 33014 35692
rect 41230 35680 41236 35692
rect 33008 35652 41236 35680
rect 33008 35640 33014 35652
rect 41230 35640 41236 35652
rect 41288 35640 41294 35692
rect 41386 35680 41414 35720
rect 46750 35708 46756 35760
rect 46808 35748 46814 35760
rect 62117 35751 62175 35757
rect 62117 35748 62129 35751
rect 46808 35720 62129 35748
rect 46808 35708 46814 35720
rect 62117 35717 62129 35720
rect 62163 35748 62175 35751
rect 63586 35748 63592 35760
rect 62163 35720 63592 35748
rect 62163 35717 62175 35720
rect 62117 35711 62175 35717
rect 63586 35708 63592 35720
rect 63644 35708 63650 35760
rect 70486 35708 70492 35760
rect 70544 35748 70550 35760
rect 112070 35748 112076 35760
rect 70544 35720 112076 35748
rect 70544 35708 70550 35720
rect 112070 35708 112076 35720
rect 112128 35708 112134 35760
rect 57422 35680 57428 35692
rect 41386 35652 57428 35680
rect 57422 35640 57428 35652
rect 57480 35640 57486 35692
rect 63773 35683 63831 35689
rect 63773 35649 63785 35683
rect 63819 35680 63831 35683
rect 63862 35680 63868 35692
rect 63819 35652 63868 35680
rect 63819 35649 63831 35652
rect 63773 35643 63831 35649
rect 63862 35640 63868 35652
rect 63920 35680 63926 35692
rect 64782 35680 64788 35692
rect 63920 35652 64788 35680
rect 63920 35640 63926 35652
rect 64782 35640 64788 35652
rect 64840 35640 64846 35692
rect 65242 35640 65248 35692
rect 65300 35680 65306 35692
rect 65337 35683 65395 35689
rect 65337 35680 65349 35683
rect 65300 35652 65349 35680
rect 65300 35640 65306 35652
rect 65337 35649 65349 35652
rect 65383 35680 65395 35683
rect 65981 35683 66039 35689
rect 65981 35680 65993 35683
rect 65383 35652 65993 35680
rect 65383 35649 65395 35652
rect 65337 35643 65395 35649
rect 65981 35649 65993 35652
rect 66027 35649 66039 35683
rect 80422 35680 80428 35692
rect 80383 35652 80428 35680
rect 65981 35643 66039 35649
rect 80422 35640 80428 35652
rect 80480 35680 80486 35692
rect 80977 35683 81035 35689
rect 80977 35680 80989 35683
rect 80480 35652 80989 35680
rect 80480 35640 80486 35652
rect 80977 35649 80989 35652
rect 81023 35649 81035 35683
rect 80977 35643 81035 35649
rect 81894 35640 81900 35692
rect 81952 35680 81958 35692
rect 83090 35680 83096 35692
rect 81952 35652 83096 35680
rect 81952 35640 81958 35652
rect 83090 35640 83096 35652
rect 83148 35640 83154 35692
rect 25130 35572 25136 35624
rect 25188 35612 25194 35624
rect 41138 35612 41144 35624
rect 25188 35584 41144 35612
rect 25188 35572 25194 35584
rect 41138 35572 41144 35584
rect 41196 35572 41202 35624
rect 41414 35572 41420 35624
rect 41472 35612 41478 35624
rect 48406 35612 48412 35624
rect 41472 35584 48412 35612
rect 41472 35572 41478 35584
rect 48406 35572 48412 35584
rect 48464 35572 48470 35624
rect 78953 35615 79011 35621
rect 78953 35581 78965 35615
rect 78999 35612 79011 35615
rect 79502 35612 79508 35624
rect 78999 35584 79508 35612
rect 78999 35581 79011 35584
rect 78953 35575 79011 35581
rect 79502 35572 79508 35584
rect 79560 35612 79566 35624
rect 81342 35612 81348 35624
rect 79560 35584 81348 35612
rect 79560 35572 79566 35584
rect 81342 35572 81348 35584
rect 81400 35572 81406 35624
rect 83642 35572 83648 35624
rect 83700 35612 83706 35624
rect 123478 35612 123484 35624
rect 83700 35584 123484 35612
rect 83700 35572 83706 35584
rect 123478 35572 123484 35584
rect 123536 35572 123542 35624
rect 25777 35547 25835 35553
rect 25777 35544 25789 35547
rect 24596 35516 25789 35544
rect 24596 35488 24624 35516
rect 25777 35513 25789 35516
rect 25823 35513 25835 35547
rect 25777 35507 25835 35513
rect 27890 35504 27896 35556
rect 27948 35544 27954 35556
rect 28077 35547 28135 35553
rect 28077 35544 28089 35547
rect 27948 35516 28089 35544
rect 27948 35504 27954 35516
rect 28077 35513 28089 35516
rect 28123 35544 28135 35547
rect 28123 35516 31064 35544
rect 28123 35513 28135 35516
rect 28077 35507 28135 35513
rect 24213 35479 24271 35485
rect 24213 35445 24225 35479
rect 24259 35476 24271 35479
rect 24578 35476 24584 35488
rect 24259 35448 24584 35476
rect 24259 35445 24271 35448
rect 24213 35439 24271 35445
rect 24578 35436 24584 35448
rect 24636 35436 24642 35488
rect 24765 35479 24823 35485
rect 24765 35445 24777 35479
rect 24811 35476 24823 35479
rect 24854 35476 24860 35488
rect 24811 35448 24860 35476
rect 24811 35445 24823 35448
rect 24765 35439 24823 35445
rect 24854 35436 24860 35448
rect 24912 35436 24918 35488
rect 30834 35436 30840 35488
rect 30892 35476 30898 35488
rect 30929 35479 30987 35485
rect 30929 35476 30941 35479
rect 30892 35448 30941 35476
rect 30892 35436 30898 35448
rect 30929 35445 30941 35448
rect 30975 35445 30987 35479
rect 31036 35476 31064 35516
rect 31294 35504 31300 35556
rect 31352 35544 31358 35556
rect 31938 35544 31944 35556
rect 31352 35516 31944 35544
rect 31352 35504 31358 35516
rect 31938 35504 31944 35516
rect 31996 35544 32002 35556
rect 34698 35544 34704 35556
rect 31996 35516 34704 35544
rect 31996 35504 32002 35516
rect 34698 35504 34704 35516
rect 34756 35504 34762 35556
rect 35802 35544 35808 35556
rect 35763 35516 35808 35544
rect 35802 35504 35808 35516
rect 35860 35504 35866 35556
rect 40865 35547 40923 35553
rect 40865 35544 40877 35547
rect 40236 35516 40877 35544
rect 40236 35488 40264 35516
rect 40865 35513 40877 35516
rect 40911 35513 40923 35547
rect 40865 35507 40923 35513
rect 42518 35504 42524 35556
rect 42576 35544 42582 35556
rect 52086 35544 52092 35556
rect 42576 35516 52092 35544
rect 42576 35504 42582 35516
rect 52086 35504 52092 35516
rect 52144 35504 52150 35556
rect 59357 35547 59415 35553
rect 59357 35513 59369 35547
rect 59403 35544 59415 35547
rect 65521 35547 65579 35553
rect 59403 35516 60504 35544
rect 59403 35513 59415 35516
rect 59357 35507 59415 35513
rect 32950 35476 32956 35488
rect 31036 35448 32956 35476
rect 30929 35439 30987 35445
rect 32950 35436 32956 35448
rect 33008 35436 33014 35488
rect 33134 35476 33140 35488
rect 33095 35448 33140 35476
rect 33134 35436 33140 35448
rect 33192 35436 33198 35488
rect 36909 35479 36967 35485
rect 36909 35445 36921 35479
rect 36955 35476 36967 35479
rect 37274 35476 37280 35488
rect 36955 35448 37280 35476
rect 36955 35445 36967 35448
rect 36909 35439 36967 35445
rect 37274 35436 37280 35448
rect 37332 35476 37338 35488
rect 38102 35476 38108 35488
rect 37332 35448 38108 35476
rect 37332 35436 37338 35448
rect 38102 35436 38108 35448
rect 38160 35436 38166 35488
rect 39853 35479 39911 35485
rect 39853 35445 39865 35479
rect 39899 35476 39911 35479
rect 40218 35476 40224 35488
rect 39899 35448 40224 35476
rect 39899 35445 39911 35448
rect 39853 35439 39911 35445
rect 40218 35436 40224 35448
rect 40276 35436 40282 35488
rect 40405 35479 40463 35485
rect 40405 35445 40417 35479
rect 40451 35476 40463 35479
rect 40954 35476 40960 35488
rect 40451 35448 40960 35476
rect 40451 35445 40463 35448
rect 40405 35439 40463 35445
rect 40954 35436 40960 35448
rect 41012 35476 41018 35488
rect 41417 35479 41475 35485
rect 41417 35476 41429 35479
rect 41012 35448 41429 35476
rect 41012 35436 41018 35448
rect 41417 35445 41429 35448
rect 41463 35445 41475 35479
rect 41417 35439 41475 35445
rect 42061 35479 42119 35485
rect 42061 35445 42073 35479
rect 42107 35476 42119 35479
rect 42794 35476 42800 35488
rect 42107 35448 42800 35476
rect 42107 35445 42119 35448
rect 42061 35439 42119 35445
rect 42794 35436 42800 35448
rect 42852 35436 42858 35488
rect 43441 35479 43499 35485
rect 43441 35445 43453 35479
rect 43487 35476 43499 35479
rect 44358 35476 44364 35488
rect 43487 35448 44364 35476
rect 43487 35445 43499 35448
rect 43441 35439 43499 35445
rect 44358 35436 44364 35448
rect 44416 35476 44422 35488
rect 44453 35479 44511 35485
rect 44453 35476 44465 35479
rect 44416 35448 44465 35476
rect 44416 35436 44422 35448
rect 44453 35445 44465 35448
rect 44499 35445 44511 35479
rect 47118 35476 47124 35488
rect 47079 35448 47124 35476
rect 44453 35439 44511 35445
rect 47118 35436 47124 35448
rect 47176 35436 47182 35488
rect 48130 35476 48136 35488
rect 48091 35448 48136 35476
rect 48130 35436 48136 35448
rect 48188 35436 48194 35488
rect 48590 35476 48596 35488
rect 48551 35448 48596 35476
rect 48590 35436 48596 35448
rect 48648 35436 48654 35488
rect 49694 35436 49700 35488
rect 49752 35476 49758 35488
rect 49881 35479 49939 35485
rect 49881 35476 49893 35479
rect 49752 35448 49893 35476
rect 49752 35436 49758 35448
rect 49881 35445 49893 35448
rect 49927 35445 49939 35479
rect 49881 35439 49939 35445
rect 51626 35436 51632 35488
rect 51684 35476 51690 35488
rect 51813 35479 51871 35485
rect 51813 35476 51825 35479
rect 51684 35448 51825 35476
rect 51684 35436 51690 35448
rect 51813 35445 51825 35448
rect 51859 35476 51871 35479
rect 52730 35476 52736 35488
rect 51859 35448 52736 35476
rect 51859 35445 51871 35448
rect 51813 35439 51871 35445
rect 52730 35436 52736 35448
rect 52788 35476 52794 35488
rect 53098 35476 53104 35488
rect 52788 35448 53104 35476
rect 52788 35436 52794 35448
rect 53098 35436 53104 35448
rect 53156 35436 53162 35488
rect 53926 35436 53932 35488
rect 53984 35476 53990 35488
rect 54021 35479 54079 35485
rect 54021 35476 54033 35479
rect 53984 35448 54033 35476
rect 53984 35436 53990 35448
rect 54021 35445 54033 35448
rect 54067 35445 54079 35479
rect 54021 35439 54079 35445
rect 56045 35479 56103 35485
rect 56045 35445 56057 35479
rect 56091 35476 56103 35479
rect 56594 35476 56600 35488
rect 56091 35448 56600 35476
rect 56091 35445 56103 35448
rect 56045 35439 56103 35445
rect 56594 35436 56600 35448
rect 56652 35436 56658 35488
rect 56965 35479 57023 35485
rect 56965 35445 56977 35479
rect 57011 35476 57023 35479
rect 57330 35476 57336 35488
rect 57011 35448 57336 35476
rect 57011 35445 57023 35448
rect 56965 35439 57023 35445
rect 57330 35436 57336 35448
rect 57388 35476 57394 35488
rect 58713 35479 58771 35485
rect 58713 35476 58725 35479
rect 57388 35448 58725 35476
rect 57388 35436 57394 35448
rect 58713 35445 58725 35448
rect 58759 35476 58771 35479
rect 58894 35476 58900 35488
rect 58759 35448 58900 35476
rect 58759 35445 58771 35448
rect 58713 35439 58771 35445
rect 58894 35436 58900 35448
rect 58952 35436 58958 35488
rect 60476 35476 60504 35516
rect 65521 35513 65533 35547
rect 65567 35544 65579 35547
rect 81434 35544 81440 35556
rect 65567 35516 81440 35544
rect 65567 35513 65579 35516
rect 65521 35507 65579 35513
rect 81434 35504 81440 35516
rect 81492 35504 81498 35556
rect 90450 35504 90456 35556
rect 90508 35544 90514 35556
rect 121546 35544 121552 35556
rect 90508 35516 121552 35544
rect 90508 35504 90514 35516
rect 121546 35504 121552 35516
rect 121604 35504 121610 35556
rect 60734 35476 60740 35488
rect 60476 35448 60740 35476
rect 60734 35436 60740 35448
rect 60792 35436 60798 35488
rect 61565 35479 61623 35485
rect 61565 35445 61577 35479
rect 61611 35476 61623 35479
rect 62022 35476 62028 35488
rect 61611 35448 62028 35476
rect 61611 35445 61623 35448
rect 61565 35439 61623 35445
rect 62022 35436 62028 35448
rect 62080 35436 62086 35488
rect 69198 35476 69204 35488
rect 69159 35448 69204 35476
rect 69198 35436 69204 35448
rect 69256 35476 69262 35488
rect 69753 35479 69811 35485
rect 69753 35476 69765 35479
rect 69256 35448 69765 35476
rect 69256 35436 69262 35448
rect 69753 35445 69765 35448
rect 69799 35445 69811 35479
rect 75086 35476 75092 35488
rect 75047 35448 75092 35476
rect 69753 35439 69811 35445
rect 75086 35436 75092 35448
rect 75144 35436 75150 35488
rect 79965 35479 80023 35485
rect 79965 35445 79977 35479
rect 80011 35476 80023 35479
rect 80054 35476 80060 35488
rect 80011 35448 80060 35476
rect 80011 35445 80023 35448
rect 79965 35439 80023 35445
rect 80054 35436 80060 35448
rect 80112 35436 80118 35488
rect 82906 35476 82912 35488
rect 82867 35448 82912 35476
rect 82906 35436 82912 35448
rect 82964 35476 82970 35488
rect 83918 35476 83924 35488
rect 82964 35448 83924 35476
rect 82964 35436 82970 35448
rect 83918 35436 83924 35448
rect 83976 35476 83982 35488
rect 84381 35479 84439 35485
rect 84381 35476 84393 35479
rect 83976 35448 84393 35476
rect 83976 35436 83982 35448
rect 84381 35445 84393 35448
rect 84427 35445 84439 35479
rect 84381 35439 84439 35445
rect 1104 35386 148856 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 65654 35386
rect 65706 35334 65718 35386
rect 65770 35334 65782 35386
rect 65834 35334 65846 35386
rect 65898 35334 65910 35386
rect 65962 35334 96374 35386
rect 96426 35334 96438 35386
rect 96490 35334 96502 35386
rect 96554 35334 96566 35386
rect 96618 35334 96630 35386
rect 96682 35334 127094 35386
rect 127146 35334 127158 35386
rect 127210 35334 127222 35386
rect 127274 35334 127286 35386
rect 127338 35334 127350 35386
rect 127402 35334 148856 35386
rect 1104 35312 148856 35334
rect 19978 35232 19984 35284
rect 20036 35272 20042 35284
rect 20530 35272 20536 35284
rect 20036 35244 20536 35272
rect 20036 35232 20042 35244
rect 20530 35232 20536 35244
rect 20588 35272 20594 35284
rect 20993 35275 21051 35281
rect 20993 35272 21005 35275
rect 20588 35244 21005 35272
rect 20588 35232 20594 35244
rect 20993 35241 21005 35244
rect 21039 35241 21051 35275
rect 20993 35235 21051 35241
rect 24486 35232 24492 35284
rect 24544 35272 24550 35284
rect 24765 35275 24823 35281
rect 24765 35272 24777 35275
rect 24544 35244 24777 35272
rect 24544 35232 24550 35244
rect 24765 35241 24777 35244
rect 24811 35241 24823 35275
rect 24765 35235 24823 35241
rect 24854 35232 24860 35284
rect 24912 35272 24918 35284
rect 25498 35272 25504 35284
rect 24912 35244 25504 35272
rect 24912 35232 24918 35244
rect 25498 35232 25504 35244
rect 25556 35272 25562 35284
rect 25961 35275 26019 35281
rect 25961 35272 25973 35275
rect 25556 35244 25973 35272
rect 25556 35232 25562 35244
rect 25961 35241 25973 35244
rect 26007 35241 26019 35275
rect 28718 35272 28724 35284
rect 28679 35244 28724 35272
rect 25961 35235 26019 35241
rect 28718 35232 28724 35244
rect 28776 35232 28782 35284
rect 75914 35272 75920 35284
rect 30300 35244 75920 35272
rect 25222 35164 25228 35216
rect 25280 35204 25286 35216
rect 30300 35204 30328 35244
rect 75914 35232 75920 35244
rect 75972 35232 75978 35284
rect 79502 35272 79508 35284
rect 79463 35244 79508 35272
rect 79502 35232 79508 35244
rect 79560 35232 79566 35284
rect 79594 35232 79600 35284
rect 79652 35272 79658 35284
rect 80057 35275 80115 35281
rect 80057 35272 80069 35275
rect 79652 35244 80069 35272
rect 79652 35232 79658 35244
rect 80057 35241 80069 35244
rect 80103 35241 80115 35275
rect 80057 35235 80115 35241
rect 80238 35232 80244 35284
rect 80296 35272 80302 35284
rect 80609 35275 80667 35281
rect 80609 35272 80621 35275
rect 80296 35244 80621 35272
rect 80296 35232 80302 35244
rect 80609 35241 80621 35244
rect 80655 35241 80667 35275
rect 81342 35272 81348 35284
rect 81303 35244 81348 35272
rect 80609 35235 80667 35241
rect 81342 35232 81348 35244
rect 81400 35272 81406 35284
rect 81805 35275 81863 35281
rect 81805 35272 81817 35275
rect 81400 35244 81817 35272
rect 81400 35232 81406 35244
rect 81805 35241 81817 35244
rect 81851 35272 81863 35275
rect 82357 35275 82415 35281
rect 82357 35272 82369 35275
rect 81851 35244 82369 35272
rect 81851 35241 81863 35244
rect 81805 35235 81863 35241
rect 82357 35241 82369 35244
rect 82403 35241 82415 35275
rect 82357 35235 82415 35241
rect 84746 35232 84752 35284
rect 84804 35272 84810 35284
rect 140682 35272 140688 35284
rect 84804 35244 140688 35272
rect 84804 35232 84810 35244
rect 140682 35232 140688 35244
rect 140740 35232 140746 35284
rect 25280 35176 30328 35204
rect 25280 35164 25286 35176
rect 35526 35164 35532 35216
rect 35584 35204 35590 35216
rect 35989 35207 36047 35213
rect 35989 35204 36001 35207
rect 35584 35176 36001 35204
rect 35584 35164 35590 35176
rect 35989 35173 36001 35176
rect 36035 35173 36047 35207
rect 35989 35167 36047 35173
rect 36630 35164 36636 35216
rect 36688 35204 36694 35216
rect 37553 35207 37611 35213
rect 37553 35204 37565 35207
rect 36688 35176 37565 35204
rect 36688 35164 36694 35176
rect 37553 35173 37565 35176
rect 37599 35173 37611 35207
rect 41690 35204 41696 35216
rect 41651 35176 41696 35204
rect 37553 35167 37611 35173
rect 41690 35164 41696 35176
rect 41748 35164 41754 35216
rect 43070 35164 43076 35216
rect 43128 35204 43134 35216
rect 43441 35207 43499 35213
rect 43441 35204 43453 35207
rect 43128 35176 43453 35204
rect 43128 35164 43134 35176
rect 43441 35173 43453 35176
rect 43487 35173 43499 35207
rect 43441 35167 43499 35173
rect 43990 35164 43996 35216
rect 44048 35204 44054 35216
rect 44177 35207 44235 35213
rect 44177 35204 44189 35207
rect 44048 35176 44189 35204
rect 44048 35164 44054 35176
rect 44177 35173 44189 35176
rect 44223 35173 44235 35207
rect 44177 35167 44235 35173
rect 44284 35176 70394 35204
rect 35342 35096 35348 35148
rect 35400 35136 35406 35148
rect 44284 35136 44312 35176
rect 35400 35108 44312 35136
rect 35400 35096 35406 35108
rect 44450 35096 44456 35148
rect 44508 35136 44514 35148
rect 57054 35136 57060 35148
rect 44508 35108 57060 35136
rect 44508 35096 44514 35108
rect 57054 35096 57060 35108
rect 57112 35096 57118 35148
rect 58526 35096 58532 35148
rect 58584 35136 58590 35148
rect 58897 35139 58955 35145
rect 58897 35136 58909 35139
rect 58584 35108 58909 35136
rect 58584 35096 58590 35108
rect 58897 35105 58909 35108
rect 58943 35105 58955 35139
rect 59906 35136 59912 35148
rect 59867 35108 59912 35136
rect 58897 35099 58955 35105
rect 59906 35096 59912 35108
rect 59964 35096 59970 35148
rect 62114 35096 62120 35148
rect 62172 35136 62178 35148
rect 62301 35139 62359 35145
rect 62301 35136 62313 35139
rect 62172 35108 62313 35136
rect 62172 35096 62178 35108
rect 62301 35105 62313 35108
rect 62347 35105 62359 35139
rect 62301 35099 62359 35105
rect 62850 35096 62856 35148
rect 62908 35136 62914 35148
rect 62945 35139 63003 35145
rect 62945 35136 62957 35139
rect 62908 35108 62957 35136
rect 62908 35096 62914 35108
rect 62945 35105 62957 35108
rect 62991 35105 63003 35139
rect 62945 35099 63003 35105
rect 64138 35096 64144 35148
rect 64196 35136 64202 35148
rect 64233 35139 64291 35145
rect 64233 35136 64245 35139
rect 64196 35108 64245 35136
rect 64196 35096 64202 35108
rect 64233 35105 64245 35108
rect 64279 35105 64291 35139
rect 64233 35099 64291 35105
rect 65334 35096 65340 35148
rect 65392 35136 65398 35148
rect 65889 35139 65947 35145
rect 65889 35136 65901 35139
rect 65392 35108 65901 35136
rect 65392 35096 65398 35108
rect 65889 35105 65901 35108
rect 65935 35105 65947 35139
rect 65889 35099 65947 35105
rect 68554 35096 68560 35148
rect 68612 35136 68618 35148
rect 69201 35139 69259 35145
rect 69201 35136 69213 35139
rect 68612 35108 69213 35136
rect 68612 35096 68618 35108
rect 69201 35105 69213 35108
rect 69247 35105 69259 35139
rect 69201 35099 69259 35105
rect 17954 35028 17960 35080
rect 18012 35068 18018 35080
rect 36538 35068 36544 35080
rect 18012 35040 36544 35068
rect 18012 35028 18018 35040
rect 36538 35028 36544 35040
rect 36596 35028 36602 35080
rect 36906 35028 36912 35080
rect 36964 35068 36970 35080
rect 37001 35071 37059 35077
rect 37001 35068 37013 35071
rect 36964 35040 37013 35068
rect 36964 35028 36970 35040
rect 37001 35037 37013 35040
rect 37047 35068 37059 35071
rect 43346 35068 43352 35080
rect 37047 35040 43352 35068
rect 37047 35037 37059 35040
rect 37001 35031 37059 35037
rect 43346 35028 43352 35040
rect 43404 35028 43410 35080
rect 44542 35028 44548 35080
rect 44600 35068 44606 35080
rect 63678 35068 63684 35080
rect 44600 35040 63684 35068
rect 44600 35028 44606 35040
rect 63678 35028 63684 35040
rect 63736 35028 63742 35080
rect 65242 35068 65248 35080
rect 65203 35040 65248 35068
rect 65242 35028 65248 35040
rect 65300 35028 65306 35080
rect 70366 35068 70394 35176
rect 75196 35176 80054 35204
rect 75196 35068 75224 35176
rect 80026 35148 80054 35176
rect 80026 35108 80060 35148
rect 80054 35096 80060 35108
rect 80112 35096 80118 35148
rect 70366 35040 75224 35068
rect 30650 34960 30656 35012
rect 30708 35000 30714 35012
rect 44450 35000 44456 35012
rect 30708 34972 44456 35000
rect 30708 34960 30714 34972
rect 44450 34960 44456 34972
rect 44508 34960 44514 35012
rect 47118 35000 47124 35012
rect 44652 34972 47124 35000
rect 25314 34892 25320 34944
rect 25372 34932 25378 34944
rect 25501 34935 25559 34941
rect 25501 34932 25513 34935
rect 25372 34904 25513 34932
rect 25372 34892 25378 34904
rect 25501 34901 25513 34904
rect 25547 34932 25559 34935
rect 25682 34932 25688 34944
rect 25547 34904 25688 34932
rect 25547 34901 25559 34904
rect 25501 34895 25559 34901
rect 25682 34892 25688 34904
rect 25740 34892 25746 34944
rect 38841 34935 38899 34941
rect 38841 34901 38853 34935
rect 38887 34932 38899 34935
rect 40681 34935 40739 34941
rect 40681 34932 40693 34935
rect 38887 34904 40693 34932
rect 38887 34901 38899 34904
rect 38841 34895 38899 34901
rect 40681 34901 40693 34904
rect 40727 34932 40739 34935
rect 40862 34932 40868 34944
rect 40727 34904 40868 34932
rect 40727 34901 40739 34904
rect 40681 34895 40739 34901
rect 40862 34892 40868 34904
rect 40920 34932 40926 34944
rect 42794 34932 42800 34944
rect 40920 34904 42800 34932
rect 40920 34892 40926 34904
rect 42794 34892 42800 34904
rect 42852 34932 42858 34944
rect 44652 34932 44680 34972
rect 47118 34960 47124 34972
rect 47176 35000 47182 35012
rect 47673 35003 47731 35009
rect 47673 35000 47685 35003
rect 47176 34972 47685 35000
rect 47176 34960 47182 34972
rect 47673 34969 47685 34972
rect 47719 34969 47731 35003
rect 47673 34963 47731 34969
rect 48222 34960 48228 35012
rect 48280 35000 48286 35012
rect 48593 35003 48651 35009
rect 48593 35000 48605 35003
rect 48280 34972 48605 35000
rect 48280 34960 48286 34972
rect 48593 34969 48605 34972
rect 48639 34969 48651 35003
rect 48593 34963 48651 34969
rect 49786 34960 49792 35012
rect 49844 35000 49850 35012
rect 50341 35003 50399 35009
rect 50341 35000 50353 35003
rect 49844 34972 50353 35000
rect 49844 34960 49850 34972
rect 50341 34969 50353 34972
rect 50387 34969 50399 35003
rect 50341 34963 50399 34969
rect 51166 34960 51172 35012
rect 51224 35000 51230 35012
rect 51261 35003 51319 35009
rect 51261 35000 51273 35003
rect 51224 34972 51273 35000
rect 51224 34960 51230 34972
rect 51261 34969 51273 34972
rect 51307 34969 51319 35003
rect 51261 34963 51319 34969
rect 53190 34960 53196 35012
rect 53248 35000 53254 35012
rect 53837 35003 53895 35009
rect 53837 35000 53849 35003
rect 53248 34972 53849 35000
rect 53248 34960 53254 34972
rect 53837 34969 53849 34972
rect 53883 34969 53895 35003
rect 53837 34963 53895 34969
rect 54386 34960 54392 35012
rect 54444 35000 54450 35012
rect 92382 35000 92388 35012
rect 54444 34972 92388 35000
rect 54444 34960 54450 34972
rect 92382 34960 92388 34972
rect 92440 34960 92446 35012
rect 45646 34932 45652 34944
rect 42852 34904 44680 34932
rect 45559 34904 45652 34932
rect 42852 34892 42858 34904
rect 45646 34892 45652 34904
rect 45704 34932 45710 34944
rect 46014 34932 46020 34944
rect 45704 34904 46020 34932
rect 45704 34892 45710 34904
rect 46014 34892 46020 34904
rect 46072 34892 46078 34944
rect 60734 34892 60740 34944
rect 60792 34932 60798 34944
rect 61194 34932 61200 34944
rect 60792 34904 60837 34932
rect 61155 34904 61200 34932
rect 60792 34892 60798 34904
rect 61194 34892 61200 34904
rect 61252 34932 61258 34944
rect 61746 34932 61752 34944
rect 61252 34904 61752 34932
rect 61252 34892 61258 34904
rect 61746 34892 61752 34904
rect 61804 34892 61810 34944
rect 61841 34935 61899 34941
rect 61841 34901 61853 34935
rect 61887 34932 61899 34935
rect 62022 34932 62028 34944
rect 61887 34904 62028 34932
rect 61887 34901 61899 34904
rect 61841 34895 61899 34901
rect 62022 34892 62028 34904
rect 62080 34892 62086 34944
rect 62574 34892 62580 34944
rect 62632 34932 62638 34944
rect 63681 34935 63739 34941
rect 63681 34932 63693 34935
rect 62632 34904 63693 34932
rect 62632 34892 62638 34904
rect 63681 34901 63693 34904
rect 63727 34932 63739 34935
rect 64230 34932 64236 34944
rect 63727 34904 64236 34932
rect 63727 34901 63739 34904
rect 63681 34895 63739 34901
rect 64230 34892 64236 34904
rect 64288 34892 64294 34944
rect 1104 34842 148856 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 81014 34842
rect 81066 34790 81078 34842
rect 81130 34790 81142 34842
rect 81194 34790 81206 34842
rect 81258 34790 81270 34842
rect 81322 34790 111734 34842
rect 111786 34790 111798 34842
rect 111850 34790 111862 34842
rect 111914 34790 111926 34842
rect 111978 34790 111990 34842
rect 112042 34790 142454 34842
rect 142506 34790 142518 34842
rect 142570 34790 142582 34842
rect 142634 34790 142646 34842
rect 142698 34790 142710 34842
rect 142762 34790 148856 34842
rect 1104 34768 148856 34790
rect 29086 34688 29092 34740
rect 29144 34728 29150 34740
rect 47026 34728 47032 34740
rect 29144 34700 47032 34728
rect 29144 34688 29150 34700
rect 47026 34688 47032 34700
rect 47084 34688 47090 34740
rect 59262 34688 59268 34740
rect 59320 34728 59326 34740
rect 102870 34728 102876 34740
rect 59320 34700 102876 34728
rect 59320 34688 59326 34700
rect 102870 34688 102876 34700
rect 102928 34688 102934 34740
rect 43806 34660 43812 34672
rect 43767 34632 43812 34660
rect 43806 34620 43812 34632
rect 43864 34620 43870 34672
rect 24578 34484 24584 34536
rect 24636 34524 24642 34536
rect 24762 34524 24768 34536
rect 24636 34496 24768 34524
rect 24636 34484 24642 34496
rect 24762 34484 24768 34496
rect 24820 34484 24826 34536
rect 69014 34484 69020 34536
rect 69072 34524 69078 34536
rect 69198 34524 69204 34536
rect 69072 34496 69204 34524
rect 69072 34484 69078 34496
rect 69198 34484 69204 34496
rect 69256 34484 69262 34536
rect 57514 34416 57520 34468
rect 57572 34456 57578 34468
rect 124030 34456 124036 34468
rect 57572 34428 124036 34456
rect 57572 34416 57578 34428
rect 124030 34416 124036 34428
rect 124088 34416 124094 34468
rect 83090 34348 83096 34400
rect 83148 34388 83154 34400
rect 143994 34388 144000 34400
rect 83148 34360 144000 34388
rect 83148 34348 83154 34360
rect 143994 34348 144000 34360
rect 144052 34348 144058 34400
rect 1104 34298 148856 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 65654 34298
rect 65706 34246 65718 34298
rect 65770 34246 65782 34298
rect 65834 34246 65846 34298
rect 65898 34246 65910 34298
rect 65962 34246 96374 34298
rect 96426 34246 96438 34298
rect 96490 34246 96502 34298
rect 96554 34246 96566 34298
rect 96618 34246 96630 34298
rect 96682 34246 127094 34298
rect 127146 34246 127158 34298
rect 127210 34246 127222 34298
rect 127274 34246 127286 34298
rect 127338 34246 127350 34298
rect 127402 34246 148856 34298
rect 1104 34224 148856 34246
rect 75822 34144 75828 34196
rect 75880 34184 75886 34196
rect 113450 34184 113456 34196
rect 75880 34156 113456 34184
rect 75880 34144 75886 34156
rect 113450 34144 113456 34156
rect 113508 34144 113514 34196
rect 38838 34076 38844 34128
rect 38896 34116 38902 34128
rect 81894 34116 81900 34128
rect 38896 34088 81900 34116
rect 38896 34076 38902 34088
rect 81894 34076 81900 34088
rect 81952 34076 81958 34128
rect 81986 34076 81992 34128
rect 82044 34116 82050 34128
rect 83826 34116 83832 34128
rect 82044 34088 83832 34116
rect 82044 34076 82050 34088
rect 83826 34076 83832 34088
rect 83884 34076 83890 34128
rect 61010 34008 61016 34060
rect 61068 34048 61074 34060
rect 107746 34048 107752 34060
rect 61068 34020 107752 34048
rect 61068 34008 61074 34020
rect 107746 34008 107752 34020
rect 107804 34008 107810 34060
rect 66070 33940 66076 33992
rect 66128 33980 66134 33992
rect 109586 33980 109592 33992
rect 66128 33952 109592 33980
rect 66128 33940 66134 33952
rect 109586 33940 109592 33952
rect 109644 33940 109650 33992
rect 69658 33872 69664 33924
rect 69716 33912 69722 33924
rect 112162 33912 112168 33924
rect 69716 33884 112168 33912
rect 69716 33872 69722 33884
rect 112162 33872 112168 33884
rect 112220 33872 112226 33924
rect 72602 33804 72608 33856
rect 72660 33844 72666 33856
rect 105906 33844 105912 33856
rect 72660 33816 105912 33844
rect 72660 33804 72666 33816
rect 105906 33804 105912 33816
rect 105964 33804 105970 33856
rect 1104 33754 148856 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 81014 33754
rect 81066 33702 81078 33754
rect 81130 33702 81142 33754
rect 81194 33702 81206 33754
rect 81258 33702 81270 33754
rect 81322 33702 111734 33754
rect 111786 33702 111798 33754
rect 111850 33702 111862 33754
rect 111914 33702 111926 33754
rect 111978 33702 111990 33754
rect 112042 33702 142454 33754
rect 142506 33702 142518 33754
rect 142570 33702 142582 33754
rect 142634 33702 142646 33754
rect 142698 33702 142710 33754
rect 142762 33702 148856 33754
rect 1104 33680 148856 33702
rect 46198 33600 46204 33652
rect 46256 33640 46262 33652
rect 79134 33640 79140 33652
rect 46256 33612 79140 33640
rect 46256 33600 46262 33612
rect 79134 33600 79140 33612
rect 79192 33600 79198 33652
rect 81894 33600 81900 33652
rect 81952 33640 81958 33652
rect 89622 33640 89628 33652
rect 81952 33612 89628 33640
rect 81952 33600 81958 33612
rect 89622 33600 89628 33612
rect 89680 33600 89686 33652
rect 25958 33532 25964 33584
rect 26016 33572 26022 33584
rect 86862 33572 86868 33584
rect 26016 33544 86868 33572
rect 26016 33532 26022 33544
rect 86862 33532 86868 33544
rect 86920 33532 86926 33584
rect 21358 33464 21364 33516
rect 21416 33504 21422 33516
rect 83182 33504 83188 33516
rect 21416 33476 83188 33504
rect 21416 33464 21422 33476
rect 83182 33464 83188 33476
rect 83240 33464 83246 33516
rect 1104 33210 148856 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 65654 33210
rect 65706 33158 65718 33210
rect 65770 33158 65782 33210
rect 65834 33158 65846 33210
rect 65898 33158 65910 33210
rect 65962 33158 96374 33210
rect 96426 33158 96438 33210
rect 96490 33158 96502 33210
rect 96554 33158 96566 33210
rect 96618 33158 96630 33210
rect 96682 33158 127094 33210
rect 127146 33158 127158 33210
rect 127210 33158 127222 33210
rect 127274 33158 127286 33210
rect 127338 33158 127350 33210
rect 127402 33158 148856 33210
rect 1104 33136 148856 33158
rect 55858 33056 55864 33108
rect 55916 33096 55922 33108
rect 56778 33096 56784 33108
rect 55916 33068 56784 33096
rect 55916 33056 55922 33068
rect 56778 33056 56784 33068
rect 56836 33056 56842 33108
rect 77754 33056 77760 33108
rect 77812 33096 77818 33108
rect 147398 33096 147404 33108
rect 77812 33068 147404 33096
rect 77812 33056 77818 33068
rect 147398 33056 147404 33068
rect 147456 33056 147462 33108
rect 51534 32988 51540 33040
rect 51592 33028 51598 33040
rect 114554 33028 114560 33040
rect 51592 33000 114560 33028
rect 51592 32988 51598 33000
rect 114554 32988 114560 33000
rect 114612 32988 114618 33040
rect 26510 32920 26516 32972
rect 26568 32960 26574 32972
rect 88058 32960 88064 32972
rect 26568 32932 88064 32960
rect 26568 32920 26574 32932
rect 88058 32920 88064 32932
rect 88116 32920 88122 32972
rect 48130 32852 48136 32904
rect 48188 32892 48194 32904
rect 108758 32892 108764 32904
rect 48188 32864 108764 32892
rect 48188 32852 48194 32864
rect 108758 32852 108764 32864
rect 108816 32852 108822 32904
rect 32490 32784 32496 32836
rect 32548 32824 32554 32836
rect 91554 32824 91560 32836
rect 32548 32796 91560 32824
rect 32548 32784 32554 32796
rect 91554 32784 91560 32796
rect 91612 32784 91618 32836
rect 44818 32716 44824 32768
rect 44876 32756 44882 32768
rect 97994 32756 98000 32768
rect 44876 32728 98000 32756
rect 44876 32716 44882 32728
rect 97994 32716 98000 32728
rect 98052 32716 98058 32768
rect 1104 32666 148856 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 81014 32666
rect 81066 32614 81078 32666
rect 81130 32614 81142 32666
rect 81194 32614 81206 32666
rect 81258 32614 81270 32666
rect 81322 32614 111734 32666
rect 111786 32614 111798 32666
rect 111850 32614 111862 32666
rect 111914 32614 111926 32666
rect 111978 32614 111990 32666
rect 112042 32614 142454 32666
rect 142506 32614 142518 32666
rect 142570 32614 142582 32666
rect 142634 32614 142646 32666
rect 142698 32614 142710 32666
rect 142762 32614 148856 32666
rect 1104 32592 148856 32614
rect 100754 32552 100760 32564
rect 51046 32524 100760 32552
rect 49142 32376 49148 32428
rect 49200 32416 49206 32428
rect 51046 32416 51074 32524
rect 100754 32512 100760 32524
rect 100812 32512 100818 32564
rect 52914 32444 52920 32496
rect 52972 32484 52978 32496
rect 104434 32484 104440 32496
rect 52972 32456 104440 32484
rect 52972 32444 52978 32456
rect 104434 32444 104440 32456
rect 104492 32444 104498 32496
rect 106274 32416 106280 32428
rect 49200 32388 51074 32416
rect 60706 32388 106280 32416
rect 49200 32376 49206 32388
rect 57146 32308 57152 32360
rect 57204 32348 57210 32360
rect 60706 32348 60734 32388
rect 106274 32376 106280 32388
rect 106332 32376 106338 32428
rect 57204 32320 60734 32348
rect 57204 32308 57210 32320
rect 1104 32122 148856 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 65654 32122
rect 65706 32070 65718 32122
rect 65770 32070 65782 32122
rect 65834 32070 65846 32122
rect 65898 32070 65910 32122
rect 65962 32070 96374 32122
rect 96426 32070 96438 32122
rect 96490 32070 96502 32122
rect 96554 32070 96566 32122
rect 96618 32070 96630 32122
rect 96682 32070 127094 32122
rect 127146 32070 127158 32122
rect 127210 32070 127222 32122
rect 127274 32070 127286 32122
rect 127338 32070 127350 32122
rect 127402 32070 148856 32122
rect 1104 32048 148856 32070
rect 62666 31696 62672 31748
rect 62724 31736 62730 31748
rect 96154 31736 96160 31748
rect 62724 31708 96160 31736
rect 62724 31696 62730 31708
rect 96154 31696 96160 31708
rect 96212 31696 96218 31748
rect 1104 31578 148856 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 81014 31578
rect 81066 31526 81078 31578
rect 81130 31526 81142 31578
rect 81194 31526 81206 31578
rect 81258 31526 81270 31578
rect 81322 31526 111734 31578
rect 111786 31526 111798 31578
rect 111850 31526 111862 31578
rect 111914 31526 111926 31578
rect 111978 31526 111990 31578
rect 112042 31526 142454 31578
rect 142506 31526 142518 31578
rect 142570 31526 142582 31578
rect 142634 31526 142646 31578
rect 142698 31526 142710 31578
rect 142762 31526 148856 31578
rect 1104 31504 148856 31526
rect 1104 31034 148856 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 65654 31034
rect 65706 30982 65718 31034
rect 65770 30982 65782 31034
rect 65834 30982 65846 31034
rect 65898 30982 65910 31034
rect 65962 30982 96374 31034
rect 96426 30982 96438 31034
rect 96490 30982 96502 31034
rect 96554 30982 96566 31034
rect 96618 30982 96630 31034
rect 96682 30982 127094 31034
rect 127146 30982 127158 31034
rect 127210 30982 127222 31034
rect 127274 30982 127286 31034
rect 127338 30982 127350 31034
rect 127402 30982 148856 31034
rect 1104 30960 148856 30982
rect 1104 30490 148856 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 81014 30490
rect 81066 30438 81078 30490
rect 81130 30438 81142 30490
rect 81194 30438 81206 30490
rect 81258 30438 81270 30490
rect 81322 30438 111734 30490
rect 111786 30438 111798 30490
rect 111850 30438 111862 30490
rect 111914 30438 111926 30490
rect 111978 30438 111990 30490
rect 112042 30438 142454 30490
rect 142506 30438 142518 30490
rect 142570 30438 142582 30490
rect 142634 30438 142646 30490
rect 142698 30438 142710 30490
rect 142762 30438 148856 30490
rect 1104 30416 148856 30438
rect 1104 29946 148856 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 65654 29946
rect 65706 29894 65718 29946
rect 65770 29894 65782 29946
rect 65834 29894 65846 29946
rect 65898 29894 65910 29946
rect 65962 29894 96374 29946
rect 96426 29894 96438 29946
rect 96490 29894 96502 29946
rect 96554 29894 96566 29946
rect 96618 29894 96630 29946
rect 96682 29894 127094 29946
rect 127146 29894 127158 29946
rect 127210 29894 127222 29946
rect 127274 29894 127286 29946
rect 127338 29894 127350 29946
rect 127402 29894 148856 29946
rect 1104 29872 148856 29894
rect 31754 29588 31760 29640
rect 31812 29628 31818 29640
rect 61194 29628 61200 29640
rect 31812 29600 61200 29628
rect 31812 29588 31818 29600
rect 61194 29588 61200 29600
rect 61252 29588 61258 29640
rect 1104 29402 148856 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 81014 29402
rect 81066 29350 81078 29402
rect 81130 29350 81142 29402
rect 81194 29350 81206 29402
rect 81258 29350 81270 29402
rect 81322 29350 111734 29402
rect 111786 29350 111798 29402
rect 111850 29350 111862 29402
rect 111914 29350 111926 29402
rect 111978 29350 111990 29402
rect 112042 29350 142454 29402
rect 142506 29350 142518 29402
rect 142570 29350 142582 29402
rect 142634 29350 142646 29402
rect 142698 29350 142710 29402
rect 142762 29350 148856 29402
rect 1104 29328 148856 29350
rect 1104 28858 148856 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 65654 28858
rect 65706 28806 65718 28858
rect 65770 28806 65782 28858
rect 65834 28806 65846 28858
rect 65898 28806 65910 28858
rect 65962 28806 96374 28858
rect 96426 28806 96438 28858
rect 96490 28806 96502 28858
rect 96554 28806 96566 28858
rect 96618 28806 96630 28858
rect 96682 28806 127094 28858
rect 127146 28806 127158 28858
rect 127210 28806 127222 28858
rect 127274 28806 127286 28858
rect 127338 28806 127350 28858
rect 127402 28806 148856 28858
rect 1104 28784 148856 28806
rect 1104 28314 148856 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 81014 28314
rect 81066 28262 81078 28314
rect 81130 28262 81142 28314
rect 81194 28262 81206 28314
rect 81258 28262 81270 28314
rect 81322 28262 111734 28314
rect 111786 28262 111798 28314
rect 111850 28262 111862 28314
rect 111914 28262 111926 28314
rect 111978 28262 111990 28314
rect 112042 28262 142454 28314
rect 142506 28262 142518 28314
rect 142570 28262 142582 28314
rect 142634 28262 142646 28314
rect 142698 28262 142710 28314
rect 142762 28262 148856 28314
rect 1104 28240 148856 28262
rect 1104 27770 148856 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 65654 27770
rect 65706 27718 65718 27770
rect 65770 27718 65782 27770
rect 65834 27718 65846 27770
rect 65898 27718 65910 27770
rect 65962 27718 96374 27770
rect 96426 27718 96438 27770
rect 96490 27718 96502 27770
rect 96554 27718 96566 27770
rect 96618 27718 96630 27770
rect 96682 27718 127094 27770
rect 127146 27718 127158 27770
rect 127210 27718 127222 27770
rect 127274 27718 127286 27770
rect 127338 27718 127350 27770
rect 127402 27718 148856 27770
rect 1104 27696 148856 27718
rect 1104 27226 148856 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 81014 27226
rect 81066 27174 81078 27226
rect 81130 27174 81142 27226
rect 81194 27174 81206 27226
rect 81258 27174 81270 27226
rect 81322 27174 111734 27226
rect 111786 27174 111798 27226
rect 111850 27174 111862 27226
rect 111914 27174 111926 27226
rect 111978 27174 111990 27226
rect 112042 27174 142454 27226
rect 142506 27174 142518 27226
rect 142570 27174 142582 27226
rect 142634 27174 142646 27226
rect 142698 27174 142710 27226
rect 142762 27174 148856 27226
rect 1104 27152 148856 27174
rect 1104 26682 148856 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 65654 26682
rect 65706 26630 65718 26682
rect 65770 26630 65782 26682
rect 65834 26630 65846 26682
rect 65898 26630 65910 26682
rect 65962 26630 96374 26682
rect 96426 26630 96438 26682
rect 96490 26630 96502 26682
rect 96554 26630 96566 26682
rect 96618 26630 96630 26682
rect 96682 26630 127094 26682
rect 127146 26630 127158 26682
rect 127210 26630 127222 26682
rect 127274 26630 127286 26682
rect 127338 26630 127350 26682
rect 127402 26630 148856 26682
rect 1104 26608 148856 26630
rect 1104 26138 148856 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 81014 26138
rect 81066 26086 81078 26138
rect 81130 26086 81142 26138
rect 81194 26086 81206 26138
rect 81258 26086 81270 26138
rect 81322 26086 111734 26138
rect 111786 26086 111798 26138
rect 111850 26086 111862 26138
rect 111914 26086 111926 26138
rect 111978 26086 111990 26138
rect 112042 26086 142454 26138
rect 142506 26086 142518 26138
rect 142570 26086 142582 26138
rect 142634 26086 142646 26138
rect 142698 26086 142710 26138
rect 142762 26086 148856 26138
rect 1104 26064 148856 26086
rect 1104 25594 148856 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 65654 25594
rect 65706 25542 65718 25594
rect 65770 25542 65782 25594
rect 65834 25542 65846 25594
rect 65898 25542 65910 25594
rect 65962 25542 96374 25594
rect 96426 25542 96438 25594
rect 96490 25542 96502 25594
rect 96554 25542 96566 25594
rect 96618 25542 96630 25594
rect 96682 25542 127094 25594
rect 127146 25542 127158 25594
rect 127210 25542 127222 25594
rect 127274 25542 127286 25594
rect 127338 25542 127350 25594
rect 127402 25542 148856 25594
rect 1104 25520 148856 25542
rect 1104 25050 148856 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 81014 25050
rect 81066 24998 81078 25050
rect 81130 24998 81142 25050
rect 81194 24998 81206 25050
rect 81258 24998 81270 25050
rect 81322 24998 111734 25050
rect 111786 24998 111798 25050
rect 111850 24998 111862 25050
rect 111914 24998 111926 25050
rect 111978 24998 111990 25050
rect 112042 24998 142454 25050
rect 142506 24998 142518 25050
rect 142570 24998 142582 25050
rect 142634 24998 142646 25050
rect 142698 24998 142710 25050
rect 142762 24998 148856 25050
rect 1104 24976 148856 24998
rect 1104 24506 148856 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 65654 24506
rect 65706 24454 65718 24506
rect 65770 24454 65782 24506
rect 65834 24454 65846 24506
rect 65898 24454 65910 24506
rect 65962 24454 96374 24506
rect 96426 24454 96438 24506
rect 96490 24454 96502 24506
rect 96554 24454 96566 24506
rect 96618 24454 96630 24506
rect 96682 24454 127094 24506
rect 127146 24454 127158 24506
rect 127210 24454 127222 24506
rect 127274 24454 127286 24506
rect 127338 24454 127350 24506
rect 127402 24454 148856 24506
rect 1104 24432 148856 24454
rect 73706 24148 73712 24200
rect 73764 24188 73770 24200
rect 75086 24188 75092 24200
rect 73764 24160 75092 24188
rect 73764 24148 73770 24160
rect 75086 24148 75092 24160
rect 75144 24148 75150 24200
rect 1104 23962 148856 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 81014 23962
rect 81066 23910 81078 23962
rect 81130 23910 81142 23962
rect 81194 23910 81206 23962
rect 81258 23910 81270 23962
rect 81322 23910 111734 23962
rect 111786 23910 111798 23962
rect 111850 23910 111862 23962
rect 111914 23910 111926 23962
rect 111978 23910 111990 23962
rect 112042 23910 142454 23962
rect 142506 23910 142518 23962
rect 142570 23910 142582 23962
rect 142634 23910 142646 23962
rect 142698 23910 142710 23962
rect 142762 23910 148856 23962
rect 1104 23888 148856 23910
rect 1104 23418 148856 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 65654 23418
rect 65706 23366 65718 23418
rect 65770 23366 65782 23418
rect 65834 23366 65846 23418
rect 65898 23366 65910 23418
rect 65962 23366 96374 23418
rect 96426 23366 96438 23418
rect 96490 23366 96502 23418
rect 96554 23366 96566 23418
rect 96618 23366 96630 23418
rect 96682 23366 127094 23418
rect 127146 23366 127158 23418
rect 127210 23366 127222 23418
rect 127274 23366 127286 23418
rect 127338 23366 127350 23418
rect 127402 23366 148856 23418
rect 1104 23344 148856 23366
rect 1104 22874 148856 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 81014 22874
rect 81066 22822 81078 22874
rect 81130 22822 81142 22874
rect 81194 22822 81206 22874
rect 81258 22822 81270 22874
rect 81322 22822 111734 22874
rect 111786 22822 111798 22874
rect 111850 22822 111862 22874
rect 111914 22822 111926 22874
rect 111978 22822 111990 22874
rect 112042 22822 142454 22874
rect 142506 22822 142518 22874
rect 142570 22822 142582 22874
rect 142634 22822 142646 22874
rect 142698 22822 142710 22874
rect 142762 22822 148856 22874
rect 1104 22800 148856 22822
rect 1104 22330 148856 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 65654 22330
rect 65706 22278 65718 22330
rect 65770 22278 65782 22330
rect 65834 22278 65846 22330
rect 65898 22278 65910 22330
rect 65962 22278 96374 22330
rect 96426 22278 96438 22330
rect 96490 22278 96502 22330
rect 96554 22278 96566 22330
rect 96618 22278 96630 22330
rect 96682 22278 127094 22330
rect 127146 22278 127158 22330
rect 127210 22278 127222 22330
rect 127274 22278 127286 22330
rect 127338 22278 127350 22330
rect 127402 22278 148856 22330
rect 1104 22256 148856 22278
rect 1104 21786 148856 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 81014 21786
rect 81066 21734 81078 21786
rect 81130 21734 81142 21786
rect 81194 21734 81206 21786
rect 81258 21734 81270 21786
rect 81322 21734 111734 21786
rect 111786 21734 111798 21786
rect 111850 21734 111862 21786
rect 111914 21734 111926 21786
rect 111978 21734 111990 21786
rect 112042 21734 142454 21786
rect 142506 21734 142518 21786
rect 142570 21734 142582 21786
rect 142634 21734 142646 21786
rect 142698 21734 142710 21786
rect 142762 21734 148856 21786
rect 1104 21712 148856 21734
rect 1104 21242 148856 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 65654 21242
rect 65706 21190 65718 21242
rect 65770 21190 65782 21242
rect 65834 21190 65846 21242
rect 65898 21190 65910 21242
rect 65962 21190 96374 21242
rect 96426 21190 96438 21242
rect 96490 21190 96502 21242
rect 96554 21190 96566 21242
rect 96618 21190 96630 21242
rect 96682 21190 127094 21242
rect 127146 21190 127158 21242
rect 127210 21190 127222 21242
rect 127274 21190 127286 21242
rect 127338 21190 127350 21242
rect 127402 21190 148856 21242
rect 1104 21168 148856 21190
rect 1104 20698 148856 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 81014 20698
rect 81066 20646 81078 20698
rect 81130 20646 81142 20698
rect 81194 20646 81206 20698
rect 81258 20646 81270 20698
rect 81322 20646 111734 20698
rect 111786 20646 111798 20698
rect 111850 20646 111862 20698
rect 111914 20646 111926 20698
rect 111978 20646 111990 20698
rect 112042 20646 142454 20698
rect 142506 20646 142518 20698
rect 142570 20646 142582 20698
rect 142634 20646 142646 20698
rect 142698 20646 142710 20698
rect 142762 20646 148856 20698
rect 1104 20624 148856 20646
rect 1104 20154 148856 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 65654 20154
rect 65706 20102 65718 20154
rect 65770 20102 65782 20154
rect 65834 20102 65846 20154
rect 65898 20102 65910 20154
rect 65962 20102 96374 20154
rect 96426 20102 96438 20154
rect 96490 20102 96502 20154
rect 96554 20102 96566 20154
rect 96618 20102 96630 20154
rect 96682 20102 127094 20154
rect 127146 20102 127158 20154
rect 127210 20102 127222 20154
rect 127274 20102 127286 20154
rect 127338 20102 127350 20154
rect 127402 20102 148856 20154
rect 1104 20080 148856 20102
rect 1104 19610 148856 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 81014 19610
rect 81066 19558 81078 19610
rect 81130 19558 81142 19610
rect 81194 19558 81206 19610
rect 81258 19558 81270 19610
rect 81322 19558 111734 19610
rect 111786 19558 111798 19610
rect 111850 19558 111862 19610
rect 111914 19558 111926 19610
rect 111978 19558 111990 19610
rect 112042 19558 142454 19610
rect 142506 19558 142518 19610
rect 142570 19558 142582 19610
rect 142634 19558 142646 19610
rect 142698 19558 142710 19610
rect 142762 19558 148856 19610
rect 1104 19536 148856 19558
rect 1104 19066 148856 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 65654 19066
rect 65706 19014 65718 19066
rect 65770 19014 65782 19066
rect 65834 19014 65846 19066
rect 65898 19014 65910 19066
rect 65962 19014 96374 19066
rect 96426 19014 96438 19066
rect 96490 19014 96502 19066
rect 96554 19014 96566 19066
rect 96618 19014 96630 19066
rect 96682 19014 127094 19066
rect 127146 19014 127158 19066
rect 127210 19014 127222 19066
rect 127274 19014 127286 19066
rect 127338 19014 127350 19066
rect 127402 19014 148856 19066
rect 1104 18992 148856 19014
rect 1104 18522 148856 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 81014 18522
rect 81066 18470 81078 18522
rect 81130 18470 81142 18522
rect 81194 18470 81206 18522
rect 81258 18470 81270 18522
rect 81322 18470 111734 18522
rect 111786 18470 111798 18522
rect 111850 18470 111862 18522
rect 111914 18470 111926 18522
rect 111978 18470 111990 18522
rect 112042 18470 142454 18522
rect 142506 18470 142518 18522
rect 142570 18470 142582 18522
rect 142634 18470 142646 18522
rect 142698 18470 142710 18522
rect 142762 18470 148856 18522
rect 1104 18448 148856 18470
rect 1104 17978 148856 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 65654 17978
rect 65706 17926 65718 17978
rect 65770 17926 65782 17978
rect 65834 17926 65846 17978
rect 65898 17926 65910 17978
rect 65962 17926 96374 17978
rect 96426 17926 96438 17978
rect 96490 17926 96502 17978
rect 96554 17926 96566 17978
rect 96618 17926 96630 17978
rect 96682 17926 127094 17978
rect 127146 17926 127158 17978
rect 127210 17926 127222 17978
rect 127274 17926 127286 17978
rect 127338 17926 127350 17978
rect 127402 17926 148856 17978
rect 1104 17904 148856 17926
rect 1104 17434 148856 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 81014 17434
rect 81066 17382 81078 17434
rect 81130 17382 81142 17434
rect 81194 17382 81206 17434
rect 81258 17382 81270 17434
rect 81322 17382 111734 17434
rect 111786 17382 111798 17434
rect 111850 17382 111862 17434
rect 111914 17382 111926 17434
rect 111978 17382 111990 17434
rect 112042 17382 142454 17434
rect 142506 17382 142518 17434
rect 142570 17382 142582 17434
rect 142634 17382 142646 17434
rect 142698 17382 142710 17434
rect 142762 17382 148856 17434
rect 1104 17360 148856 17382
rect 1104 16890 148856 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 65654 16890
rect 65706 16838 65718 16890
rect 65770 16838 65782 16890
rect 65834 16838 65846 16890
rect 65898 16838 65910 16890
rect 65962 16838 96374 16890
rect 96426 16838 96438 16890
rect 96490 16838 96502 16890
rect 96554 16838 96566 16890
rect 96618 16838 96630 16890
rect 96682 16838 127094 16890
rect 127146 16838 127158 16890
rect 127210 16838 127222 16890
rect 127274 16838 127286 16890
rect 127338 16838 127350 16890
rect 127402 16838 148856 16890
rect 1104 16816 148856 16838
rect 1104 16346 148856 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 81014 16346
rect 81066 16294 81078 16346
rect 81130 16294 81142 16346
rect 81194 16294 81206 16346
rect 81258 16294 81270 16346
rect 81322 16294 111734 16346
rect 111786 16294 111798 16346
rect 111850 16294 111862 16346
rect 111914 16294 111926 16346
rect 111978 16294 111990 16346
rect 112042 16294 142454 16346
rect 142506 16294 142518 16346
rect 142570 16294 142582 16346
rect 142634 16294 142646 16346
rect 142698 16294 142710 16346
rect 142762 16294 148856 16346
rect 1104 16272 148856 16294
rect 1104 15802 148856 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 65654 15802
rect 65706 15750 65718 15802
rect 65770 15750 65782 15802
rect 65834 15750 65846 15802
rect 65898 15750 65910 15802
rect 65962 15750 96374 15802
rect 96426 15750 96438 15802
rect 96490 15750 96502 15802
rect 96554 15750 96566 15802
rect 96618 15750 96630 15802
rect 96682 15750 127094 15802
rect 127146 15750 127158 15802
rect 127210 15750 127222 15802
rect 127274 15750 127286 15802
rect 127338 15750 127350 15802
rect 127402 15750 148856 15802
rect 1104 15728 148856 15750
rect 1104 15258 148856 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 81014 15258
rect 81066 15206 81078 15258
rect 81130 15206 81142 15258
rect 81194 15206 81206 15258
rect 81258 15206 81270 15258
rect 81322 15206 111734 15258
rect 111786 15206 111798 15258
rect 111850 15206 111862 15258
rect 111914 15206 111926 15258
rect 111978 15206 111990 15258
rect 112042 15206 142454 15258
rect 142506 15206 142518 15258
rect 142570 15206 142582 15258
rect 142634 15206 142646 15258
rect 142698 15206 142710 15258
rect 142762 15206 148856 15258
rect 1104 15184 148856 15206
rect 1104 14714 148856 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 65654 14714
rect 65706 14662 65718 14714
rect 65770 14662 65782 14714
rect 65834 14662 65846 14714
rect 65898 14662 65910 14714
rect 65962 14662 96374 14714
rect 96426 14662 96438 14714
rect 96490 14662 96502 14714
rect 96554 14662 96566 14714
rect 96618 14662 96630 14714
rect 96682 14662 127094 14714
rect 127146 14662 127158 14714
rect 127210 14662 127222 14714
rect 127274 14662 127286 14714
rect 127338 14662 127350 14714
rect 127402 14662 148856 14714
rect 1104 14640 148856 14662
rect 1104 14170 148856 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 81014 14170
rect 81066 14118 81078 14170
rect 81130 14118 81142 14170
rect 81194 14118 81206 14170
rect 81258 14118 81270 14170
rect 81322 14118 111734 14170
rect 111786 14118 111798 14170
rect 111850 14118 111862 14170
rect 111914 14118 111926 14170
rect 111978 14118 111990 14170
rect 112042 14118 142454 14170
rect 142506 14118 142518 14170
rect 142570 14118 142582 14170
rect 142634 14118 142646 14170
rect 142698 14118 142710 14170
rect 142762 14118 148856 14170
rect 1104 14096 148856 14118
rect 1104 13626 148856 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 65654 13626
rect 65706 13574 65718 13626
rect 65770 13574 65782 13626
rect 65834 13574 65846 13626
rect 65898 13574 65910 13626
rect 65962 13574 96374 13626
rect 96426 13574 96438 13626
rect 96490 13574 96502 13626
rect 96554 13574 96566 13626
rect 96618 13574 96630 13626
rect 96682 13574 127094 13626
rect 127146 13574 127158 13626
rect 127210 13574 127222 13626
rect 127274 13574 127286 13626
rect 127338 13574 127350 13626
rect 127402 13574 148856 13626
rect 1104 13552 148856 13574
rect 1104 13082 148856 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 81014 13082
rect 81066 13030 81078 13082
rect 81130 13030 81142 13082
rect 81194 13030 81206 13082
rect 81258 13030 81270 13082
rect 81322 13030 111734 13082
rect 111786 13030 111798 13082
rect 111850 13030 111862 13082
rect 111914 13030 111926 13082
rect 111978 13030 111990 13082
rect 112042 13030 142454 13082
rect 142506 13030 142518 13082
rect 142570 13030 142582 13082
rect 142634 13030 142646 13082
rect 142698 13030 142710 13082
rect 142762 13030 148856 13082
rect 1104 13008 148856 13030
rect 1104 12538 148856 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 65654 12538
rect 65706 12486 65718 12538
rect 65770 12486 65782 12538
rect 65834 12486 65846 12538
rect 65898 12486 65910 12538
rect 65962 12486 96374 12538
rect 96426 12486 96438 12538
rect 96490 12486 96502 12538
rect 96554 12486 96566 12538
rect 96618 12486 96630 12538
rect 96682 12486 127094 12538
rect 127146 12486 127158 12538
rect 127210 12486 127222 12538
rect 127274 12486 127286 12538
rect 127338 12486 127350 12538
rect 127402 12486 148856 12538
rect 1104 12464 148856 12486
rect 9582 12248 9588 12300
rect 9640 12288 9646 12300
rect 15378 12288 15384 12300
rect 9640 12260 15384 12288
rect 9640 12248 9646 12260
rect 15378 12248 15384 12260
rect 15436 12248 15442 12300
rect 1104 11994 148856 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 81014 11994
rect 81066 11942 81078 11994
rect 81130 11942 81142 11994
rect 81194 11942 81206 11994
rect 81258 11942 81270 11994
rect 81322 11942 111734 11994
rect 111786 11942 111798 11994
rect 111850 11942 111862 11994
rect 111914 11942 111926 11994
rect 111978 11942 111990 11994
rect 112042 11942 142454 11994
rect 142506 11942 142518 11994
rect 142570 11942 142582 11994
rect 142634 11942 142646 11994
rect 142698 11942 142710 11994
rect 142762 11942 148856 11994
rect 1104 11920 148856 11942
rect 1104 11450 148856 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 65654 11450
rect 65706 11398 65718 11450
rect 65770 11398 65782 11450
rect 65834 11398 65846 11450
rect 65898 11398 65910 11450
rect 65962 11398 96374 11450
rect 96426 11398 96438 11450
rect 96490 11398 96502 11450
rect 96554 11398 96566 11450
rect 96618 11398 96630 11450
rect 96682 11398 127094 11450
rect 127146 11398 127158 11450
rect 127210 11398 127222 11450
rect 127274 11398 127286 11450
rect 127338 11398 127350 11450
rect 127402 11398 148856 11450
rect 1104 11376 148856 11398
rect 1104 10906 148856 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 81014 10906
rect 81066 10854 81078 10906
rect 81130 10854 81142 10906
rect 81194 10854 81206 10906
rect 81258 10854 81270 10906
rect 81322 10854 111734 10906
rect 111786 10854 111798 10906
rect 111850 10854 111862 10906
rect 111914 10854 111926 10906
rect 111978 10854 111990 10906
rect 112042 10854 142454 10906
rect 142506 10854 142518 10906
rect 142570 10854 142582 10906
rect 142634 10854 142646 10906
rect 142698 10854 142710 10906
rect 142762 10854 148856 10906
rect 1104 10832 148856 10854
rect 1104 10362 148856 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 65654 10362
rect 65706 10310 65718 10362
rect 65770 10310 65782 10362
rect 65834 10310 65846 10362
rect 65898 10310 65910 10362
rect 65962 10310 96374 10362
rect 96426 10310 96438 10362
rect 96490 10310 96502 10362
rect 96554 10310 96566 10362
rect 96618 10310 96630 10362
rect 96682 10310 127094 10362
rect 127146 10310 127158 10362
rect 127210 10310 127222 10362
rect 127274 10310 127286 10362
rect 127338 10310 127350 10362
rect 127402 10310 148856 10362
rect 1104 10288 148856 10310
rect 1104 9818 148856 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 81014 9818
rect 81066 9766 81078 9818
rect 81130 9766 81142 9818
rect 81194 9766 81206 9818
rect 81258 9766 81270 9818
rect 81322 9766 111734 9818
rect 111786 9766 111798 9818
rect 111850 9766 111862 9818
rect 111914 9766 111926 9818
rect 111978 9766 111990 9818
rect 112042 9766 142454 9818
rect 142506 9766 142518 9818
rect 142570 9766 142582 9818
rect 142634 9766 142646 9818
rect 142698 9766 142710 9818
rect 142762 9766 148856 9818
rect 1104 9744 148856 9766
rect 1104 9274 148856 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 65654 9274
rect 65706 9222 65718 9274
rect 65770 9222 65782 9274
rect 65834 9222 65846 9274
rect 65898 9222 65910 9274
rect 65962 9222 96374 9274
rect 96426 9222 96438 9274
rect 96490 9222 96502 9274
rect 96554 9222 96566 9274
rect 96618 9222 96630 9274
rect 96682 9222 127094 9274
rect 127146 9222 127158 9274
rect 127210 9222 127222 9274
rect 127274 9222 127286 9274
rect 127338 9222 127350 9274
rect 127402 9222 148856 9274
rect 1104 9200 148856 9222
rect 1104 8730 148856 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 81014 8730
rect 81066 8678 81078 8730
rect 81130 8678 81142 8730
rect 81194 8678 81206 8730
rect 81258 8678 81270 8730
rect 81322 8678 111734 8730
rect 111786 8678 111798 8730
rect 111850 8678 111862 8730
rect 111914 8678 111926 8730
rect 111978 8678 111990 8730
rect 112042 8678 142454 8730
rect 142506 8678 142518 8730
rect 142570 8678 142582 8730
rect 142634 8678 142646 8730
rect 142698 8678 142710 8730
rect 142762 8678 148856 8730
rect 1104 8656 148856 8678
rect 66806 8304 66812 8356
rect 66864 8344 66870 8356
rect 67634 8344 67640 8356
rect 66864 8316 67640 8344
rect 66864 8304 66870 8316
rect 67634 8304 67640 8316
rect 67692 8304 67698 8356
rect 1104 8186 148856 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 65654 8186
rect 65706 8134 65718 8186
rect 65770 8134 65782 8186
rect 65834 8134 65846 8186
rect 65898 8134 65910 8186
rect 65962 8134 96374 8186
rect 96426 8134 96438 8186
rect 96490 8134 96502 8186
rect 96554 8134 96566 8186
rect 96618 8134 96630 8186
rect 96682 8134 127094 8186
rect 127146 8134 127158 8186
rect 127210 8134 127222 8186
rect 127274 8134 127286 8186
rect 127338 8134 127350 8186
rect 127402 8134 148856 8186
rect 1104 8112 148856 8134
rect 1104 7642 148856 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 81014 7642
rect 81066 7590 81078 7642
rect 81130 7590 81142 7642
rect 81194 7590 81206 7642
rect 81258 7590 81270 7642
rect 81322 7590 111734 7642
rect 111786 7590 111798 7642
rect 111850 7590 111862 7642
rect 111914 7590 111926 7642
rect 111978 7590 111990 7642
rect 112042 7590 142454 7642
rect 142506 7590 142518 7642
rect 142570 7590 142582 7642
rect 142634 7590 142646 7642
rect 142698 7590 142710 7642
rect 142762 7590 148856 7642
rect 1104 7568 148856 7590
rect 1104 7098 148856 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 65654 7098
rect 65706 7046 65718 7098
rect 65770 7046 65782 7098
rect 65834 7046 65846 7098
rect 65898 7046 65910 7098
rect 65962 7046 96374 7098
rect 96426 7046 96438 7098
rect 96490 7046 96502 7098
rect 96554 7046 96566 7098
rect 96618 7046 96630 7098
rect 96682 7046 127094 7098
rect 127146 7046 127158 7098
rect 127210 7046 127222 7098
rect 127274 7046 127286 7098
rect 127338 7046 127350 7098
rect 127402 7046 148856 7098
rect 1104 7024 148856 7046
rect 82446 6808 82452 6860
rect 82504 6848 82510 6860
rect 83090 6848 83096 6860
rect 82504 6820 83096 6848
rect 82504 6808 82510 6820
rect 83090 6808 83096 6820
rect 83148 6808 83154 6860
rect 1104 6554 148856 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 81014 6554
rect 81066 6502 81078 6554
rect 81130 6502 81142 6554
rect 81194 6502 81206 6554
rect 81258 6502 81270 6554
rect 81322 6502 111734 6554
rect 111786 6502 111798 6554
rect 111850 6502 111862 6554
rect 111914 6502 111926 6554
rect 111978 6502 111990 6554
rect 112042 6502 142454 6554
rect 142506 6502 142518 6554
rect 142570 6502 142582 6554
rect 142634 6502 142646 6554
rect 142698 6502 142710 6554
rect 142762 6502 148856 6554
rect 1104 6480 148856 6502
rect 1104 6010 148856 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 65654 6010
rect 65706 5958 65718 6010
rect 65770 5958 65782 6010
rect 65834 5958 65846 6010
rect 65898 5958 65910 6010
rect 65962 5958 96374 6010
rect 96426 5958 96438 6010
rect 96490 5958 96502 6010
rect 96554 5958 96566 6010
rect 96618 5958 96630 6010
rect 96682 5958 127094 6010
rect 127146 5958 127158 6010
rect 127210 5958 127222 6010
rect 127274 5958 127286 6010
rect 127338 5958 127350 6010
rect 127402 5958 148856 6010
rect 1104 5936 148856 5958
rect 64046 5896 64052 5908
rect 64007 5868 64052 5896
rect 64046 5856 64052 5868
rect 64104 5856 64110 5908
rect 65518 5856 65524 5908
rect 65576 5896 65582 5908
rect 65797 5899 65855 5905
rect 65797 5896 65809 5899
rect 65576 5868 65809 5896
rect 65576 5856 65582 5868
rect 65797 5865 65809 5868
rect 65843 5865 65855 5899
rect 65797 5859 65855 5865
rect 80054 5856 80060 5908
rect 80112 5896 80118 5908
rect 80112 5868 80157 5896
rect 80112 5856 80118 5868
rect 78214 5652 78220 5704
rect 78272 5692 78278 5704
rect 79042 5692 79048 5704
rect 78272 5664 79048 5692
rect 78272 5652 78278 5664
rect 79042 5652 79048 5664
rect 79100 5652 79106 5704
rect 65150 5556 65156 5568
rect 65111 5528 65156 5556
rect 65150 5516 65156 5528
rect 65208 5516 65214 5568
rect 69474 5556 69480 5568
rect 69435 5528 69480 5556
rect 69474 5516 69480 5528
rect 69532 5516 69538 5568
rect 75730 5516 75736 5568
rect 75788 5556 75794 5568
rect 76466 5556 76472 5568
rect 75788 5528 76472 5556
rect 75788 5516 75794 5528
rect 76466 5516 76472 5528
rect 76524 5516 76530 5568
rect 77202 5516 77208 5568
rect 77260 5556 77266 5568
rect 78490 5556 78496 5568
rect 77260 5528 78496 5556
rect 77260 5516 77266 5528
rect 78490 5516 78496 5528
rect 78548 5516 78554 5568
rect 79045 5559 79103 5565
rect 79045 5525 79057 5559
rect 79091 5556 79103 5559
rect 79134 5556 79140 5568
rect 79091 5528 79140 5556
rect 79091 5525 79103 5528
rect 79045 5519 79103 5525
rect 79134 5516 79140 5528
rect 79192 5556 79198 5568
rect 79505 5559 79563 5565
rect 79505 5556 79517 5559
rect 79192 5528 79517 5556
rect 79192 5516 79198 5528
rect 79505 5525 79517 5528
rect 79551 5525 79563 5559
rect 79505 5519 79563 5525
rect 80146 5516 80152 5568
rect 80204 5556 80210 5568
rect 80609 5559 80667 5565
rect 80609 5556 80621 5559
rect 80204 5528 80621 5556
rect 80204 5516 80210 5528
rect 80609 5525 80621 5528
rect 80655 5525 80667 5559
rect 80609 5519 80667 5525
rect 1104 5466 148856 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 81014 5466
rect 81066 5414 81078 5466
rect 81130 5414 81142 5466
rect 81194 5414 81206 5466
rect 81258 5414 81270 5466
rect 81322 5414 111734 5466
rect 111786 5414 111798 5466
rect 111850 5414 111862 5466
rect 111914 5414 111926 5466
rect 111978 5414 111990 5466
rect 112042 5414 142454 5466
rect 142506 5414 142518 5466
rect 142570 5414 142582 5466
rect 142634 5414 142646 5466
rect 142698 5414 142710 5466
rect 142762 5414 148856 5466
rect 1104 5392 148856 5414
rect 28350 5352 28356 5364
rect 28311 5324 28356 5352
rect 28350 5312 28356 5324
rect 28408 5312 28414 5364
rect 36078 5352 36084 5364
rect 36039 5324 36084 5352
rect 36078 5312 36084 5324
rect 36136 5312 36142 5364
rect 38194 5312 38200 5364
rect 38252 5352 38258 5364
rect 38289 5355 38347 5361
rect 38289 5352 38301 5355
rect 38252 5324 38301 5352
rect 38252 5312 38258 5324
rect 38289 5321 38301 5324
rect 38335 5321 38347 5355
rect 38289 5315 38347 5321
rect 52086 5312 52092 5364
rect 52144 5352 52150 5364
rect 52362 5352 52368 5364
rect 52144 5324 52368 5352
rect 52144 5312 52150 5324
rect 52362 5312 52368 5324
rect 52420 5352 52426 5364
rect 53469 5355 53527 5361
rect 53469 5352 53481 5355
rect 52420 5324 53481 5352
rect 52420 5312 52426 5324
rect 53469 5321 53481 5324
rect 53515 5321 53527 5355
rect 53469 5315 53527 5321
rect 63494 5312 63500 5364
rect 63552 5352 63558 5364
rect 63681 5355 63739 5361
rect 63681 5352 63693 5355
rect 63552 5324 63693 5352
rect 63552 5312 63558 5324
rect 63681 5321 63693 5324
rect 63727 5321 63739 5355
rect 63681 5315 63739 5321
rect 65981 5355 66039 5361
rect 65981 5321 65993 5355
rect 66027 5352 66039 5355
rect 66070 5352 66076 5364
rect 66027 5324 66076 5352
rect 66027 5321 66039 5324
rect 65981 5315 66039 5321
rect 66070 5312 66076 5324
rect 66128 5312 66134 5364
rect 69017 5355 69075 5361
rect 69017 5321 69029 5355
rect 69063 5352 69075 5355
rect 69106 5352 69112 5364
rect 69063 5324 69112 5352
rect 69063 5321 69075 5324
rect 69017 5315 69075 5321
rect 69106 5312 69112 5324
rect 69164 5312 69170 5364
rect 69474 5312 69480 5364
rect 69532 5352 69538 5364
rect 69661 5355 69719 5361
rect 69661 5352 69673 5355
rect 69532 5324 69673 5352
rect 69532 5312 69538 5324
rect 69661 5321 69673 5324
rect 69707 5352 69719 5355
rect 78769 5355 78827 5361
rect 78769 5352 78781 5355
rect 69707 5324 78781 5352
rect 69707 5321 69719 5324
rect 69661 5315 69719 5321
rect 78769 5321 78781 5324
rect 78815 5321 78827 5355
rect 78769 5315 78827 5321
rect 67085 5287 67143 5293
rect 67085 5253 67097 5287
rect 67131 5284 67143 5287
rect 68186 5284 68192 5296
rect 67131 5256 68192 5284
rect 67131 5253 67143 5256
rect 67085 5247 67143 5253
rect 68186 5244 68192 5256
rect 68244 5284 68250 5296
rect 69492 5284 69520 5312
rect 68244 5256 69520 5284
rect 68244 5244 68250 5256
rect 78784 5216 78812 5315
rect 79336 5256 81480 5284
rect 79336 5225 79364 5256
rect 81452 5225 81480 5256
rect 79321 5219 79379 5225
rect 79321 5216 79333 5219
rect 78784 5188 79333 5216
rect 79321 5185 79333 5188
rect 79367 5185 79379 5219
rect 79321 5179 79379 5185
rect 80149 5219 80207 5225
rect 80149 5185 80161 5219
rect 80195 5185 80207 5219
rect 80149 5179 80207 5185
rect 80793 5219 80851 5225
rect 80793 5185 80805 5219
rect 80839 5185 80851 5219
rect 80793 5179 80851 5185
rect 81437 5219 81495 5225
rect 81437 5185 81449 5219
rect 81483 5216 81495 5219
rect 81483 5188 82032 5216
rect 81483 5185 81495 5188
rect 81437 5179 81495 5185
rect 36740 5120 41414 5148
rect 34790 5040 34796 5092
rect 34848 5080 34854 5092
rect 36740 5089 36768 5120
rect 36725 5083 36783 5089
rect 36725 5080 36737 5083
rect 34848 5052 36737 5080
rect 34848 5040 34854 5052
rect 36725 5049 36737 5052
rect 36771 5049 36783 5083
rect 36725 5043 36783 5049
rect 37553 5083 37611 5089
rect 37553 5049 37565 5083
rect 37599 5080 37611 5083
rect 38562 5080 38568 5092
rect 37599 5052 38568 5080
rect 37599 5049 37611 5052
rect 37553 5043 37611 5049
rect 38562 5040 38568 5052
rect 38620 5040 38626 5092
rect 35618 5012 35624 5024
rect 35579 4984 35624 5012
rect 35618 4972 35624 4984
rect 35676 4972 35682 5024
rect 41386 5012 41414 5120
rect 60826 5080 60832 5092
rect 60739 5052 60832 5080
rect 60826 5040 60832 5052
rect 60884 5080 60890 5092
rect 62577 5083 62635 5089
rect 62577 5080 62589 5083
rect 60884 5052 62589 5080
rect 60884 5040 60890 5052
rect 62577 5049 62589 5052
rect 62623 5049 62635 5083
rect 62577 5043 62635 5049
rect 66533 5083 66591 5089
rect 66533 5049 66545 5083
rect 66579 5080 66591 5083
rect 78125 5083 78183 5089
rect 66579 5052 70394 5080
rect 66579 5049 66591 5052
rect 66533 5043 66591 5049
rect 70366 5024 70394 5052
rect 78125 5049 78137 5083
rect 78171 5080 78183 5083
rect 79134 5080 79140 5092
rect 78171 5052 79140 5080
rect 78171 5049 78183 5052
rect 78125 5043 78183 5049
rect 79134 5040 79140 5052
rect 79192 5040 79198 5092
rect 80164 5080 80192 5179
rect 80808 5148 80836 5179
rect 81710 5148 81716 5160
rect 80808 5120 81716 5148
rect 81710 5108 81716 5120
rect 81768 5108 81774 5160
rect 81434 5080 81440 5092
rect 80164 5052 81440 5080
rect 81434 5040 81440 5052
rect 81492 5040 81498 5092
rect 82004 5024 82032 5188
rect 82541 5083 82599 5089
rect 82541 5049 82553 5083
rect 82587 5080 82599 5083
rect 83366 5080 83372 5092
rect 82587 5052 83372 5080
rect 82587 5049 82599 5052
rect 82541 5043 82599 5049
rect 83366 5040 83372 5052
rect 83424 5040 83430 5092
rect 42702 5012 42708 5024
rect 41386 4984 42708 5012
rect 42702 4972 42708 4984
rect 42760 4972 42766 5024
rect 47118 5012 47124 5024
rect 47079 4984 47124 5012
rect 47118 4972 47124 4984
rect 47176 4972 47182 5024
rect 48130 5012 48136 5024
rect 48091 4984 48136 5012
rect 48130 4972 48136 4984
rect 48188 4972 48194 5024
rect 48314 4972 48320 5024
rect 48372 5012 48378 5024
rect 48593 5015 48651 5021
rect 48593 5012 48605 5015
rect 48372 4984 48605 5012
rect 48372 4972 48378 4984
rect 48593 4981 48605 4984
rect 48639 4981 48651 5015
rect 48593 4975 48651 4981
rect 49050 4972 49056 5024
rect 49108 5012 49114 5024
rect 49145 5015 49203 5021
rect 49145 5012 49157 5015
rect 49108 4984 49157 5012
rect 49108 4972 49114 4984
rect 49145 4981 49157 4984
rect 49191 5012 49203 5015
rect 49602 5012 49608 5024
rect 49191 4984 49608 5012
rect 49191 4981 49203 4984
rect 49145 4975 49203 4981
rect 49602 4972 49608 4984
rect 49660 4972 49666 5024
rect 53006 5012 53012 5024
rect 52967 4984 53012 5012
rect 53006 4972 53012 4984
rect 53064 4972 53070 5024
rect 58066 5012 58072 5024
rect 58027 4984 58072 5012
rect 58066 4972 58072 4984
rect 58124 4972 58130 5024
rect 58710 5012 58716 5024
rect 58671 4984 58716 5012
rect 58710 4972 58716 4984
rect 58768 4972 58774 5024
rect 61838 5012 61844 5024
rect 61799 4984 61844 5012
rect 61838 4972 61844 4984
rect 61896 4972 61902 5024
rect 64322 5012 64328 5024
rect 64283 4984 64328 5012
rect 64322 4972 64328 4984
rect 64380 4972 64386 5024
rect 64874 5012 64880 5024
rect 64835 4984 64880 5012
rect 64874 4972 64880 4984
rect 64932 4972 64938 5024
rect 65334 5012 65340 5024
rect 65295 4984 65340 5012
rect 65334 4972 65340 4984
rect 65392 4972 65398 5024
rect 68465 5015 68523 5021
rect 68465 4981 68477 5015
rect 68511 5012 68523 5015
rect 68922 5012 68928 5024
rect 68511 4984 68928 5012
rect 68511 4981 68523 4984
rect 68465 4975 68523 4981
rect 68922 4972 68928 4984
rect 68980 4972 68986 5024
rect 69658 4972 69664 5024
rect 69716 5012 69722 5024
rect 70121 5015 70179 5021
rect 70121 5012 70133 5015
rect 69716 4984 70133 5012
rect 69716 4972 69722 4984
rect 70121 4981 70133 4984
rect 70167 4981 70179 5015
rect 70121 4975 70179 4981
rect 70302 4972 70308 5024
rect 70360 5012 70394 5024
rect 70673 5015 70731 5021
rect 70673 5012 70685 5015
rect 70360 4984 70685 5012
rect 70360 4972 70366 4984
rect 70673 4981 70685 4984
rect 70719 4981 70731 5015
rect 79410 5012 79416 5024
rect 79371 4984 79416 5012
rect 70673 4975 70731 4981
rect 79410 4972 79416 4984
rect 79468 4972 79474 5024
rect 79502 4972 79508 5024
rect 79560 5012 79566 5024
rect 79965 5015 80023 5021
rect 79965 5012 79977 5015
rect 79560 4984 79977 5012
rect 79560 4972 79566 4984
rect 79965 4981 79977 4984
rect 80011 4981 80023 5015
rect 79965 4975 80023 4981
rect 80238 4972 80244 5024
rect 80296 5012 80302 5024
rect 80609 5015 80667 5021
rect 80609 5012 80621 5015
rect 80296 4984 80621 5012
rect 80296 4972 80302 4984
rect 80609 4981 80621 4984
rect 80655 4981 80667 5015
rect 80609 4975 80667 4981
rect 80790 4972 80796 5024
rect 80848 5012 80854 5024
rect 81345 5015 81403 5021
rect 81345 5012 81357 5015
rect 80848 4984 81357 5012
rect 80848 4972 80854 4984
rect 81345 4981 81357 4984
rect 81391 4981 81403 5015
rect 81986 5012 81992 5024
rect 81947 4984 81992 5012
rect 81345 4975 81403 4981
rect 81986 4972 81992 4984
rect 82044 4972 82050 5024
rect 82998 5012 83004 5024
rect 82959 4984 83004 5012
rect 82998 4972 83004 4984
rect 83056 4972 83062 5024
rect 1104 4922 148856 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 65654 4922
rect 65706 4870 65718 4922
rect 65770 4870 65782 4922
rect 65834 4870 65846 4922
rect 65898 4870 65910 4922
rect 65962 4870 96374 4922
rect 96426 4870 96438 4922
rect 96490 4870 96502 4922
rect 96554 4870 96566 4922
rect 96618 4870 96630 4922
rect 96682 4870 127094 4922
rect 127146 4870 127158 4922
rect 127210 4870 127222 4922
rect 127274 4870 127286 4922
rect 127338 4870 127350 4922
rect 127402 4870 148856 4922
rect 1104 4848 148856 4870
rect 40586 4808 40592 4820
rect 40547 4780 40592 4808
rect 40586 4768 40592 4780
rect 40644 4768 40650 4820
rect 42702 4768 42708 4820
rect 42760 4808 42766 4820
rect 45281 4811 45339 4817
rect 45281 4808 45293 4811
rect 42760 4780 45293 4808
rect 42760 4768 42766 4780
rect 45281 4777 45293 4780
rect 45327 4777 45339 4811
rect 45281 4771 45339 4777
rect 48317 4811 48375 4817
rect 48317 4777 48329 4811
rect 48363 4808 48375 4811
rect 48590 4808 48596 4820
rect 48363 4780 48596 4808
rect 48363 4777 48375 4780
rect 48317 4771 48375 4777
rect 48590 4768 48596 4780
rect 48648 4768 48654 4820
rect 48958 4808 48964 4820
rect 48919 4780 48964 4808
rect 48958 4768 48964 4780
rect 49016 4768 49022 4820
rect 49510 4808 49516 4820
rect 49471 4780 49516 4808
rect 49510 4768 49516 4780
rect 49568 4768 49574 4820
rect 53834 4808 53840 4820
rect 53795 4780 53840 4808
rect 53834 4768 53840 4780
rect 53892 4768 53898 4820
rect 57974 4808 57980 4820
rect 57887 4780 57980 4808
rect 57974 4768 57980 4780
rect 58032 4808 58038 4820
rect 58618 4808 58624 4820
rect 58032 4780 58624 4808
rect 58032 4768 58038 4780
rect 58618 4768 58624 4780
rect 58676 4768 58682 4820
rect 59078 4808 59084 4820
rect 59039 4780 59084 4808
rect 59078 4768 59084 4780
rect 59136 4768 59142 4820
rect 61102 4808 61108 4820
rect 61063 4780 61108 4808
rect 61102 4768 61108 4780
rect 61160 4768 61166 4820
rect 67634 4808 67640 4820
rect 67595 4780 67640 4808
rect 67634 4768 67640 4780
rect 67692 4768 67698 4820
rect 68186 4808 68192 4820
rect 68147 4780 68192 4808
rect 68186 4768 68192 4780
rect 68244 4768 68250 4820
rect 78214 4808 78220 4820
rect 78175 4780 78220 4808
rect 78214 4768 78220 4780
rect 78272 4768 78278 4820
rect 83090 4808 83096 4820
rect 83051 4780 83096 4808
rect 83090 4768 83096 4780
rect 83148 4768 83154 4820
rect 43438 4740 43444 4752
rect 43399 4712 43444 4740
rect 43438 4700 43444 4712
rect 43496 4700 43502 4752
rect 49528 4740 49556 4768
rect 47504 4712 49556 4740
rect 33689 4675 33747 4681
rect 33689 4641 33701 4675
rect 33735 4672 33747 4675
rect 34333 4675 34391 4681
rect 34333 4672 34345 4675
rect 33735 4644 34345 4672
rect 33735 4641 33747 4644
rect 33689 4635 33747 4641
rect 34333 4641 34345 4644
rect 34379 4672 34391 4675
rect 36906 4672 36912 4684
rect 34379 4644 36912 4672
rect 34379 4641 34391 4644
rect 34333 4635 34391 4641
rect 36906 4632 36912 4644
rect 36964 4632 36970 4684
rect 47504 4681 47532 4712
rect 49602 4700 49608 4752
rect 49660 4740 49666 4752
rect 66073 4743 66131 4749
rect 66073 4740 66085 4743
rect 49660 4712 66085 4740
rect 49660 4700 49666 4712
rect 66073 4709 66085 4712
rect 66119 4740 66131 4743
rect 66162 4740 66168 4752
rect 66119 4712 66168 4740
rect 66119 4709 66131 4712
rect 66073 4703 66131 4709
rect 66162 4700 66168 4712
rect 66220 4700 66226 4752
rect 66530 4700 66536 4752
rect 66588 4740 66594 4752
rect 66717 4743 66775 4749
rect 66717 4740 66729 4743
rect 66588 4712 66729 4740
rect 66588 4700 66594 4712
rect 66717 4709 66729 4712
rect 66763 4740 66775 4743
rect 68204 4740 68232 4768
rect 66763 4712 68232 4740
rect 80609 4743 80667 4749
rect 66763 4709 66775 4712
rect 66717 4703 66775 4709
rect 80609 4709 80621 4743
rect 80655 4740 80667 4743
rect 81526 4740 81532 4752
rect 80655 4712 81532 4740
rect 80655 4709 80667 4712
rect 80609 4703 80667 4709
rect 81526 4700 81532 4712
rect 81584 4700 81590 4752
rect 47489 4675 47547 4681
rect 47489 4641 47501 4675
rect 47535 4641 47547 4675
rect 47489 4635 47547 4641
rect 47578 4632 47584 4684
rect 47636 4672 47642 4684
rect 47636 4644 47681 4672
rect 47636 4632 47642 4644
rect 48130 4632 48136 4684
rect 48188 4672 48194 4684
rect 62945 4675 63003 4681
rect 62945 4672 62957 4675
rect 48188 4644 62957 4672
rect 48188 4632 48194 4644
rect 62945 4641 62957 4644
rect 62991 4672 63003 4675
rect 63310 4672 63316 4684
rect 62991 4644 63316 4672
rect 62991 4641 63003 4644
rect 62945 4635 63003 4641
rect 63310 4632 63316 4644
rect 63368 4632 63374 4684
rect 78674 4632 78680 4684
rect 78732 4672 78738 4684
rect 79778 4672 79784 4684
rect 78732 4644 79784 4672
rect 78732 4632 78738 4644
rect 79778 4632 79784 4644
rect 79836 4632 79842 4684
rect 81986 4672 81992 4684
rect 81452 4644 81992 4672
rect 26234 4564 26240 4616
rect 26292 4604 26298 4616
rect 28169 4607 28227 4613
rect 28169 4604 28181 4607
rect 26292 4576 28181 4604
rect 26292 4564 26298 4576
rect 28169 4573 28181 4576
rect 28215 4604 28227 4607
rect 29089 4607 29147 4613
rect 29089 4604 29101 4607
rect 28215 4576 29101 4604
rect 28215 4573 28227 4576
rect 28169 4567 28227 4573
rect 29089 4573 29101 4576
rect 29135 4604 29147 4607
rect 30282 4604 30288 4616
rect 29135 4576 30288 4604
rect 29135 4573 29147 4576
rect 29089 4567 29147 4573
rect 30282 4564 30288 4576
rect 30340 4564 30346 4616
rect 35345 4607 35403 4613
rect 35345 4573 35357 4607
rect 35391 4604 35403 4607
rect 35805 4607 35863 4613
rect 35805 4604 35817 4607
rect 35391 4576 35817 4604
rect 35391 4573 35403 4576
rect 35345 4567 35403 4573
rect 35805 4573 35817 4576
rect 35851 4604 35863 4607
rect 38010 4604 38016 4616
rect 35851 4576 38016 4604
rect 35851 4573 35863 4576
rect 35805 4567 35863 4573
rect 29733 4539 29791 4545
rect 29733 4536 29745 4539
rect 27632 4508 29745 4536
rect 27632 4480 27660 4508
rect 29733 4505 29745 4508
rect 29779 4505 29791 4539
rect 29733 4499 29791 4505
rect 33686 4496 33692 4548
rect 33744 4536 33750 4548
rect 35360 4536 35388 4567
rect 38010 4564 38016 4576
rect 38068 4604 38074 4616
rect 39850 4604 39856 4616
rect 38068 4576 39856 4604
rect 38068 4564 38074 4576
rect 39850 4564 39856 4576
rect 39908 4604 39914 4616
rect 40037 4607 40095 4613
rect 40037 4604 40049 4607
rect 39908 4576 40049 4604
rect 39908 4564 39914 4576
rect 40037 4573 40049 4576
rect 40083 4604 40095 4607
rect 41969 4607 42027 4613
rect 41969 4604 41981 4607
rect 40083 4576 41981 4604
rect 40083 4573 40095 4576
rect 40037 4567 40095 4573
rect 41969 4573 41981 4576
rect 42015 4604 42027 4607
rect 42426 4604 42432 4616
rect 42015 4576 42432 4604
rect 42015 4573 42027 4576
rect 41969 4567 42027 4573
rect 42426 4564 42432 4576
rect 42484 4564 42490 4616
rect 47210 4564 47216 4616
rect 47268 4604 47274 4616
rect 47397 4607 47455 4613
rect 47397 4604 47409 4607
rect 47268 4576 47409 4604
rect 47268 4564 47274 4576
rect 47397 4573 47409 4576
rect 47443 4604 47455 4607
rect 48148 4604 48176 4632
rect 47443 4576 48176 4604
rect 47443 4573 47455 4576
rect 47397 4567 47455 4573
rect 51442 4564 51448 4616
rect 51500 4604 51506 4616
rect 51629 4607 51687 4613
rect 51629 4604 51641 4607
rect 51500 4576 51641 4604
rect 51500 4564 51506 4576
rect 51629 4573 51641 4576
rect 51675 4573 51687 4607
rect 51629 4567 51687 4573
rect 57057 4607 57115 4613
rect 57057 4573 57069 4607
rect 57103 4604 57115 4607
rect 58158 4604 58164 4616
rect 57103 4576 58164 4604
rect 57103 4573 57115 4576
rect 57057 4567 57115 4573
rect 58158 4564 58164 4576
rect 58216 4564 58222 4616
rect 62206 4604 62212 4616
rect 62167 4576 62212 4604
rect 62206 4564 62212 4576
rect 62264 4564 62270 4616
rect 65058 4604 65064 4616
rect 65019 4576 65064 4604
rect 65058 4564 65064 4576
rect 65116 4564 65122 4616
rect 69842 4604 69848 4616
rect 69803 4576 69848 4604
rect 69842 4564 69848 4576
rect 69900 4564 69906 4616
rect 70949 4607 71007 4613
rect 70949 4604 70961 4607
rect 70228 4576 70961 4604
rect 33744 4508 35388 4536
rect 36817 4539 36875 4545
rect 33744 4496 33750 4508
rect 36817 4505 36829 4539
rect 36863 4536 36875 4539
rect 36906 4536 36912 4548
rect 36863 4508 36912 4536
rect 36863 4505 36875 4508
rect 36817 4499 36875 4505
rect 36906 4496 36912 4508
rect 36964 4536 36970 4548
rect 47118 4536 47124 4548
rect 36964 4508 39528 4536
rect 36964 4496 36970 4508
rect 6362 4468 6368 4480
rect 6323 4440 6368 4468
rect 6362 4428 6368 4440
rect 6420 4428 6426 4480
rect 22649 4471 22707 4477
rect 22649 4437 22661 4471
rect 22695 4468 22707 4471
rect 23290 4468 23296 4480
rect 22695 4440 23296 4468
rect 22695 4437 22707 4440
rect 22649 4431 22707 4437
rect 23290 4428 23296 4440
rect 23348 4428 23354 4480
rect 23842 4468 23848 4480
rect 23803 4440 23848 4468
rect 23842 4428 23848 4440
rect 23900 4428 23906 4480
rect 27614 4468 27620 4480
rect 27575 4440 27620 4468
rect 27614 4428 27620 4440
rect 27672 4428 27678 4480
rect 30190 4428 30196 4480
rect 30248 4468 30254 4480
rect 30377 4471 30435 4477
rect 30377 4468 30389 4471
rect 30248 4440 30389 4468
rect 30248 4428 30254 4440
rect 30377 4437 30389 4440
rect 30423 4437 30435 4471
rect 30377 4431 30435 4437
rect 31941 4471 31999 4477
rect 31941 4437 31953 4471
rect 31987 4468 31999 4471
rect 32306 4468 32312 4480
rect 31987 4440 32312 4468
rect 31987 4437 31999 4440
rect 31941 4431 31999 4437
rect 32306 4428 32312 4440
rect 32364 4428 32370 4480
rect 32766 4468 32772 4480
rect 32727 4440 32772 4468
rect 32766 4428 32772 4440
rect 32824 4428 32830 4480
rect 35894 4428 35900 4480
rect 35952 4468 35958 4480
rect 37274 4468 37280 4480
rect 35952 4440 35997 4468
rect 37235 4440 37280 4468
rect 35952 4428 35958 4440
rect 37274 4428 37280 4440
rect 37332 4428 37338 4480
rect 38562 4428 38568 4480
rect 38620 4468 38626 4480
rect 39500 4477 39528 4508
rect 46492 4508 47124 4536
rect 38749 4471 38807 4477
rect 38749 4468 38761 4471
rect 38620 4440 38761 4468
rect 38620 4428 38626 4440
rect 38749 4437 38761 4440
rect 38795 4437 38807 4471
rect 38749 4431 38807 4437
rect 39485 4471 39543 4477
rect 39485 4437 39497 4471
rect 39531 4468 39543 4471
rect 41233 4471 41291 4477
rect 41233 4468 41245 4471
rect 39531 4440 41245 4468
rect 39531 4437 39543 4440
rect 39485 4431 39543 4437
rect 41233 4437 41245 4440
rect 41279 4468 41291 4471
rect 41322 4468 41328 4480
rect 41279 4440 41328 4468
rect 41279 4437 41291 4440
rect 41233 4431 41291 4437
rect 41322 4428 41328 4440
rect 41380 4428 41386 4480
rect 42521 4471 42579 4477
rect 42521 4437 42533 4471
rect 42567 4468 42579 4471
rect 42978 4468 42984 4480
rect 42567 4440 42984 4468
rect 42567 4437 42579 4440
rect 42521 4431 42579 4437
rect 42978 4428 42984 4440
rect 43036 4428 43042 4480
rect 45922 4428 45928 4480
rect 45980 4468 45986 4480
rect 46492 4477 46520 4508
rect 47118 4496 47124 4508
rect 47176 4536 47182 4548
rect 47578 4536 47584 4548
rect 47176 4508 47584 4536
rect 47176 4496 47182 4508
rect 47578 4496 47584 4508
rect 47636 4496 47642 4548
rect 48314 4496 48320 4548
rect 48372 4536 48378 4548
rect 48409 4539 48467 4545
rect 48409 4536 48421 4539
rect 48372 4508 48421 4536
rect 48372 4496 48378 4508
rect 48409 4505 48421 4508
rect 48455 4505 48467 4539
rect 48409 4499 48467 4505
rect 57790 4496 57796 4548
rect 57848 4536 57854 4548
rect 58437 4539 58495 4545
rect 58437 4536 58449 4539
rect 57848 4508 58449 4536
rect 57848 4496 57854 4508
rect 58437 4505 58449 4508
rect 58483 4505 58495 4539
rect 58437 4499 58495 4505
rect 64141 4539 64199 4545
rect 64141 4505 64153 4539
rect 64187 4505 64199 4539
rect 70228 4536 70256 4576
rect 70949 4573 70961 4576
rect 70995 4604 71007 4607
rect 71590 4604 71596 4616
rect 70995 4576 71596 4604
rect 70995 4573 71007 4576
rect 70949 4567 71007 4573
rect 71590 4564 71596 4576
rect 71648 4564 71654 4616
rect 79689 4607 79747 4613
rect 79689 4573 79701 4607
rect 79735 4604 79747 4607
rect 80054 4604 80060 4616
rect 79735 4576 80060 4604
rect 79735 4573 79747 4576
rect 79689 4567 79747 4573
rect 80054 4564 80060 4576
rect 80112 4564 80118 4616
rect 80422 4604 80428 4616
rect 80383 4576 80428 4604
rect 80422 4564 80428 4576
rect 80480 4564 80486 4616
rect 81452 4613 81480 4644
rect 81986 4632 81992 4644
rect 82044 4672 82050 4684
rect 82044 4644 82676 4672
rect 82044 4632 82050 4644
rect 81437 4607 81495 4613
rect 81437 4573 81449 4607
rect 81483 4573 81495 4607
rect 82078 4604 82084 4616
rect 82039 4576 82084 4604
rect 81437 4567 81495 4573
rect 82078 4564 82084 4576
rect 82136 4564 82142 4616
rect 64141 4499 64199 4505
rect 68664 4508 70256 4536
rect 46477 4471 46535 4477
rect 46477 4468 46489 4471
rect 45980 4440 46489 4468
rect 45980 4428 45986 4440
rect 46477 4437 46489 4440
rect 46523 4437 46535 4471
rect 47026 4468 47032 4480
rect 46987 4440 47032 4468
rect 46477 4431 46535 4437
rect 47026 4428 47032 4440
rect 47084 4428 47090 4480
rect 50433 4471 50491 4477
rect 50433 4437 50445 4471
rect 50479 4468 50491 4471
rect 50614 4468 50620 4480
rect 50479 4440 50620 4468
rect 50479 4437 50491 4440
rect 50433 4431 50491 4437
rect 50614 4428 50620 4440
rect 50672 4428 50678 4480
rect 51626 4428 51632 4480
rect 51684 4468 51690 4480
rect 51721 4471 51779 4477
rect 51721 4468 51733 4471
rect 51684 4440 51733 4468
rect 51684 4428 51690 4440
rect 51721 4437 51733 4440
rect 51767 4437 51779 4471
rect 51721 4431 51779 4437
rect 52454 4428 52460 4480
rect 52512 4468 52518 4480
rect 52733 4471 52791 4477
rect 52733 4468 52745 4471
rect 52512 4440 52745 4468
rect 52512 4428 52518 4440
rect 52733 4437 52745 4440
rect 52779 4437 52791 4471
rect 54294 4468 54300 4480
rect 54255 4440 54300 4468
rect 52733 4431 52791 4437
rect 54294 4428 54300 4440
rect 54352 4428 54358 4480
rect 56045 4471 56103 4477
rect 56045 4437 56057 4471
rect 56091 4468 56103 4471
rect 56318 4468 56324 4480
rect 56091 4440 56324 4468
rect 56091 4437 56103 4440
rect 56045 4431 56103 4437
rect 56318 4428 56324 4440
rect 56376 4428 56382 4480
rect 56410 4428 56416 4480
rect 56468 4468 56474 4480
rect 56597 4471 56655 4477
rect 56597 4468 56609 4471
rect 56468 4440 56609 4468
rect 56468 4428 56474 4440
rect 56597 4437 56609 4440
rect 56643 4437 56655 4471
rect 56597 4431 56655 4437
rect 57241 4471 57299 4477
rect 57241 4437 57253 4471
rect 57287 4468 57299 4471
rect 58342 4468 58348 4480
rect 57287 4440 58348 4468
rect 57287 4437 57299 4440
rect 57241 4431 57299 4437
rect 58342 4428 58348 4440
rect 58400 4428 58406 4480
rect 61470 4428 61476 4480
rect 61528 4468 61534 4480
rect 61657 4471 61715 4477
rect 61657 4468 61669 4471
rect 61528 4440 61669 4468
rect 61528 4428 61534 4440
rect 61657 4437 61669 4440
rect 61703 4437 61715 4471
rect 62298 4468 62304 4480
rect 62259 4440 62304 4468
rect 61657 4431 61715 4437
rect 62298 4428 62304 4440
rect 62356 4428 62362 4480
rect 63402 4428 63408 4480
rect 63460 4468 63466 4480
rect 63497 4471 63555 4477
rect 63497 4468 63509 4471
rect 63460 4440 63509 4468
rect 63460 4428 63466 4440
rect 63497 4437 63509 4440
rect 63543 4468 63555 4471
rect 64156 4468 64184 4499
rect 68664 4480 68692 4508
rect 70302 4496 70308 4548
rect 70360 4536 70366 4548
rect 71501 4539 71559 4545
rect 71501 4536 71513 4539
rect 70360 4508 71513 4536
rect 70360 4496 70366 4508
rect 71501 4505 71513 4508
rect 71547 4505 71559 4539
rect 71501 4499 71559 4505
rect 80330 4496 80336 4548
rect 80388 4536 80394 4548
rect 82648 4545 82676 4644
rect 82633 4539 82691 4545
rect 80388 4508 81940 4536
rect 80388 4496 80394 4508
rect 64414 4468 64420 4480
rect 63543 4440 64184 4468
rect 64375 4440 64420 4468
rect 63543 4437 63555 4440
rect 63497 4431 63555 4437
rect 64414 4428 64420 4440
rect 64472 4428 64478 4480
rect 65242 4468 65248 4480
rect 65203 4440 65248 4468
rect 65242 4428 65248 4440
rect 65300 4428 65306 4480
rect 68646 4468 68652 4480
rect 68607 4440 68652 4468
rect 68646 4428 68652 4440
rect 68704 4428 68710 4480
rect 69198 4468 69204 4480
rect 69159 4440 69204 4468
rect 69198 4428 69204 4440
rect 69256 4428 69262 4480
rect 70029 4471 70087 4477
rect 70029 4437 70041 4471
rect 70075 4468 70087 4471
rect 70394 4468 70400 4480
rect 70075 4440 70400 4468
rect 70075 4437 70087 4440
rect 70029 4431 70087 4437
rect 70394 4428 70400 4440
rect 70452 4428 70458 4480
rect 74997 4471 75055 4477
rect 74997 4437 75009 4471
rect 75043 4468 75055 4471
rect 75086 4468 75092 4480
rect 75043 4440 75092 4468
rect 75043 4437 75055 4440
rect 74997 4431 75055 4437
rect 75086 4428 75092 4440
rect 75144 4428 75150 4480
rect 77662 4468 77668 4480
rect 77623 4440 77668 4468
rect 77662 4428 77668 4440
rect 77720 4428 77726 4480
rect 78674 4468 78680 4480
rect 78635 4440 78680 4468
rect 78674 4428 78680 4440
rect 78732 4428 78738 4480
rect 78766 4428 78772 4480
rect 78824 4468 78830 4480
rect 79229 4471 79287 4477
rect 79229 4468 79241 4471
rect 78824 4440 79241 4468
rect 78824 4428 78830 4440
rect 79229 4437 79241 4440
rect 79275 4437 79287 4471
rect 79229 4431 79287 4437
rect 79597 4471 79655 4477
rect 79597 4437 79609 4471
rect 79643 4468 79655 4471
rect 80146 4468 80152 4480
rect 79643 4440 80152 4468
rect 79643 4437 79655 4440
rect 79597 4431 79655 4437
rect 80146 4428 80152 4440
rect 80204 4428 80210 4480
rect 81342 4468 81348 4480
rect 81303 4440 81348 4468
rect 81342 4428 81348 4440
rect 81400 4428 81406 4480
rect 81912 4477 81940 4508
rect 82633 4505 82645 4539
rect 82679 4536 82691 4539
rect 84194 4536 84200 4548
rect 82679 4508 84200 4536
rect 82679 4505 82691 4508
rect 82633 4499 82691 4505
rect 84194 4496 84200 4508
rect 84252 4496 84258 4548
rect 81897 4471 81955 4477
rect 81897 4437 81909 4471
rect 81943 4437 81955 4471
rect 81897 4431 81955 4437
rect 82814 4428 82820 4480
rect 82872 4468 82878 4480
rect 83645 4471 83703 4477
rect 83645 4468 83657 4471
rect 82872 4440 83657 4468
rect 82872 4428 82878 4440
rect 83645 4437 83657 4440
rect 83691 4437 83703 4471
rect 83645 4431 83703 4437
rect 1104 4378 148856 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 81014 4378
rect 81066 4326 81078 4378
rect 81130 4326 81142 4378
rect 81194 4326 81206 4378
rect 81258 4326 81270 4378
rect 81322 4326 111734 4378
rect 111786 4326 111798 4378
rect 111850 4326 111862 4378
rect 111914 4326 111926 4378
rect 111978 4326 111990 4378
rect 112042 4326 142454 4378
rect 142506 4326 142518 4378
rect 142570 4326 142582 4378
rect 142634 4326 142646 4378
rect 142698 4326 142710 4378
rect 142762 4326 148856 4378
rect 1104 4304 148856 4326
rect 32766 4224 32772 4276
rect 32824 4264 32830 4276
rect 49050 4264 49056 4276
rect 32824 4236 49056 4264
rect 32824 4224 32830 4236
rect 49050 4224 49056 4236
rect 49108 4224 49114 4276
rect 54294 4224 54300 4276
rect 54352 4264 54358 4276
rect 63402 4264 63408 4276
rect 54352 4236 63408 4264
rect 54352 4224 54358 4236
rect 63402 4224 63408 4236
rect 63460 4224 63466 4276
rect 64414 4224 64420 4276
rect 64472 4264 64478 4276
rect 67177 4267 67235 4273
rect 67177 4264 67189 4267
rect 64472 4236 67189 4264
rect 64472 4224 64478 4236
rect 67177 4233 67189 4236
rect 67223 4264 67235 4267
rect 68278 4264 68284 4276
rect 67223 4236 68284 4264
rect 67223 4233 67235 4236
rect 67177 4227 67235 4233
rect 68278 4224 68284 4236
rect 68336 4264 68342 4276
rect 68646 4264 68652 4276
rect 68336 4236 68652 4264
rect 68336 4224 68342 4236
rect 68646 4224 68652 4236
rect 68704 4224 68710 4276
rect 81434 4264 81440 4276
rect 81395 4236 81440 4264
rect 81434 4224 81440 4236
rect 81492 4224 81498 4276
rect 81805 4267 81863 4273
rect 81805 4233 81817 4267
rect 81851 4264 81863 4267
rect 82722 4264 82728 4276
rect 81851 4236 82728 4264
rect 81851 4233 81863 4236
rect 81805 4227 81863 4233
rect 82722 4224 82728 4236
rect 82780 4224 82786 4276
rect 26326 4156 26332 4208
rect 26384 4196 26390 4208
rect 26605 4199 26663 4205
rect 26605 4196 26617 4199
rect 26384 4168 26617 4196
rect 26384 4156 26390 4168
rect 26605 4165 26617 4168
rect 26651 4196 26663 4199
rect 26651 4168 28028 4196
rect 26651 4165 26663 4168
rect 26605 4159 26663 4165
rect 5994 4088 6000 4140
rect 6052 4128 6058 4140
rect 6549 4131 6607 4137
rect 6549 4128 6561 4131
rect 6052 4100 6561 4128
rect 6052 4088 6058 4100
rect 6549 4097 6561 4100
rect 6595 4097 6607 4131
rect 6549 4091 6607 4097
rect 22465 4131 22523 4137
rect 22465 4097 22477 4131
rect 22511 4128 22523 4131
rect 22738 4128 22744 4140
rect 22511 4100 22744 4128
rect 22511 4097 22523 4100
rect 22465 4091 22523 4097
rect 22738 4088 22744 4100
rect 22796 4088 22802 4140
rect 23569 4131 23627 4137
rect 23569 4097 23581 4131
rect 23615 4097 23627 4131
rect 27338 4128 27344 4140
rect 27299 4100 27344 4128
rect 23569 4091 23627 4097
rect 23584 4060 23612 4091
rect 27338 4088 27344 4100
rect 27396 4088 27402 4140
rect 28000 4137 28028 4168
rect 35618 4156 35624 4208
rect 35676 4196 35682 4208
rect 35805 4199 35863 4205
rect 35805 4196 35817 4199
rect 35676 4168 35817 4196
rect 35676 4156 35682 4168
rect 35805 4165 35817 4168
rect 35851 4165 35863 4199
rect 35805 4159 35863 4165
rect 37274 4156 37280 4208
rect 37332 4196 37338 4208
rect 37553 4199 37611 4205
rect 37553 4196 37565 4199
rect 37332 4168 37565 4196
rect 37332 4156 37338 4168
rect 37553 4165 37565 4168
rect 37599 4165 37611 4199
rect 44269 4199 44327 4205
rect 37553 4159 37611 4165
rect 39776 4168 40080 4196
rect 27985 4131 28043 4137
rect 27985 4097 27997 4131
rect 28031 4128 28043 4131
rect 28031 4100 28580 4128
rect 28031 4097 28043 4100
rect 27985 4091 28043 4097
rect 28442 4060 28448 4072
rect 23584 4032 28448 4060
rect 28442 4020 28448 4032
rect 28500 4020 28506 4072
rect 6638 3952 6644 4004
rect 6696 3992 6702 4004
rect 7193 3995 7251 4001
rect 7193 3992 7205 3995
rect 6696 3964 7205 3992
rect 6696 3952 6702 3964
rect 7193 3961 7205 3964
rect 7239 3961 7251 3995
rect 7193 3955 7251 3961
rect 23750 3952 23756 4004
rect 23808 3992 23814 4004
rect 24673 3995 24731 4001
rect 24673 3992 24685 3995
rect 23808 3964 24685 3992
rect 23808 3952 23814 3964
rect 24673 3961 24685 3964
rect 24719 3992 24731 3995
rect 26234 3992 26240 4004
rect 24719 3964 26240 3992
rect 24719 3961 24731 3964
rect 24673 3955 24731 3961
rect 26234 3952 26240 3964
rect 26292 3952 26298 4004
rect 28552 4001 28580 4100
rect 28810 4088 28816 4140
rect 28868 4128 28874 4140
rect 28997 4131 29055 4137
rect 28997 4128 29009 4131
rect 28868 4100 29009 4128
rect 28868 4088 28874 4100
rect 28997 4097 29009 4100
rect 29043 4097 29055 4131
rect 32769 4131 32827 4137
rect 32769 4128 32781 4131
rect 28997 4091 29055 4097
rect 29104 4100 32781 4128
rect 28537 3995 28595 4001
rect 28537 3961 28549 3995
rect 28583 3992 28595 3995
rect 29104 3992 29132 4100
rect 32769 4097 32781 4100
rect 32815 4128 32827 4131
rect 33229 4131 33287 4137
rect 33229 4128 33241 4131
rect 32815 4100 33241 4128
rect 32815 4097 32827 4100
rect 32769 4091 32827 4097
rect 33229 4097 33241 4100
rect 33275 4128 33287 4131
rect 33686 4128 33692 4140
rect 33275 4100 33692 4128
rect 33275 4097 33287 4100
rect 33229 4091 33287 4097
rect 33686 4088 33692 4100
rect 33744 4088 33750 4140
rect 33778 4088 33784 4140
rect 33836 4128 33842 4140
rect 34057 4131 34115 4137
rect 34057 4128 34069 4131
rect 33836 4100 34069 4128
rect 33836 4088 33842 4100
rect 34057 4097 34069 4100
rect 34103 4097 34115 4131
rect 34057 4091 34115 4097
rect 34146 4088 34152 4140
rect 34204 4128 34210 4140
rect 34977 4131 35035 4137
rect 34977 4128 34989 4131
rect 34204 4100 34989 4128
rect 34204 4088 34210 4100
rect 34977 4097 34989 4100
rect 35023 4097 35035 4131
rect 35986 4128 35992 4140
rect 35947 4100 35992 4128
rect 34977 4091 35035 4097
rect 35986 4088 35992 4100
rect 36044 4088 36050 4140
rect 36449 4131 36507 4137
rect 36449 4097 36461 4131
rect 36495 4128 36507 4131
rect 37458 4128 37464 4140
rect 36495 4100 37464 4128
rect 36495 4097 36507 4100
rect 36449 4091 36507 4097
rect 37458 4088 37464 4100
rect 37516 4088 37522 4140
rect 37642 4088 37648 4140
rect 37700 4128 37706 4140
rect 37737 4131 37795 4137
rect 37737 4128 37749 4131
rect 37700 4100 37749 4128
rect 37700 4088 37706 4100
rect 37737 4097 37749 4100
rect 37783 4097 37795 4131
rect 37737 4091 37795 4097
rect 38010 4088 38016 4140
rect 38068 4128 38074 4140
rect 38197 4131 38255 4137
rect 38197 4128 38209 4131
rect 38068 4100 38209 4128
rect 38068 4088 38074 4100
rect 38197 4097 38209 4100
rect 38243 4097 38255 4131
rect 38197 4091 38255 4097
rect 39393 4131 39451 4137
rect 39393 4097 39405 4131
rect 39439 4128 39451 4131
rect 39776 4128 39804 4168
rect 40052 4140 40080 4168
rect 44269 4165 44281 4199
rect 44315 4165 44327 4199
rect 44269 4159 44327 4165
rect 48133 4199 48191 4205
rect 48133 4165 48145 4199
rect 48179 4196 48191 4199
rect 49510 4196 49516 4208
rect 48179 4168 49516 4196
rect 48179 4165 48191 4168
rect 48133 4159 48191 4165
rect 39439 4100 39804 4128
rect 39439 4097 39451 4100
rect 39393 4091 39451 4097
rect 39850 4088 39856 4140
rect 39908 4128 39914 4140
rect 39908 4100 39953 4128
rect 39908 4088 39914 4100
rect 40034 4088 40040 4140
rect 40092 4088 40098 4140
rect 42061 4131 42119 4137
rect 42061 4097 42073 4131
rect 42107 4128 42119 4131
rect 42150 4128 42156 4140
rect 42107 4100 42156 4128
rect 42107 4097 42119 4100
rect 42061 4091 42119 4097
rect 42150 4088 42156 4100
rect 42208 4088 42214 4140
rect 42981 4131 43039 4137
rect 42981 4097 42993 4131
rect 43027 4128 43039 4131
rect 43806 4128 43812 4140
rect 43027 4100 43812 4128
rect 43027 4097 43039 4100
rect 42981 4091 43039 4097
rect 43806 4088 43812 4100
rect 43864 4088 43870 4140
rect 43898 4088 43904 4140
rect 43956 4128 43962 4140
rect 44284 4128 44312 4159
rect 49510 4156 49516 4168
rect 49568 4196 49574 4208
rect 49568 4168 49924 4196
rect 49568 4156 49574 4168
rect 43956 4100 44312 4128
rect 43956 4088 43962 4100
rect 44358 4088 44364 4140
rect 44416 4128 44422 4140
rect 44453 4131 44511 4137
rect 44453 4128 44465 4131
rect 44416 4100 44465 4128
rect 44416 4088 44422 4100
rect 44453 4097 44465 4100
rect 44499 4097 44511 4131
rect 44453 4091 44511 4097
rect 46293 4131 46351 4137
rect 46293 4097 46305 4131
rect 46339 4097 46351 4131
rect 47026 4128 47032 4140
rect 46987 4100 47032 4128
rect 46293 4091 46351 4097
rect 29641 4063 29699 4069
rect 29641 4029 29653 4063
rect 29687 4060 29699 4063
rect 29822 4060 29828 4072
rect 29687 4032 29828 4060
rect 29687 4029 29699 4032
rect 29641 4023 29699 4029
rect 28583 3964 29132 3992
rect 28583 3961 28595 3964
rect 28537 3955 28595 3961
rect 5997 3927 6055 3933
rect 5997 3893 6009 3927
rect 6043 3924 6055 3927
rect 6270 3924 6276 3936
rect 6043 3896 6276 3924
rect 6043 3893 6055 3896
rect 5997 3887 6055 3893
rect 6270 3884 6276 3896
rect 6328 3884 6334 3936
rect 6733 3927 6791 3933
rect 6733 3893 6745 3927
rect 6779 3924 6791 3927
rect 6822 3924 6828 3936
rect 6779 3896 6828 3924
rect 6779 3893 6791 3896
rect 6733 3887 6791 3893
rect 6822 3884 6828 3896
rect 6880 3884 6886 3936
rect 8018 3924 8024 3936
rect 7979 3896 8024 3924
rect 8018 3884 8024 3896
rect 8076 3884 8082 3936
rect 22278 3924 22284 3936
rect 22239 3896 22284 3924
rect 22278 3884 22284 3896
rect 22336 3884 22342 3936
rect 23198 3884 23204 3936
rect 23256 3924 23262 3936
rect 23385 3927 23443 3933
rect 23385 3924 23397 3927
rect 23256 3896 23397 3924
rect 23256 3884 23262 3896
rect 23385 3893 23397 3896
rect 23431 3893 23443 3927
rect 23385 3887 23443 3893
rect 24121 3927 24179 3933
rect 24121 3893 24133 3927
rect 24167 3924 24179 3927
rect 24946 3924 24952 3936
rect 24167 3896 24952 3924
rect 24167 3893 24179 3896
rect 24121 3887 24179 3893
rect 24946 3884 24952 3896
rect 25004 3884 25010 3936
rect 25958 3924 25964 3936
rect 25919 3896 25964 3924
rect 25958 3884 25964 3896
rect 26016 3884 26022 3936
rect 27154 3924 27160 3936
rect 27115 3896 27160 3924
rect 27154 3884 27160 3896
rect 27212 3884 27218 3936
rect 27890 3924 27896 3936
rect 27851 3896 27896 3924
rect 27890 3884 27896 3896
rect 27948 3884 27954 3936
rect 27982 3884 27988 3936
rect 28040 3924 28046 3936
rect 29656 3924 29684 4023
rect 29822 4020 29828 4032
rect 29880 4060 29886 4072
rect 46106 4060 46112 4072
rect 29880 4032 46112 4060
rect 29880 4020 29886 4032
rect 46106 4020 46112 4032
rect 46164 4020 46170 4072
rect 38562 3952 38568 4004
rect 38620 3992 38626 4004
rect 41417 3995 41475 4001
rect 41417 3992 41429 3995
rect 38620 3964 41429 3992
rect 38620 3952 38626 3964
rect 41417 3961 41429 3964
rect 41463 3992 41475 3995
rect 41598 3992 41604 4004
rect 41463 3964 41604 3992
rect 41463 3961 41475 3964
rect 41417 3955 41475 3961
rect 41598 3952 41604 3964
rect 41656 3952 41662 4004
rect 42426 3952 42432 4004
rect 42484 3992 42490 4004
rect 46308 3992 46336 4091
rect 47026 4088 47032 4100
rect 47084 4088 47090 4140
rect 48225 4131 48283 4137
rect 48225 4097 48237 4131
rect 48271 4128 48283 4131
rect 48958 4128 48964 4140
rect 48271 4100 48964 4128
rect 48271 4097 48283 4100
rect 48225 4091 48283 4097
rect 48958 4088 48964 4100
rect 49016 4088 49022 4140
rect 49053 4131 49111 4137
rect 49053 4097 49065 4131
rect 49099 4128 49111 4131
rect 49418 4128 49424 4140
rect 49099 4100 49424 4128
rect 49099 4097 49111 4100
rect 49053 4091 49111 4097
rect 49418 4088 49424 4100
rect 49476 4128 49482 4140
rect 49605 4131 49663 4137
rect 49605 4128 49617 4131
rect 49476 4100 49617 4128
rect 49476 4088 49482 4100
rect 49605 4097 49617 4100
rect 49651 4097 49663 4131
rect 49605 4091 49663 4097
rect 49694 4088 49700 4140
rect 49752 4128 49758 4140
rect 49789 4131 49847 4137
rect 49789 4128 49801 4131
rect 49752 4100 49801 4128
rect 49752 4088 49758 4100
rect 49789 4097 49801 4100
rect 49835 4097 49847 4131
rect 49789 4091 49847 4097
rect 47578 4020 47584 4072
rect 47636 4060 47642 4072
rect 48317 4063 48375 4069
rect 48317 4060 48329 4063
rect 47636 4032 48329 4060
rect 47636 4020 47642 4032
rect 48317 4029 48329 4032
rect 48363 4029 48375 4063
rect 49896 4060 49924 4168
rect 51442 4156 51448 4208
rect 51500 4196 51506 4208
rect 51500 4168 52408 4196
rect 51500 4156 51506 4168
rect 51077 4131 51135 4137
rect 51077 4097 51089 4131
rect 51123 4128 51135 4131
rect 51350 4128 51356 4140
rect 51123 4100 51356 4128
rect 51123 4097 51135 4100
rect 51077 4091 51135 4097
rect 51350 4088 51356 4100
rect 51408 4088 51414 4140
rect 51721 4131 51779 4137
rect 51721 4097 51733 4131
rect 51767 4128 51779 4131
rect 52178 4128 52184 4140
rect 51767 4100 52184 4128
rect 51767 4097 51779 4100
rect 51721 4091 51779 4097
rect 52178 4088 52184 4100
rect 52236 4088 52242 4140
rect 52380 4137 52408 4168
rect 52454 4156 52460 4208
rect 52512 4196 52518 4208
rect 53009 4199 53067 4205
rect 53009 4196 53021 4199
rect 52512 4168 53021 4196
rect 52512 4156 52518 4168
rect 53009 4165 53021 4168
rect 53055 4165 53067 4199
rect 53009 4159 53067 4165
rect 55048 4168 55352 4196
rect 52365 4131 52423 4137
rect 52365 4097 52377 4131
rect 52411 4097 52423 4131
rect 52365 4091 52423 4097
rect 53098 4088 53104 4140
rect 53156 4128 53162 4140
rect 53193 4131 53251 4137
rect 53193 4128 53205 4131
rect 53156 4100 53205 4128
rect 53156 4088 53162 4100
rect 53193 4097 53205 4100
rect 53239 4097 53251 4131
rect 53193 4091 53251 4097
rect 55048 4060 55076 4168
rect 55125 4131 55183 4137
rect 55125 4097 55137 4131
rect 55171 4128 55183 4131
rect 55171 4100 55260 4128
rect 55171 4097 55183 4100
rect 55125 4091 55183 4097
rect 49896 4032 55076 4060
rect 48317 4023 48375 4029
rect 49326 3992 49332 4004
rect 42484 3964 45140 3992
rect 46308 3964 49332 3992
rect 42484 3952 42490 3964
rect 45112 3936 45140 3964
rect 49326 3952 49332 3964
rect 49384 3992 49390 4004
rect 51442 3992 51448 4004
rect 49384 3964 51448 3992
rect 49384 3952 49390 3964
rect 51442 3952 51448 3964
rect 51500 3992 51506 4004
rect 55140 3992 55168 4091
rect 51500 3964 55168 3992
rect 55232 3992 55260 4100
rect 55324 4060 55352 4168
rect 56318 4156 56324 4208
rect 56376 4196 56382 4208
rect 56505 4199 56563 4205
rect 56505 4196 56517 4199
rect 56376 4168 56517 4196
rect 56376 4156 56382 4168
rect 56505 4165 56517 4168
rect 56551 4165 56563 4199
rect 64693 4199 64751 4205
rect 64693 4196 64705 4199
rect 56505 4159 56563 4165
rect 64524 4168 64705 4196
rect 55858 4128 55864 4140
rect 55819 4100 55864 4128
rect 55858 4088 55864 4100
rect 55916 4088 55922 4140
rect 56594 4088 56600 4140
rect 56652 4128 56658 4140
rect 56689 4131 56747 4137
rect 56689 4128 56701 4131
rect 56652 4100 56701 4128
rect 56652 4088 56658 4100
rect 56689 4097 56701 4100
rect 56735 4097 56747 4131
rect 56689 4091 56747 4097
rect 57333 4131 57391 4137
rect 57333 4097 57345 4131
rect 57379 4128 57391 4131
rect 57422 4128 57428 4140
rect 57379 4100 57428 4128
rect 57379 4097 57391 4100
rect 57333 4091 57391 4097
rect 57422 4088 57428 4100
rect 57480 4088 57486 4140
rect 58069 4131 58127 4137
rect 58069 4128 58081 4131
rect 57992 4100 58081 4128
rect 57146 4060 57152 4072
rect 55324 4032 57152 4060
rect 57146 4020 57152 4032
rect 57204 4020 57210 4072
rect 56502 3992 56508 4004
rect 55232 3964 56508 3992
rect 51500 3952 51506 3964
rect 56502 3952 56508 3964
rect 56560 3992 56566 4004
rect 57992 3992 58020 4100
rect 58069 4097 58081 4100
rect 58115 4128 58127 4131
rect 60093 4131 60151 4137
rect 58115 4100 60044 4128
rect 58115 4097 58127 4100
rect 58069 4091 58127 4097
rect 60016 4060 60044 4100
rect 60093 4097 60105 4131
rect 60139 4128 60151 4131
rect 60458 4128 60464 4140
rect 60139 4100 60464 4128
rect 60139 4097 60151 4100
rect 60093 4091 60151 4097
rect 60458 4088 60464 4100
rect 60516 4128 60522 4140
rect 60645 4131 60703 4137
rect 60645 4128 60657 4131
rect 60516 4100 60657 4128
rect 60516 4088 60522 4100
rect 60645 4097 60657 4100
rect 60691 4097 60703 4131
rect 60645 4091 60703 4097
rect 60734 4088 60740 4140
rect 60792 4128 60798 4140
rect 60829 4131 60887 4137
rect 60829 4128 60841 4131
rect 60792 4100 60841 4128
rect 60792 4088 60798 4100
rect 60829 4097 60841 4100
rect 60875 4097 60887 4131
rect 60829 4091 60887 4097
rect 61473 4131 61531 4137
rect 61473 4097 61485 4131
rect 61519 4128 61531 4131
rect 62206 4128 62212 4140
rect 61519 4100 62212 4128
rect 61519 4097 61531 4100
rect 61473 4091 61531 4097
rect 61488 4060 61516 4091
rect 62206 4088 62212 4100
rect 62264 4128 62270 4140
rect 62301 4131 62359 4137
rect 62301 4128 62313 4131
rect 62264 4100 62313 4128
rect 62264 4088 62270 4100
rect 62301 4097 62313 4100
rect 62347 4097 62359 4131
rect 63310 4128 63316 4140
rect 63271 4100 63316 4128
rect 62301 4091 62359 4097
rect 63310 4088 63316 4100
rect 63368 4088 63374 4140
rect 60016 4032 61516 4060
rect 63862 4020 63868 4072
rect 63920 4060 63926 4072
rect 64417 4063 64475 4069
rect 64417 4060 64429 4063
rect 63920 4032 64429 4060
rect 63920 4020 63926 4032
rect 64417 4029 64429 4032
rect 64463 4029 64475 4063
rect 64417 4023 64475 4029
rect 56560 3964 58020 3992
rect 58161 3995 58219 4001
rect 56560 3952 56566 3964
rect 58161 3961 58173 3995
rect 58207 3992 58219 3995
rect 59354 3992 59360 4004
rect 58207 3964 59360 3992
rect 58207 3961 58219 3964
rect 58161 3955 58219 3961
rect 59354 3952 59360 3964
rect 59412 3952 59418 4004
rect 62393 3995 62451 4001
rect 62393 3961 62405 3995
rect 62439 3992 62451 3995
rect 63954 3992 63960 4004
rect 62439 3964 63960 3992
rect 62439 3961 62451 3964
rect 62393 3955 62451 3961
rect 63954 3952 63960 3964
rect 64012 3952 64018 4004
rect 64524 3992 64552 4168
rect 64693 4165 64705 4168
rect 64739 4165 64751 4199
rect 66070 4196 66076 4208
rect 64693 4159 64751 4165
rect 64984 4168 66076 4196
rect 64601 4063 64659 4069
rect 64601 4029 64613 4063
rect 64647 4060 64659 4063
rect 64984 4060 65012 4168
rect 66070 4156 66076 4168
rect 66128 4156 66134 4208
rect 69290 4156 69296 4208
rect 69348 4196 69354 4208
rect 79413 4199 79471 4205
rect 69348 4168 70150 4196
rect 69348 4156 69354 4168
rect 79413 4165 79425 4199
rect 79459 4196 79471 4199
rect 79502 4196 79508 4208
rect 79459 4168 79508 4196
rect 79459 4165 79471 4168
rect 79413 4159 79471 4165
rect 79502 4156 79508 4168
rect 79560 4156 79566 4208
rect 81342 4196 81348 4208
rect 80638 4168 81348 4196
rect 81342 4156 81348 4168
rect 81400 4156 81406 4208
rect 65705 4131 65763 4137
rect 65705 4128 65717 4131
rect 64647 4032 65012 4060
rect 65076 4100 65717 4128
rect 64647 4029 64659 4032
rect 64601 4023 64659 4029
rect 65076 4001 65104 4100
rect 65705 4097 65717 4100
rect 65751 4097 65763 4131
rect 66530 4128 66536 4140
rect 66491 4100 66536 4128
rect 65705 4091 65763 4097
rect 66530 4088 66536 4100
rect 66588 4088 66594 4140
rect 68741 4131 68799 4137
rect 68741 4097 68753 4131
rect 68787 4128 68799 4131
rect 68830 4128 68836 4140
rect 68787 4100 68836 4128
rect 68787 4097 68799 4100
rect 68741 4091 68799 4097
rect 68830 4088 68836 4100
rect 68888 4088 68894 4140
rect 71406 4088 71412 4140
rect 71464 4128 71470 4140
rect 71777 4131 71835 4137
rect 71777 4128 71789 4131
rect 71464 4100 71789 4128
rect 71464 4088 71470 4100
rect 71777 4097 71789 4100
rect 71823 4097 71835 4131
rect 75730 4128 75736 4140
rect 75691 4100 75736 4128
rect 71777 4091 71835 4097
rect 75730 4088 75736 4100
rect 75788 4088 75794 4140
rect 77941 4131 77999 4137
rect 77941 4097 77953 4131
rect 77987 4128 77999 4131
rect 78766 4128 78772 4140
rect 77987 4100 78772 4128
rect 77987 4097 77999 4100
rect 77941 4091 77999 4097
rect 78766 4088 78772 4100
rect 78824 4088 78830 4140
rect 81897 4131 81955 4137
rect 81897 4097 81909 4131
rect 81943 4128 81955 4131
rect 83090 4128 83096 4140
rect 81943 4100 83096 4128
rect 81943 4097 81955 4100
rect 81897 4091 81955 4097
rect 83090 4088 83096 4100
rect 83148 4088 83154 4140
rect 83826 4128 83832 4140
rect 83787 4100 83832 4128
rect 83826 4088 83832 4100
rect 83884 4088 83890 4140
rect 65150 4020 65156 4072
rect 65208 4060 65214 4072
rect 69198 4060 69204 4072
rect 65208 4032 69204 4060
rect 65208 4020 65214 4032
rect 69198 4020 69204 4032
rect 69256 4060 69262 4072
rect 69385 4063 69443 4069
rect 69385 4060 69397 4063
rect 69256 4032 69397 4060
rect 69256 4020 69262 4032
rect 69385 4029 69397 4032
rect 69431 4029 69443 4063
rect 69661 4063 69719 4069
rect 69661 4060 69673 4063
rect 69385 4023 69443 4029
rect 69492 4032 69673 4060
rect 65061 3995 65119 4001
rect 64524 3964 64920 3992
rect 28040 3896 29684 3924
rect 28040 3884 28046 3896
rect 30282 3884 30288 3936
rect 30340 3924 30346 3936
rect 30469 3927 30527 3933
rect 30469 3924 30481 3927
rect 30340 3896 30481 3924
rect 30340 3884 30346 3896
rect 30469 3893 30481 3896
rect 30515 3893 30527 3927
rect 31662 3924 31668 3936
rect 31623 3896 31668 3924
rect 30469 3887 30527 3893
rect 31662 3884 31668 3896
rect 31720 3884 31726 3936
rect 33318 3924 33324 3936
rect 33279 3896 33324 3924
rect 33318 3884 33324 3896
rect 33376 3884 33382 3936
rect 33870 3924 33876 3936
rect 33831 3896 33876 3924
rect 33870 3884 33876 3896
rect 33928 3884 33934 3936
rect 34238 3884 34244 3936
rect 34296 3924 34302 3936
rect 35161 3927 35219 3933
rect 35161 3924 35173 3927
rect 34296 3896 35173 3924
rect 34296 3884 34302 3896
rect 35161 3893 35173 3896
rect 35207 3893 35219 3927
rect 35161 3887 35219 3893
rect 36633 3927 36691 3933
rect 36633 3893 36645 3927
rect 36679 3924 36691 3927
rect 37734 3924 37740 3936
rect 36679 3896 37740 3924
rect 36679 3893 36691 3896
rect 36633 3887 36691 3893
rect 37734 3884 37740 3896
rect 37792 3884 37798 3936
rect 38289 3927 38347 3933
rect 38289 3893 38301 3927
rect 38335 3924 38347 3927
rect 38746 3924 38752 3936
rect 38335 3896 38752 3924
rect 38335 3893 38347 3896
rect 38289 3887 38347 3893
rect 38746 3884 38752 3896
rect 38804 3884 38810 3936
rect 39206 3924 39212 3936
rect 39167 3896 39212 3924
rect 39206 3884 39212 3896
rect 39264 3884 39270 3936
rect 39942 3924 39948 3936
rect 39903 3896 39948 3924
rect 39942 3884 39948 3896
rect 40000 3884 40006 3936
rect 40865 3927 40923 3933
rect 40865 3893 40877 3927
rect 40911 3924 40923 3927
rect 41138 3924 41144 3936
rect 40911 3896 41144 3924
rect 40911 3893 40923 3896
rect 40865 3887 40923 3893
rect 41138 3884 41144 3896
rect 41196 3884 41202 3936
rect 41874 3924 41880 3936
rect 41835 3896 41880 3924
rect 41874 3884 41880 3896
rect 41932 3884 41938 3936
rect 42797 3927 42855 3933
rect 42797 3893 42809 3927
rect 42843 3924 42855 3927
rect 42886 3924 42892 3936
rect 42843 3896 42892 3924
rect 42843 3893 42855 3896
rect 42797 3887 42855 3893
rect 42886 3884 42892 3896
rect 42944 3884 42950 3936
rect 43717 3927 43775 3933
rect 43717 3893 43729 3927
rect 43763 3924 43775 3927
rect 43898 3924 43904 3936
rect 43763 3896 43904 3924
rect 43763 3893 43775 3896
rect 43717 3887 43775 3893
rect 43898 3884 43904 3896
rect 43956 3884 43962 3936
rect 45094 3924 45100 3936
rect 45055 3896 45100 3924
rect 45094 3884 45100 3896
rect 45152 3884 45158 3936
rect 45462 3884 45468 3936
rect 45520 3924 45526 3936
rect 45557 3927 45615 3933
rect 45557 3924 45569 3927
rect 45520 3896 45569 3924
rect 45520 3884 45526 3896
rect 45557 3893 45569 3896
rect 45603 3893 45615 3927
rect 46198 3924 46204 3936
rect 46159 3896 46204 3924
rect 45557 3887 45615 3893
rect 46198 3884 46204 3896
rect 46256 3884 46262 3936
rect 46290 3884 46296 3936
rect 46348 3924 46354 3936
rect 46845 3927 46903 3933
rect 46845 3924 46857 3927
rect 46348 3896 46857 3924
rect 46348 3884 46354 3896
rect 46845 3893 46857 3896
rect 46891 3893 46903 3927
rect 46845 3887 46903 3893
rect 46934 3884 46940 3936
rect 46992 3924 46998 3936
rect 47765 3927 47823 3933
rect 47765 3924 47777 3927
rect 46992 3896 47777 3924
rect 46992 3884 46998 3896
rect 47765 3893 47777 3896
rect 47811 3893 47823 3927
rect 47765 3887 47823 3893
rect 50433 3927 50491 3933
rect 50433 3893 50445 3927
rect 50479 3924 50491 3927
rect 50614 3924 50620 3936
rect 50479 3896 50620 3924
rect 50479 3893 50491 3896
rect 50433 3887 50491 3893
rect 50614 3884 50620 3896
rect 50672 3884 50678 3936
rect 50890 3924 50896 3936
rect 50851 3896 50896 3924
rect 50890 3884 50896 3896
rect 50948 3884 50954 3936
rect 51534 3924 51540 3936
rect 51495 3896 51540 3924
rect 51534 3884 51540 3896
rect 51592 3884 51598 3936
rect 52270 3924 52276 3936
rect 52231 3896 52276 3924
rect 52270 3884 52276 3896
rect 52328 3884 52334 3936
rect 54018 3924 54024 3936
rect 53979 3896 54024 3924
rect 54018 3884 54024 3896
rect 54076 3924 54082 3936
rect 54573 3927 54631 3933
rect 54573 3924 54585 3927
rect 54076 3896 54585 3924
rect 54076 3884 54082 3896
rect 54573 3893 54585 3896
rect 54619 3893 54631 3927
rect 54573 3887 54631 3893
rect 55214 3884 55220 3936
rect 55272 3924 55278 3936
rect 55272 3896 55317 3924
rect 55272 3884 55278 3896
rect 56594 3884 56600 3936
rect 56652 3924 56658 3936
rect 57149 3927 57207 3933
rect 57149 3924 57161 3927
rect 56652 3896 57161 3924
rect 56652 3884 56658 3896
rect 57149 3893 57161 3896
rect 57195 3893 57207 3927
rect 57149 3887 57207 3893
rect 59173 3927 59231 3933
rect 59173 3893 59185 3927
rect 59219 3924 59231 3927
rect 59630 3924 59636 3936
rect 59219 3896 59636 3924
rect 59219 3893 59231 3896
rect 59173 3887 59231 3893
rect 59630 3884 59636 3896
rect 59688 3884 59694 3936
rect 61378 3924 61384 3936
rect 61339 3896 61384 3924
rect 61378 3884 61384 3896
rect 61436 3884 61442 3936
rect 63218 3884 63224 3936
rect 63276 3924 63282 3936
rect 63497 3927 63555 3933
rect 63497 3924 63509 3927
rect 63276 3896 63509 3924
rect 63276 3884 63282 3896
rect 63497 3893 63509 3896
rect 63543 3893 63555 3927
rect 64892 3924 64920 3964
rect 65061 3961 65073 3995
rect 65107 3961 65119 3995
rect 65334 3992 65340 4004
rect 65061 3955 65119 3961
rect 65168 3964 65340 3992
rect 65168 3924 65196 3964
rect 65334 3952 65340 3964
rect 65392 3992 65398 4004
rect 67358 3992 67364 4004
rect 65392 3964 67364 3992
rect 65392 3952 65398 3964
rect 67358 3952 67364 3964
rect 67416 3952 67422 4004
rect 68925 3995 68983 4001
rect 68925 3961 68937 3995
rect 68971 3992 68983 3995
rect 69492 3992 69520 4032
rect 69661 4029 69673 4032
rect 69707 4029 69719 4063
rect 69661 4023 69719 4029
rect 69750 4020 69756 4072
rect 69808 4060 69814 4072
rect 72329 4063 72387 4069
rect 72329 4060 72341 4063
rect 69808 4032 72341 4060
rect 69808 4020 69814 4032
rect 72329 4029 72341 4032
rect 72375 4060 72387 4063
rect 72418 4060 72424 4072
rect 72375 4032 72424 4060
rect 72375 4029 72387 4032
rect 72329 4023 72387 4029
rect 72418 4020 72424 4032
rect 72476 4020 72482 4072
rect 72510 4020 72516 4072
rect 72568 4060 72574 4072
rect 79134 4060 79140 4072
rect 72568 4032 78996 4060
rect 79095 4032 79140 4060
rect 72568 4020 72574 4032
rect 73522 3992 73528 4004
rect 68971 3964 69520 3992
rect 70688 3964 73528 3992
rect 68971 3961 68983 3964
rect 68925 3955 68983 3961
rect 65518 3924 65524 3936
rect 64892 3896 65196 3924
rect 65479 3896 65524 3924
rect 63497 3887 63555 3893
rect 65518 3884 65524 3896
rect 65576 3884 65582 3936
rect 66441 3927 66499 3933
rect 66441 3893 66453 3927
rect 66487 3924 66499 3927
rect 66530 3924 66536 3936
rect 66487 3896 66536 3924
rect 66487 3893 66499 3896
rect 66441 3887 66499 3893
rect 66530 3884 66536 3896
rect 66588 3884 66594 3936
rect 67821 3927 67879 3933
rect 67821 3893 67833 3927
rect 67867 3924 67879 3927
rect 68462 3924 68468 3936
rect 67867 3896 68468 3924
rect 67867 3893 67879 3896
rect 67821 3887 67879 3893
rect 68462 3884 68468 3896
rect 68520 3884 68526 3936
rect 69198 3884 69204 3936
rect 69256 3924 69262 3936
rect 70688 3924 70716 3964
rect 73522 3952 73528 3964
rect 73580 3952 73586 4004
rect 77110 3992 77116 4004
rect 75380 3964 77116 3992
rect 75380 3936 75408 3964
rect 77110 3952 77116 3964
rect 77168 3992 77174 4004
rect 78674 3992 78680 4004
rect 77168 3964 78680 3992
rect 77168 3952 77174 3964
rect 78674 3952 78680 3964
rect 78732 3952 78738 4004
rect 69256 3896 70716 3924
rect 71133 3927 71191 3933
rect 69256 3884 69262 3896
rect 71133 3893 71145 3927
rect 71179 3924 71191 3927
rect 71222 3924 71228 3936
rect 71179 3896 71228 3924
rect 71179 3893 71191 3896
rect 71133 3887 71191 3893
rect 71222 3884 71228 3896
rect 71280 3884 71286 3936
rect 71590 3884 71596 3936
rect 71648 3924 71654 3936
rect 74629 3927 74687 3933
rect 74629 3924 74641 3927
rect 71648 3896 74641 3924
rect 71648 3884 71654 3896
rect 74629 3893 74641 3896
rect 74675 3924 74687 3927
rect 75362 3924 75368 3936
rect 74675 3896 75368 3924
rect 74675 3893 74687 3896
rect 74629 3887 74687 3893
rect 75362 3884 75368 3896
rect 75420 3884 75426 3936
rect 76466 3884 76472 3936
rect 76524 3924 76530 3936
rect 76561 3927 76619 3933
rect 76561 3924 76573 3927
rect 76524 3896 76573 3924
rect 76524 3884 76530 3896
rect 76561 3893 76573 3896
rect 76607 3893 76619 3927
rect 76561 3887 76619 3893
rect 78125 3927 78183 3933
rect 78125 3893 78137 3927
rect 78171 3924 78183 3927
rect 78766 3924 78772 3936
rect 78171 3896 78772 3924
rect 78171 3893 78183 3896
rect 78125 3887 78183 3893
rect 78766 3884 78772 3896
rect 78824 3884 78830 3936
rect 78968 3924 78996 4032
rect 79134 4020 79140 4032
rect 79192 4020 79198 4072
rect 79778 4020 79784 4072
rect 79836 4060 79842 4072
rect 81986 4060 81992 4072
rect 79836 4032 81992 4060
rect 79836 4020 79842 4032
rect 81986 4020 81992 4032
rect 82044 4060 82050 4072
rect 82998 4060 83004 4072
rect 82044 4032 83004 4060
rect 82044 4020 82050 4032
rect 82998 4020 83004 4032
rect 83056 4060 83062 4072
rect 83185 4063 83243 4069
rect 83185 4060 83197 4063
rect 83056 4032 83197 4060
rect 83056 4020 83062 4032
rect 83185 4029 83197 4032
rect 83231 4060 83243 4063
rect 83642 4060 83648 4072
rect 83231 4032 83648 4060
rect 83231 4029 83243 4032
rect 83185 4023 83243 4029
rect 83642 4020 83648 4032
rect 83700 4020 83706 4072
rect 80885 3995 80943 4001
rect 80885 3961 80897 3995
rect 80931 3992 80943 3995
rect 82722 3992 82728 4004
rect 80931 3964 82728 3992
rect 80931 3961 80943 3964
rect 80885 3955 80943 3961
rect 82722 3952 82728 3964
rect 82780 3992 82786 4004
rect 82780 3964 93854 3992
rect 82780 3952 82786 3964
rect 81434 3924 81440 3936
rect 78968 3896 81440 3924
rect 81434 3884 81440 3896
rect 81492 3884 81498 3936
rect 83458 3884 83464 3936
rect 83516 3924 83522 3936
rect 84381 3927 84439 3933
rect 84381 3924 84393 3927
rect 83516 3896 84393 3924
rect 83516 3884 83522 3896
rect 84381 3893 84393 3896
rect 84427 3893 84439 3927
rect 93826 3924 93854 3964
rect 117222 3924 117228 3936
rect 93826 3896 117228 3924
rect 84381 3887 84439 3893
rect 117222 3884 117228 3896
rect 117280 3884 117286 3936
rect 1104 3834 148856 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 65654 3834
rect 65706 3782 65718 3834
rect 65770 3782 65782 3834
rect 65834 3782 65846 3834
rect 65898 3782 65910 3834
rect 65962 3782 96374 3834
rect 96426 3782 96438 3834
rect 96490 3782 96502 3834
rect 96554 3782 96566 3834
rect 96618 3782 96630 3834
rect 96682 3782 127094 3834
rect 127146 3782 127158 3834
rect 127210 3782 127222 3834
rect 127274 3782 127286 3834
rect 127338 3782 127350 3834
rect 127402 3782 148856 3834
rect 1104 3760 148856 3782
rect 8573 3723 8631 3729
rect 8573 3689 8585 3723
rect 8619 3720 8631 3723
rect 22738 3720 22744 3732
rect 8619 3692 22600 3720
rect 22699 3692 22744 3720
rect 8619 3689 8631 3692
rect 8573 3683 8631 3689
rect 7006 3584 7012 3596
rect 6288 3556 7012 3584
rect 6288 3528 6316 3556
rect 7006 3544 7012 3556
rect 7064 3584 7070 3596
rect 7064 3556 8064 3584
rect 7064 3544 7070 3556
rect 4893 3519 4951 3525
rect 4893 3485 4905 3519
rect 4939 3516 4951 3519
rect 5258 3516 5264 3528
rect 4939 3488 5264 3516
rect 4939 3485 4951 3488
rect 4893 3479 4951 3485
rect 5258 3476 5264 3488
rect 5316 3516 5322 3528
rect 5353 3519 5411 3525
rect 5353 3516 5365 3519
rect 5316 3488 5365 3516
rect 5316 3476 5322 3488
rect 5353 3485 5365 3488
rect 5399 3485 5411 3519
rect 6270 3516 6276 3528
rect 6231 3488 6276 3516
rect 5353 3479 5411 3485
rect 6270 3476 6276 3488
rect 6328 3476 6334 3528
rect 6638 3476 6644 3528
rect 6696 3516 6702 3528
rect 8036 3525 8064 3556
rect 6917 3519 6975 3525
rect 6917 3516 6929 3519
rect 6696 3488 6929 3516
rect 6696 3476 6702 3488
rect 6917 3485 6929 3488
rect 6963 3485 6975 3519
rect 6917 3479 6975 3485
rect 8021 3519 8079 3525
rect 8021 3485 8033 3519
rect 8067 3516 8079 3519
rect 8588 3516 8616 3683
rect 22572 3652 22600 3692
rect 22738 3680 22744 3692
rect 22796 3680 22802 3732
rect 23934 3720 23940 3732
rect 23032 3692 23796 3720
rect 23895 3692 23940 3720
rect 23032 3652 23060 3692
rect 22572 3624 23060 3652
rect 23768 3652 23796 3692
rect 23934 3680 23940 3692
rect 23992 3680 23998 3732
rect 24670 3720 24676 3732
rect 24631 3692 24676 3720
rect 24670 3680 24676 3692
rect 24728 3680 24734 3732
rect 30193 3723 30251 3729
rect 30193 3720 30205 3723
rect 26344 3692 30205 3720
rect 26344 3652 26372 3692
rect 30193 3689 30205 3692
rect 30239 3689 30251 3723
rect 33134 3720 33140 3732
rect 33095 3692 33140 3720
rect 30193 3683 30251 3689
rect 23768 3624 26372 3652
rect 27522 3612 27528 3664
rect 27580 3652 27586 3664
rect 27982 3652 27988 3664
rect 27580 3624 27988 3652
rect 27580 3612 27586 3624
rect 27982 3612 27988 3624
rect 28040 3612 28046 3664
rect 28718 3612 28724 3664
rect 28776 3652 28782 3664
rect 28997 3655 29055 3661
rect 28997 3652 29009 3655
rect 28776 3624 29009 3652
rect 28776 3612 28782 3624
rect 28997 3621 29009 3624
rect 29043 3621 29055 3655
rect 30208 3652 30236 3683
rect 33134 3680 33140 3692
rect 33192 3680 33198 3732
rect 40218 3720 40224 3732
rect 40179 3692 40224 3720
rect 40218 3680 40224 3692
rect 40276 3680 40282 3732
rect 40954 3720 40960 3732
rect 40915 3692 40960 3720
rect 40954 3680 40960 3692
rect 41012 3680 41018 3732
rect 43806 3720 43812 3732
rect 43767 3692 43812 3720
rect 43806 3680 43812 3692
rect 43864 3680 43870 3732
rect 46106 3680 46112 3732
rect 46164 3720 46170 3732
rect 46164 3692 51120 3720
rect 46164 3680 46170 3692
rect 36909 3655 36967 3661
rect 30208 3624 30328 3652
rect 28997 3615 29055 3621
rect 9398 3544 9404 3596
rect 9456 3584 9462 3596
rect 22002 3584 22008 3596
rect 9456 3556 22008 3584
rect 9456 3544 9462 3556
rect 22002 3544 22008 3556
rect 22060 3544 22066 3596
rect 23290 3544 23296 3596
rect 23348 3584 23354 3596
rect 23385 3587 23443 3593
rect 23385 3584 23397 3587
rect 23348 3556 23397 3584
rect 23348 3544 23354 3556
rect 23385 3553 23397 3556
rect 23431 3584 23443 3587
rect 24946 3584 24952 3596
rect 23431 3556 24952 3584
rect 23431 3553 23443 3556
rect 23385 3547 23443 3553
rect 24946 3544 24952 3556
rect 25004 3544 25010 3596
rect 26234 3584 26240 3596
rect 26195 3556 26240 3584
rect 26234 3544 26240 3556
rect 26292 3544 26298 3596
rect 26513 3587 26571 3593
rect 26513 3553 26525 3587
rect 26559 3584 26571 3587
rect 27154 3584 27160 3596
rect 26559 3556 27160 3584
rect 26559 3553 26571 3556
rect 26513 3547 26571 3553
rect 27154 3544 27160 3556
rect 27212 3544 27218 3596
rect 27890 3584 27896 3596
rect 27632 3556 27896 3584
rect 8067 3488 8616 3516
rect 21453 3519 21511 3525
rect 8067 3485 8079 3488
rect 8021 3479 8079 3485
rect 21453 3485 21465 3519
rect 21499 3485 21511 3519
rect 22094 3516 22100 3528
rect 22007 3488 22100 3516
rect 21453 3479 21511 3485
rect 5626 3408 5632 3460
rect 5684 3448 5690 3460
rect 6181 3451 6239 3457
rect 6181 3448 6193 3451
rect 5684 3420 6193 3448
rect 5684 3408 5690 3420
rect 6181 3417 6193 3420
rect 6227 3417 6239 3451
rect 21468 3448 21496 3479
rect 22094 3476 22100 3488
rect 22152 3516 22158 3528
rect 25866 3516 25872 3528
rect 22152 3488 25872 3516
rect 22152 3476 22158 3488
rect 25866 3476 25872 3488
rect 25924 3476 25930 3528
rect 27632 3502 27660 3556
rect 27890 3544 27896 3556
rect 27948 3544 27954 3596
rect 28074 3544 28080 3596
rect 28132 3584 28138 3596
rect 30190 3584 30196 3596
rect 28132 3556 30196 3584
rect 28132 3544 28138 3556
rect 30190 3544 30196 3556
rect 30248 3544 30254 3596
rect 28813 3519 28871 3525
rect 28813 3485 28825 3519
rect 28859 3485 28871 3519
rect 30300 3516 30328 3624
rect 36909 3621 36921 3655
rect 36955 3652 36967 3655
rect 38562 3652 38568 3664
rect 36955 3624 38568 3652
rect 36955 3621 36967 3624
rect 36909 3615 36967 3621
rect 30374 3544 30380 3596
rect 30432 3584 30438 3596
rect 35710 3584 35716 3596
rect 30432 3556 34284 3584
rect 35671 3556 35716 3584
rect 30432 3544 30438 3556
rect 30745 3519 30803 3525
rect 30745 3516 30757 3519
rect 30300 3488 30757 3516
rect 28813 3479 28871 3485
rect 30745 3485 30757 3488
rect 30791 3516 30803 3519
rect 32766 3516 32772 3528
rect 30791 3488 32772 3516
rect 30791 3485 30803 3488
rect 30745 3479 30803 3485
rect 24210 3448 24216 3460
rect 21468 3420 24216 3448
rect 6181 3411 6239 3417
rect 24210 3408 24216 3420
rect 24268 3408 24274 3460
rect 5537 3383 5595 3389
rect 5537 3349 5549 3383
rect 5583 3380 5595 3383
rect 5718 3380 5724 3392
rect 5583 3352 5724 3380
rect 5583 3349 5595 3352
rect 5537 3343 5595 3349
rect 5718 3340 5724 3352
rect 5776 3340 5782 3392
rect 6730 3380 6736 3392
rect 6691 3352 6736 3380
rect 6730 3340 6736 3352
rect 6788 3340 6794 3392
rect 7926 3380 7932 3392
rect 7887 3352 7932 3380
rect 7926 3340 7932 3352
rect 7984 3340 7990 3392
rect 9214 3380 9220 3392
rect 9175 3352 9220 3380
rect 9214 3340 9220 3352
rect 9272 3340 9278 3392
rect 20438 3380 20444 3392
rect 20399 3352 20444 3380
rect 20438 3340 20444 3352
rect 20496 3340 20502 3392
rect 20990 3380 20996 3392
rect 20951 3352 20996 3380
rect 20990 3340 20996 3352
rect 21048 3340 21054 3392
rect 21634 3380 21640 3392
rect 21595 3352 21640 3380
rect 21634 3340 21640 3352
rect 21692 3340 21698 3392
rect 22189 3383 22247 3389
rect 22189 3349 22201 3383
rect 22235 3380 22247 3383
rect 22738 3380 22744 3392
rect 22235 3352 22744 3380
rect 22235 3349 22247 3352
rect 22189 3343 22247 3349
rect 22738 3340 22744 3352
rect 22796 3340 22802 3392
rect 23014 3340 23020 3392
rect 23072 3380 23078 3392
rect 23109 3383 23167 3389
rect 23109 3380 23121 3383
rect 23072 3352 23121 3380
rect 23072 3340 23078 3352
rect 23109 3349 23121 3352
rect 23155 3349 23167 3383
rect 23109 3343 23167 3349
rect 23201 3383 23259 3389
rect 23201 3349 23213 3383
rect 23247 3380 23259 3383
rect 23934 3380 23940 3392
rect 23247 3352 23940 3380
rect 23247 3349 23259 3352
rect 23201 3343 23259 3349
rect 23934 3340 23940 3352
rect 23992 3340 23998 3392
rect 24854 3340 24860 3392
rect 24912 3380 24918 3392
rect 25133 3383 25191 3389
rect 25133 3380 25145 3383
rect 24912 3352 25145 3380
rect 24912 3340 24918 3352
rect 25133 3349 25145 3352
rect 25179 3349 25191 3383
rect 25133 3343 25191 3349
rect 25777 3383 25835 3389
rect 25777 3349 25789 3383
rect 25823 3380 25835 3383
rect 26418 3380 26424 3392
rect 25823 3352 26424 3380
rect 25823 3349 25835 3352
rect 25777 3343 25835 3349
rect 26418 3340 26424 3352
rect 26476 3340 26482 3392
rect 27982 3340 27988 3392
rect 28040 3380 28046 3392
rect 28828 3380 28856 3479
rect 32766 3476 32772 3488
rect 32824 3476 32830 3528
rect 34149 3519 34207 3525
rect 34149 3485 34161 3519
rect 34195 3485 34207 3519
rect 34256 3516 34284 3556
rect 35710 3544 35716 3556
rect 35768 3544 35774 3596
rect 35805 3587 35863 3593
rect 35805 3553 35817 3587
rect 35851 3584 35863 3587
rect 35986 3584 35992 3596
rect 35851 3556 35992 3584
rect 35851 3553 35863 3556
rect 35805 3547 35863 3553
rect 35986 3544 35992 3556
rect 36044 3544 36050 3596
rect 36924 3516 36952 3615
rect 38562 3612 38568 3624
rect 38620 3612 38626 3664
rect 43346 3652 43352 3664
rect 43259 3624 43352 3652
rect 43346 3612 43352 3624
rect 43404 3652 43410 3664
rect 51092 3652 51120 3692
rect 51350 3680 51356 3732
rect 51408 3720 51414 3732
rect 51905 3723 51963 3729
rect 51905 3720 51917 3723
rect 51408 3692 51917 3720
rect 51408 3680 51414 3692
rect 51905 3689 51917 3692
rect 51951 3689 51963 3723
rect 51905 3683 51963 3689
rect 53282 3680 53288 3732
rect 53340 3720 53346 3732
rect 57422 3720 57428 3732
rect 53340 3692 55214 3720
rect 57383 3692 57428 3720
rect 53340 3680 53346 3692
rect 53926 3652 53932 3664
rect 43404 3624 45416 3652
rect 51092 3624 52040 3652
rect 53887 3624 53932 3652
rect 43404 3612 43410 3624
rect 41598 3584 41604 3596
rect 41559 3556 41604 3584
rect 41598 3544 41604 3556
rect 41656 3544 41662 3596
rect 41874 3584 41880 3596
rect 41835 3556 41880 3584
rect 41874 3544 41880 3556
rect 41932 3544 41938 3596
rect 43438 3544 43444 3596
rect 43496 3584 43502 3596
rect 44269 3587 44327 3593
rect 44269 3584 44281 3587
rect 43496 3556 44281 3584
rect 43496 3544 43502 3556
rect 44269 3553 44281 3556
rect 44315 3553 44327 3587
rect 44269 3547 44327 3553
rect 44361 3587 44419 3593
rect 44361 3553 44373 3587
rect 44407 3584 44419 3587
rect 45388 3584 45416 3624
rect 44407 3556 45324 3584
rect 45388 3556 51074 3584
rect 44407 3553 44419 3556
rect 44361 3547 44419 3553
rect 34256 3488 36952 3516
rect 34149 3479 34207 3485
rect 31941 3451 31999 3457
rect 31941 3417 31953 3451
rect 31987 3448 31999 3451
rect 32858 3448 32864 3460
rect 31987 3420 32864 3448
rect 31987 3417 31999 3420
rect 31941 3411 31999 3417
rect 32858 3408 32864 3420
rect 32916 3448 32922 3460
rect 33045 3451 33103 3457
rect 33045 3448 33057 3451
rect 32916 3420 33057 3448
rect 32916 3408 32922 3420
rect 33045 3417 33057 3420
rect 33091 3417 33103 3451
rect 34164 3448 34192 3479
rect 37090 3476 37096 3528
rect 37148 3516 37154 3528
rect 38657 3519 38715 3525
rect 38657 3516 38669 3519
rect 37148 3488 38669 3516
rect 37148 3476 37154 3488
rect 38657 3485 38669 3488
rect 38703 3485 38715 3519
rect 38657 3479 38715 3485
rect 42978 3476 42984 3528
rect 43036 3476 43042 3528
rect 44376 3516 44404 3547
rect 44008 3488 44404 3516
rect 35621 3451 35679 3457
rect 34164 3420 35296 3448
rect 33045 3411 33103 3417
rect 28040 3352 28856 3380
rect 28040 3340 28046 3352
rect 30742 3340 30748 3392
rect 30800 3380 30806 3392
rect 30837 3383 30895 3389
rect 30837 3380 30849 3383
rect 30800 3352 30849 3380
rect 30800 3340 30806 3352
rect 30837 3349 30849 3352
rect 30883 3349 30895 3383
rect 30837 3343 30895 3349
rect 32306 3340 32312 3392
rect 32364 3380 32370 3392
rect 32401 3383 32459 3389
rect 32401 3380 32413 3383
rect 32364 3352 32413 3380
rect 32364 3340 32370 3352
rect 32401 3349 32413 3352
rect 32447 3349 32459 3383
rect 32401 3343 32459 3349
rect 34333 3383 34391 3389
rect 34333 3349 34345 3383
rect 34379 3380 34391 3383
rect 34698 3380 34704 3392
rect 34379 3352 34704 3380
rect 34379 3349 34391 3352
rect 34333 3343 34391 3349
rect 34698 3340 34704 3352
rect 34756 3340 34762 3392
rect 35268 3389 35296 3420
rect 35621 3417 35633 3451
rect 35667 3417 35679 3451
rect 35621 3411 35679 3417
rect 35253 3383 35311 3389
rect 35253 3349 35265 3383
rect 35299 3349 35311 3383
rect 35636 3380 35664 3411
rect 35802 3408 35808 3460
rect 35860 3448 35866 3460
rect 36078 3448 36084 3460
rect 35860 3420 36084 3448
rect 35860 3408 35866 3420
rect 36078 3408 36084 3420
rect 36136 3408 36142 3460
rect 38194 3448 38200 3460
rect 38155 3420 38200 3448
rect 38194 3408 38200 3420
rect 38252 3408 38258 3460
rect 40129 3451 40187 3457
rect 40129 3417 40141 3451
rect 40175 3417 40187 3451
rect 40129 3411 40187 3417
rect 41049 3451 41107 3457
rect 41049 3417 41061 3451
rect 41095 3448 41107 3451
rect 41138 3448 41144 3460
rect 41095 3420 41144 3448
rect 41095 3417 41107 3420
rect 41049 3411 41107 3417
rect 37090 3380 37096 3392
rect 35636 3352 37096 3380
rect 35253 3343 35311 3349
rect 37090 3340 37096 3352
rect 37148 3340 37154 3392
rect 38378 3340 38384 3392
rect 38436 3380 38442 3392
rect 38841 3383 38899 3389
rect 38841 3380 38853 3383
rect 38436 3352 38853 3380
rect 38436 3340 38442 3352
rect 38841 3349 38853 3352
rect 38887 3349 38899 3383
rect 38841 3343 38899 3349
rect 39485 3383 39543 3389
rect 39485 3349 39497 3383
rect 39531 3380 39543 3383
rect 39758 3380 39764 3392
rect 39531 3352 39764 3380
rect 39531 3349 39543 3352
rect 39485 3343 39543 3349
rect 39758 3340 39764 3352
rect 39816 3380 39822 3392
rect 40144 3380 40172 3411
rect 41138 3408 41144 3420
rect 41196 3408 41202 3460
rect 39816 3352 40172 3380
rect 39816 3340 39822 3352
rect 42518 3340 42524 3392
rect 42576 3380 42582 3392
rect 44008 3380 44036 3488
rect 45094 3476 45100 3528
rect 45152 3516 45158 3528
rect 45189 3519 45247 3525
rect 45189 3516 45201 3519
rect 45152 3488 45201 3516
rect 45152 3476 45158 3488
rect 45189 3485 45201 3488
rect 45235 3485 45247 3519
rect 45296 3516 45324 3556
rect 45922 3516 45928 3528
rect 45296 3488 45928 3516
rect 45189 3479 45247 3485
rect 45922 3476 45928 3488
rect 45980 3476 45986 3528
rect 46201 3519 46259 3525
rect 46201 3485 46213 3519
rect 46247 3516 46259 3519
rect 46750 3516 46756 3528
rect 46247 3488 46756 3516
rect 46247 3485 46259 3488
rect 46201 3479 46259 3485
rect 46750 3476 46756 3488
rect 46808 3476 46814 3528
rect 46842 3476 46848 3528
rect 46900 3516 46906 3528
rect 49050 3516 49056 3528
rect 46900 3488 46945 3516
rect 49011 3488 49056 3516
rect 46900 3476 46906 3488
rect 49050 3476 49056 3488
rect 49108 3476 49114 3528
rect 49326 3516 49332 3528
rect 49287 3488 49332 3516
rect 49326 3476 49332 3488
rect 49384 3476 49390 3528
rect 50893 3519 50951 3525
rect 50893 3485 50905 3519
rect 50939 3485 50951 3519
rect 50893 3479 50951 3485
rect 44174 3448 44180 3460
rect 44087 3420 44180 3448
rect 44174 3408 44180 3420
rect 44232 3448 44238 3460
rect 50908 3448 50936 3479
rect 44232 3420 50936 3448
rect 51046 3448 51074 3556
rect 51902 3448 51908 3460
rect 51046 3420 51908 3448
rect 44232 3408 44238 3420
rect 51902 3408 51908 3420
rect 51960 3408 51966 3460
rect 45278 3380 45284 3392
rect 42576 3352 44036 3380
rect 45239 3352 45284 3380
rect 42576 3340 42582 3352
rect 45278 3340 45284 3352
rect 45336 3340 45342 3392
rect 46385 3383 46443 3389
rect 46385 3349 46397 3383
rect 46431 3380 46443 3383
rect 47670 3380 47676 3392
rect 46431 3352 47676 3380
rect 46431 3349 46443 3352
rect 46385 3343 46443 3349
rect 47670 3340 47676 3352
rect 47728 3340 47734 3392
rect 47762 3340 47768 3392
rect 47820 3380 47826 3392
rect 48133 3383 48191 3389
rect 48133 3380 48145 3383
rect 47820 3352 48145 3380
rect 47820 3340 47826 3352
rect 48133 3349 48145 3352
rect 48179 3380 48191 3383
rect 50341 3383 50399 3389
rect 50341 3380 50353 3383
rect 48179 3352 50353 3380
rect 48179 3349 48191 3352
rect 48133 3343 48191 3349
rect 50341 3349 50353 3352
rect 50387 3380 50399 3383
rect 50614 3380 50620 3392
rect 50387 3352 50620 3380
rect 50387 3349 50399 3352
rect 50341 3343 50399 3349
rect 50614 3340 50620 3352
rect 50672 3340 50678 3392
rect 50798 3340 50804 3392
rect 50856 3380 50862 3392
rect 51077 3383 51135 3389
rect 51077 3380 51089 3383
rect 50856 3352 51089 3380
rect 50856 3340 50862 3352
rect 51077 3349 51089 3352
rect 51123 3349 51135 3383
rect 52012 3380 52040 3624
rect 53926 3612 53932 3624
rect 53984 3612 53990 3664
rect 55186 3652 55214 3692
rect 57422 3680 57428 3692
rect 57480 3680 57486 3732
rect 57698 3680 57704 3732
rect 57756 3720 57762 3732
rect 57756 3692 65012 3720
rect 57756 3680 57762 3692
rect 63313 3655 63371 3661
rect 63313 3652 63325 3655
rect 55186 3624 62252 3652
rect 52086 3544 52092 3596
rect 52144 3584 52150 3596
rect 52365 3587 52423 3593
rect 52365 3584 52377 3587
rect 52144 3556 52377 3584
rect 52144 3544 52150 3556
rect 52365 3553 52377 3556
rect 52411 3553 52423 3587
rect 52365 3547 52423 3553
rect 52549 3587 52607 3593
rect 52549 3553 52561 3587
rect 52595 3584 52607 3587
rect 54202 3584 54208 3596
rect 52595 3556 54208 3584
rect 52595 3553 52607 3556
rect 52549 3547 52607 3553
rect 54202 3544 54208 3556
rect 54260 3544 54266 3596
rect 54312 3556 55076 3584
rect 52273 3519 52331 3525
rect 52273 3485 52285 3519
rect 52319 3516 52331 3519
rect 52454 3516 52460 3528
rect 52319 3488 52460 3516
rect 52319 3485 52331 3488
rect 52273 3479 52331 3485
rect 52454 3476 52460 3488
rect 52512 3516 52518 3528
rect 53006 3516 53012 3528
rect 52512 3488 53012 3516
rect 52512 3476 52518 3488
rect 53006 3476 53012 3488
rect 53064 3516 53070 3528
rect 54312 3516 54340 3556
rect 53064 3488 54340 3516
rect 54941 3519 54999 3525
rect 53064 3476 53070 3488
rect 54941 3485 54953 3519
rect 54987 3485 54999 3519
rect 54941 3479 54999 3485
rect 53193 3451 53251 3457
rect 53193 3417 53205 3451
rect 53239 3448 53251 3451
rect 53558 3448 53564 3460
rect 53239 3420 53564 3448
rect 53239 3417 53251 3420
rect 53193 3411 53251 3417
rect 53558 3408 53564 3420
rect 53616 3448 53622 3460
rect 53745 3451 53803 3457
rect 53745 3448 53757 3451
rect 53616 3420 53757 3448
rect 53616 3408 53622 3420
rect 53745 3417 53757 3420
rect 53791 3417 53803 3451
rect 53745 3411 53803 3417
rect 54294 3380 54300 3392
rect 52012 3352 54300 3380
rect 51077 3343 51135 3349
rect 54294 3340 54300 3352
rect 54352 3340 54358 3392
rect 54570 3340 54576 3392
rect 54628 3380 54634 3392
rect 54757 3383 54815 3389
rect 54757 3380 54769 3383
rect 54628 3352 54769 3380
rect 54628 3340 54634 3352
rect 54757 3349 54769 3352
rect 54803 3349 54815 3383
rect 54956 3380 54984 3479
rect 55048 3448 55076 3556
rect 55858 3544 55864 3596
rect 55916 3584 55922 3596
rect 56413 3587 56471 3593
rect 56413 3584 56425 3587
rect 55916 3556 56425 3584
rect 55916 3544 55922 3556
rect 56413 3553 56425 3556
rect 56459 3553 56471 3587
rect 56413 3547 56471 3553
rect 56505 3587 56563 3593
rect 56505 3553 56517 3587
rect 56551 3584 56563 3587
rect 57977 3587 58035 3593
rect 57977 3584 57989 3587
rect 56551 3556 57989 3584
rect 56551 3553 56563 3556
rect 56505 3547 56563 3553
rect 57977 3553 57989 3556
rect 58023 3584 58035 3587
rect 58618 3584 58624 3596
rect 58023 3556 58624 3584
rect 58023 3553 58035 3556
rect 57977 3547 58035 3553
rect 55122 3476 55128 3528
rect 55180 3516 55186 3528
rect 56520 3516 56548 3547
rect 58618 3544 58624 3556
rect 58676 3584 58682 3596
rect 61102 3584 61108 3596
rect 58676 3556 60964 3584
rect 61063 3556 61108 3584
rect 58676 3544 58682 3556
rect 55180 3488 56548 3516
rect 55180 3476 55186 3488
rect 57146 3476 57152 3528
rect 57204 3516 57210 3528
rect 59173 3519 59231 3525
rect 59173 3516 59185 3519
rect 57204 3488 59185 3516
rect 57204 3476 57210 3488
rect 59173 3485 59185 3488
rect 59219 3485 59231 3519
rect 59173 3479 59231 3485
rect 60093 3519 60151 3525
rect 60093 3485 60105 3519
rect 60139 3516 60151 3519
rect 60936 3516 60964 3556
rect 61102 3544 61108 3556
rect 61160 3544 61166 3596
rect 61197 3587 61255 3593
rect 61197 3553 61209 3587
rect 61243 3553 61255 3587
rect 61197 3547 61255 3553
rect 61212 3516 61240 3547
rect 62022 3516 62028 3528
rect 60139 3488 60688 3516
rect 60936 3488 61884 3516
rect 61983 3488 62028 3516
rect 60139 3485 60151 3488
rect 60093 3479 60151 3485
rect 57698 3448 57704 3460
rect 55048 3420 57704 3448
rect 57698 3408 57704 3420
rect 57756 3408 57762 3460
rect 57885 3451 57943 3457
rect 57885 3417 57897 3451
rect 57931 3448 57943 3451
rect 57974 3448 57980 3460
rect 57931 3420 57980 3448
rect 57931 3417 57943 3420
rect 57885 3411 57943 3417
rect 57974 3408 57980 3420
rect 58032 3408 58038 3460
rect 55953 3383 56011 3389
rect 55953 3380 55965 3383
rect 54956 3352 55965 3380
rect 54757 3343 54815 3349
rect 55953 3349 55965 3352
rect 55999 3349 56011 3383
rect 55953 3343 56011 3349
rect 56042 3340 56048 3392
rect 56100 3380 56106 3392
rect 56321 3383 56379 3389
rect 56321 3380 56333 3383
rect 56100 3352 56333 3380
rect 56100 3340 56106 3352
rect 56321 3349 56333 3352
rect 56367 3380 56379 3383
rect 56410 3380 56416 3392
rect 56367 3352 56416 3380
rect 56367 3349 56379 3352
rect 56321 3343 56379 3349
rect 56410 3340 56416 3352
rect 56468 3340 56474 3392
rect 57422 3340 57428 3392
rect 57480 3380 57486 3392
rect 57790 3380 57796 3392
rect 57480 3352 57796 3380
rect 57480 3340 57486 3352
rect 57790 3340 57796 3352
rect 57848 3340 57854 3392
rect 58710 3380 58716 3392
rect 58671 3352 58716 3380
rect 58710 3340 58716 3352
rect 58768 3340 58774 3392
rect 59078 3340 59084 3392
rect 59136 3380 59142 3392
rect 59357 3383 59415 3389
rect 59357 3380 59369 3383
rect 59136 3352 59369 3380
rect 59136 3340 59142 3352
rect 59357 3349 59369 3352
rect 59403 3349 59415 3383
rect 59357 3343 59415 3349
rect 59909 3383 59967 3389
rect 59909 3349 59921 3383
rect 59955 3380 59967 3383
rect 59998 3380 60004 3392
rect 59955 3352 60004 3380
rect 59955 3349 59967 3352
rect 59909 3343 59967 3349
rect 59998 3340 60004 3352
rect 60056 3340 60062 3392
rect 60660 3389 60688 3488
rect 61013 3451 61071 3457
rect 61013 3417 61025 3451
rect 61059 3448 61071 3451
rect 61470 3448 61476 3460
rect 61059 3420 61476 3448
rect 61059 3417 61071 3420
rect 61013 3411 61071 3417
rect 61470 3408 61476 3420
rect 61528 3408 61534 3460
rect 61856 3448 61884 3488
rect 62022 3476 62028 3488
rect 62080 3476 62086 3528
rect 62224 3516 62252 3624
rect 62408 3624 63325 3652
rect 62408 3516 62436 3624
rect 63313 3621 63325 3624
rect 63359 3621 63371 3655
rect 64984 3652 65012 3692
rect 65058 3680 65064 3732
rect 65116 3720 65122 3732
rect 65245 3723 65303 3729
rect 65245 3720 65257 3723
rect 65116 3692 65257 3720
rect 65116 3680 65122 3692
rect 65245 3689 65257 3692
rect 65291 3689 65303 3723
rect 65245 3683 65303 3689
rect 66438 3680 66444 3732
rect 66496 3720 66502 3732
rect 68830 3720 68836 3732
rect 66496 3692 67404 3720
rect 68791 3692 68836 3720
rect 66496 3680 66502 3692
rect 63313 3615 63371 3621
rect 63420 3624 63908 3652
rect 64984 3624 66668 3652
rect 62574 3544 62580 3596
rect 62632 3584 62638 3596
rect 63420 3584 63448 3624
rect 63880 3596 63908 3624
rect 62632 3556 63448 3584
rect 62632 3544 62638 3556
rect 63494 3544 63500 3596
rect 63552 3584 63558 3596
rect 63773 3587 63831 3593
rect 63773 3584 63785 3587
rect 63552 3556 63785 3584
rect 63552 3544 63558 3556
rect 63773 3553 63785 3556
rect 63819 3553 63831 3587
rect 63773 3547 63831 3553
rect 63862 3544 63868 3596
rect 63920 3584 63926 3596
rect 64601 3587 64659 3593
rect 64601 3584 64613 3587
rect 63920 3556 64613 3584
rect 63920 3544 63926 3556
rect 64601 3553 64613 3556
rect 64647 3553 64659 3587
rect 64601 3547 64659 3553
rect 64785 3587 64843 3593
rect 64785 3553 64797 3587
rect 64831 3584 64843 3587
rect 65426 3584 65432 3596
rect 64831 3556 65432 3584
rect 64831 3553 64843 3556
rect 64785 3547 64843 3553
rect 65426 3544 65432 3556
rect 65484 3544 65490 3596
rect 66438 3584 66444 3596
rect 66399 3556 66444 3584
rect 66438 3544 66444 3556
rect 66496 3544 66502 3596
rect 62485 3519 62543 3525
rect 62485 3516 62497 3519
rect 62224 3488 62344 3516
rect 62408 3488 62497 3516
rect 62316 3448 62344 3488
rect 62485 3485 62497 3488
rect 62531 3485 62543 3519
rect 62485 3479 62543 3485
rect 63681 3519 63739 3525
rect 63681 3485 63693 3519
rect 63727 3485 63739 3519
rect 64874 3516 64880 3528
rect 64835 3488 64880 3516
rect 63681 3479 63739 3485
rect 63696 3448 63724 3479
rect 64874 3476 64880 3488
rect 64932 3476 64938 3528
rect 66162 3476 66168 3528
rect 66220 3516 66226 3528
rect 66257 3519 66315 3525
rect 66257 3516 66269 3519
rect 66220 3488 66269 3516
rect 66220 3476 66226 3488
rect 66257 3485 66269 3488
rect 66303 3485 66315 3519
rect 66257 3479 66315 3485
rect 65058 3448 65064 3460
rect 61856 3420 62252 3448
rect 62316 3420 63632 3448
rect 63696 3420 65064 3448
rect 60645 3383 60703 3389
rect 60645 3349 60657 3383
rect 60691 3349 60703 3383
rect 60645 3343 60703 3349
rect 61194 3340 61200 3392
rect 61252 3380 61258 3392
rect 61841 3383 61899 3389
rect 61841 3380 61853 3383
rect 61252 3352 61853 3380
rect 61252 3340 61258 3352
rect 61841 3349 61853 3352
rect 61887 3349 61899 3383
rect 62224 3380 62252 3420
rect 62574 3380 62580 3392
rect 62224 3352 62580 3380
rect 61841 3343 61899 3349
rect 62574 3340 62580 3352
rect 62632 3340 62638 3392
rect 62669 3383 62727 3389
rect 62669 3349 62681 3383
rect 62715 3380 62727 3383
rect 63494 3380 63500 3392
rect 62715 3352 63500 3380
rect 62715 3349 62727 3352
rect 62669 3343 62727 3349
rect 63494 3340 63500 3352
rect 63552 3340 63558 3392
rect 63604 3380 63632 3420
rect 65058 3408 65064 3420
rect 65116 3408 65122 3460
rect 66640 3448 66668 3624
rect 67376 3584 67404 3692
rect 68830 3680 68836 3692
rect 68888 3680 68894 3732
rect 69842 3680 69848 3732
rect 69900 3720 69906 3732
rect 70029 3723 70087 3729
rect 70029 3720 70041 3723
rect 69900 3692 70041 3720
rect 69900 3680 69906 3692
rect 70029 3689 70041 3692
rect 70075 3689 70087 3723
rect 70029 3683 70087 3689
rect 70118 3680 70124 3732
rect 70176 3720 70182 3732
rect 70176 3692 79824 3720
rect 70176 3680 70182 3692
rect 76466 3612 76472 3664
rect 76524 3652 76530 3664
rect 79796 3652 79824 3692
rect 80422 3680 80428 3732
rect 80480 3720 80486 3732
rect 81253 3723 81311 3729
rect 81253 3720 81265 3723
rect 80480 3692 81265 3720
rect 80480 3680 80486 3692
rect 81253 3689 81265 3692
rect 81299 3689 81311 3723
rect 81253 3683 81311 3689
rect 81820 3692 82032 3720
rect 81820 3652 81848 3692
rect 76524 3624 78536 3652
rect 79796 3624 81848 3652
rect 82004 3652 82032 3692
rect 82078 3680 82084 3732
rect 82136 3720 82142 3732
rect 82449 3723 82507 3729
rect 82449 3720 82461 3723
rect 82136 3692 82461 3720
rect 82136 3680 82142 3692
rect 82449 3689 82461 3692
rect 82495 3689 82507 3723
rect 82449 3683 82507 3689
rect 82722 3680 82728 3732
rect 82780 3720 82786 3732
rect 84749 3723 84807 3729
rect 84749 3720 84761 3723
rect 82780 3692 84761 3720
rect 82780 3680 82786 3692
rect 84749 3689 84761 3692
rect 84795 3689 84807 3723
rect 84749 3683 84807 3689
rect 84838 3680 84844 3732
rect 84896 3720 84902 3732
rect 145926 3720 145932 3732
rect 84896 3692 145932 3720
rect 84896 3680 84902 3692
rect 145926 3680 145932 3692
rect 145984 3680 145990 3732
rect 104526 3652 104532 3664
rect 82004 3624 89714 3652
rect 76524 3612 76530 3624
rect 68002 3584 68008 3596
rect 67376 3556 68008 3584
rect 67376 3525 67404 3556
rect 68002 3544 68008 3556
rect 68060 3544 68066 3596
rect 68278 3584 68284 3596
rect 68239 3556 68284 3584
rect 68278 3544 68284 3556
rect 68336 3584 68342 3596
rect 69385 3587 69443 3593
rect 69385 3584 69397 3587
rect 68336 3556 69397 3584
rect 68336 3544 68342 3556
rect 69385 3553 69397 3556
rect 69431 3553 69443 3587
rect 71406 3584 71412 3596
rect 71367 3556 71412 3584
rect 69385 3547 69443 3553
rect 71406 3544 71412 3556
rect 71464 3544 71470 3596
rect 71590 3584 71596 3596
rect 71551 3556 71596 3584
rect 71590 3544 71596 3556
rect 71648 3544 71654 3596
rect 75362 3584 75368 3596
rect 75323 3556 75368 3584
rect 75362 3544 75368 3556
rect 75420 3544 75426 3596
rect 77110 3544 77116 3596
rect 77168 3584 77174 3596
rect 78508 3593 78536 3624
rect 77849 3587 77907 3593
rect 77849 3584 77861 3587
rect 77168 3556 77861 3584
rect 77168 3544 77174 3556
rect 77849 3553 77861 3556
rect 77895 3553 77907 3587
rect 77849 3547 77907 3553
rect 78493 3587 78551 3593
rect 78493 3553 78505 3587
rect 78539 3553 78551 3587
rect 78766 3584 78772 3596
rect 78727 3556 78772 3584
rect 78493 3547 78551 3553
rect 78766 3544 78772 3556
rect 78824 3544 78830 3596
rect 80146 3544 80152 3596
rect 80204 3584 80210 3596
rect 80241 3587 80299 3593
rect 80241 3584 80253 3587
rect 80204 3556 80253 3584
rect 80204 3544 80210 3556
rect 80241 3553 80253 3556
rect 80287 3584 80299 3587
rect 81342 3584 81348 3596
rect 80287 3556 81348 3584
rect 80287 3553 80299 3556
rect 80241 3547 80299 3553
rect 81342 3544 81348 3556
rect 81400 3544 81406 3596
rect 81897 3587 81955 3593
rect 81897 3553 81909 3587
rect 81943 3584 81955 3587
rect 81986 3584 81992 3596
rect 81943 3556 81992 3584
rect 81943 3553 81955 3556
rect 81897 3547 81955 3553
rect 81986 3544 81992 3556
rect 82044 3584 82050 3596
rect 83001 3587 83059 3593
rect 83001 3584 83013 3587
rect 82044 3556 83013 3584
rect 82044 3544 82050 3556
rect 83001 3553 83013 3556
rect 83047 3553 83059 3587
rect 83001 3547 83059 3553
rect 83274 3544 83280 3596
rect 83332 3584 83338 3596
rect 89686 3584 89714 3624
rect 93826 3624 104532 3652
rect 93826 3584 93854 3624
rect 104526 3612 104532 3624
rect 104584 3612 104590 3664
rect 83332 3556 83964 3584
rect 89686 3556 93854 3584
rect 83332 3544 83338 3556
rect 67361 3519 67419 3525
rect 67361 3485 67373 3519
rect 67407 3485 67419 3519
rect 67361 3479 67419 3485
rect 67634 3476 67640 3528
rect 67692 3516 67698 3528
rect 68373 3519 68431 3525
rect 68373 3516 68385 3519
rect 67692 3488 68385 3516
rect 67692 3476 67698 3488
rect 68373 3485 68385 3488
rect 68419 3485 68431 3519
rect 68373 3479 68431 3485
rect 68462 3476 68468 3528
rect 68520 3516 68526 3528
rect 68520 3488 68565 3516
rect 68520 3476 68526 3488
rect 69106 3476 69112 3528
rect 69164 3516 69170 3528
rect 69569 3519 69627 3525
rect 69569 3516 69581 3519
rect 69164 3488 69581 3516
rect 69164 3476 69170 3488
rect 69569 3485 69581 3488
rect 69615 3485 69627 3519
rect 69569 3479 69627 3485
rect 69658 3476 69664 3528
rect 69716 3516 69722 3528
rect 69716 3488 69761 3516
rect 69716 3476 69722 3488
rect 69934 3476 69940 3528
rect 69992 3476 69998 3528
rect 70026 3476 70032 3528
rect 70084 3516 70090 3528
rect 73525 3519 73583 3525
rect 73525 3516 73537 3519
rect 70084 3488 73537 3516
rect 70084 3476 70090 3488
rect 73525 3485 73537 3488
rect 73571 3516 73583 3519
rect 74074 3516 74080 3528
rect 73571 3488 74080 3516
rect 73571 3485 73583 3488
rect 73525 3479 73583 3485
rect 74074 3476 74080 3488
rect 74132 3476 74138 3528
rect 74169 3519 74227 3525
rect 74169 3485 74181 3519
rect 74215 3516 74227 3519
rect 74534 3516 74540 3528
rect 74215 3488 74540 3516
rect 74215 3485 74227 3488
rect 74169 3479 74227 3485
rect 74534 3476 74540 3488
rect 74592 3476 74598 3528
rect 75273 3519 75331 3525
rect 75273 3485 75285 3519
rect 75319 3516 75331 3519
rect 75730 3516 75736 3528
rect 75319 3488 75736 3516
rect 75319 3485 75331 3488
rect 75273 3479 75331 3485
rect 75730 3476 75736 3488
rect 75788 3476 75794 3528
rect 75822 3476 75828 3528
rect 75880 3516 75886 3528
rect 76101 3519 76159 3525
rect 76101 3516 76113 3519
rect 75880 3488 76113 3516
rect 75880 3476 75886 3488
rect 76101 3485 76113 3488
rect 76147 3516 76159 3519
rect 76558 3516 76564 3528
rect 76147 3488 76564 3516
rect 76147 3485 76159 3488
rect 76101 3479 76159 3485
rect 76558 3476 76564 3488
rect 76616 3476 76622 3528
rect 76837 3519 76895 3525
rect 76837 3485 76849 3519
rect 76883 3516 76895 3519
rect 77757 3519 77815 3525
rect 76883 3488 77340 3516
rect 76883 3485 76895 3488
rect 76837 3479 76895 3485
rect 69750 3448 69756 3460
rect 66640 3420 69756 3448
rect 69750 3408 69756 3420
rect 69808 3408 69814 3460
rect 69952 3448 69980 3476
rect 69860 3420 69980 3448
rect 66806 3380 66812 3392
rect 63604 3352 66812 3380
rect 66806 3340 66812 3352
rect 66864 3340 66870 3392
rect 67266 3380 67272 3392
rect 67227 3352 67272 3380
rect 67266 3340 67272 3352
rect 67324 3340 67330 3392
rect 67358 3340 67364 3392
rect 67416 3380 67422 3392
rect 69860 3380 69888 3420
rect 70118 3408 70124 3460
rect 70176 3448 70182 3460
rect 76190 3448 76196 3460
rect 70176 3420 76196 3448
rect 70176 3408 70182 3420
rect 76190 3408 76196 3420
rect 76248 3408 76254 3460
rect 67416 3352 69888 3380
rect 67416 3340 67422 3352
rect 69934 3340 69940 3392
rect 69992 3380 69998 3392
rect 70949 3383 71007 3389
rect 70949 3380 70961 3383
rect 69992 3352 70961 3380
rect 69992 3340 69998 3352
rect 70949 3349 70961 3352
rect 70995 3349 71007 3383
rect 70949 3343 71007 3349
rect 71317 3383 71375 3389
rect 71317 3349 71329 3383
rect 71363 3380 71375 3383
rect 72237 3383 72295 3389
rect 72237 3380 72249 3383
rect 71363 3352 72249 3380
rect 71363 3349 71375 3352
rect 71317 3343 71375 3349
rect 72237 3349 72249 3352
rect 72283 3380 72295 3383
rect 72694 3380 72700 3392
rect 72283 3352 72700 3380
rect 72283 3349 72295 3352
rect 72237 3343 72295 3349
rect 72694 3340 72700 3352
rect 72752 3340 72758 3392
rect 72878 3340 72884 3392
rect 72936 3380 72942 3392
rect 72973 3383 73031 3389
rect 72973 3380 72985 3383
rect 72936 3352 72985 3380
rect 72936 3340 72942 3352
rect 72973 3349 72985 3352
rect 73019 3349 73031 3383
rect 72973 3343 73031 3349
rect 74442 3340 74448 3392
rect 74500 3380 74506 3392
rect 74813 3383 74871 3389
rect 74813 3380 74825 3383
rect 74500 3352 74825 3380
rect 74500 3340 74506 3352
rect 74813 3349 74825 3352
rect 74859 3349 74871 3383
rect 74813 3343 74871 3349
rect 75181 3383 75239 3389
rect 75181 3349 75193 3383
rect 75227 3380 75239 3383
rect 75822 3380 75828 3392
rect 75227 3352 75828 3380
rect 75227 3349 75239 3352
rect 75181 3343 75239 3349
rect 75822 3340 75828 3352
rect 75880 3340 75886 3392
rect 76374 3340 76380 3392
rect 76432 3380 76438 3392
rect 77312 3389 77340 3488
rect 77757 3485 77769 3519
rect 77803 3516 77815 3519
rect 78214 3516 78220 3528
rect 77803 3488 78220 3516
rect 77803 3485 77815 3488
rect 77757 3479 77815 3485
rect 78214 3476 78220 3488
rect 78272 3476 78278 3528
rect 81621 3519 81679 3525
rect 81621 3485 81633 3519
rect 81667 3516 81679 3519
rect 82814 3516 82820 3528
rect 81667 3488 82820 3516
rect 81667 3485 81679 3488
rect 81621 3479 81679 3485
rect 82814 3476 82820 3488
rect 82872 3476 82878 3528
rect 82909 3519 82967 3525
rect 82909 3485 82921 3519
rect 82955 3516 82967 3519
rect 83826 3516 83832 3528
rect 82955 3488 83832 3516
rect 82955 3485 82967 3488
rect 82909 3479 82967 3485
rect 83826 3476 83832 3488
rect 83884 3476 83890 3528
rect 83936 3516 83964 3556
rect 83936 3488 89714 3516
rect 79410 3408 79416 3460
rect 79468 3408 79474 3460
rect 81713 3451 81771 3457
rect 81713 3417 81725 3451
rect 81759 3448 81771 3451
rect 81802 3448 81808 3460
rect 81759 3420 81808 3448
rect 81759 3417 81771 3420
rect 81713 3411 81771 3417
rect 81802 3408 81808 3420
rect 81860 3408 81866 3460
rect 82354 3408 82360 3460
rect 82412 3448 82418 3460
rect 84197 3451 84255 3457
rect 84197 3448 84209 3451
rect 82412 3420 84209 3448
rect 82412 3408 82418 3420
rect 84197 3417 84209 3420
rect 84243 3417 84255 3451
rect 89686 3448 89714 3488
rect 108298 3448 108304 3460
rect 89686 3420 108304 3448
rect 84197 3411 84255 3417
rect 108298 3408 108304 3420
rect 108356 3408 108362 3460
rect 76653 3383 76711 3389
rect 76653 3380 76665 3383
rect 76432 3352 76665 3380
rect 76432 3340 76438 3352
rect 76653 3349 76665 3352
rect 76699 3349 76711 3383
rect 76653 3343 76711 3349
rect 77297 3383 77355 3389
rect 77297 3349 77309 3383
rect 77343 3349 77355 3383
rect 77662 3380 77668 3392
rect 77575 3352 77668 3380
rect 77297 3343 77355 3349
rect 77662 3340 77668 3352
rect 77720 3380 77726 3392
rect 78122 3380 78128 3392
rect 77720 3352 78128 3380
rect 77720 3340 77726 3352
rect 78122 3340 78128 3352
rect 78180 3340 78186 3392
rect 81820 3380 81848 3408
rect 82722 3380 82728 3392
rect 81820 3352 82728 3380
rect 82722 3340 82728 3352
rect 82780 3340 82786 3392
rect 82817 3383 82875 3389
rect 82817 3349 82829 3383
rect 82863 3380 82875 3383
rect 83366 3380 83372 3392
rect 82863 3352 83372 3380
rect 82863 3349 82875 3352
rect 82817 3343 82875 3349
rect 83366 3340 83372 3352
rect 83424 3340 83430 3392
rect 83642 3380 83648 3392
rect 83603 3352 83648 3380
rect 83642 3340 83648 3352
rect 83700 3340 83706 3392
rect 85390 3380 85396 3392
rect 85351 3352 85396 3380
rect 85390 3340 85396 3352
rect 85448 3340 85454 3392
rect 1104 3290 148856 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 81014 3290
rect 81066 3238 81078 3290
rect 81130 3238 81142 3290
rect 81194 3238 81206 3290
rect 81258 3238 81270 3290
rect 81322 3238 111734 3290
rect 111786 3238 111798 3290
rect 111850 3238 111862 3290
rect 111914 3238 111926 3290
rect 111978 3238 111990 3290
rect 112042 3238 142454 3290
rect 142506 3238 142518 3290
rect 142570 3238 142582 3290
rect 142634 3238 142646 3290
rect 142698 3238 142710 3290
rect 142762 3238 148856 3290
rect 1104 3216 148856 3238
rect 5718 3176 5724 3188
rect 5679 3148 5724 3176
rect 5718 3136 5724 3148
rect 5776 3136 5782 3188
rect 5813 3179 5871 3185
rect 5813 3145 5825 3179
rect 5859 3176 5871 3179
rect 8113 3179 8171 3185
rect 8113 3176 8125 3179
rect 5859 3148 8125 3176
rect 5859 3145 5871 3148
rect 5813 3139 5871 3145
rect 8113 3145 8125 3148
rect 8159 3145 8171 3179
rect 9398 3176 9404 3188
rect 9359 3148 9404 3176
rect 8113 3139 8171 3145
rect 9398 3136 9404 3148
rect 9456 3136 9462 3188
rect 21634 3136 21640 3188
rect 21692 3176 21698 3188
rect 24210 3176 24216 3188
rect 21692 3148 23520 3176
rect 24171 3148 24216 3176
rect 21692 3136 21698 3148
rect 4614 3068 4620 3120
rect 4672 3108 4678 3120
rect 5261 3111 5319 3117
rect 5261 3108 5273 3111
rect 4672 3080 5273 3108
rect 4672 3068 4678 3080
rect 5261 3077 5273 3080
rect 5307 3077 5319 3111
rect 5994 3108 6000 3120
rect 5955 3080 6000 3108
rect 5261 3071 5319 3077
rect 5994 3068 6000 3080
rect 6052 3068 6058 3120
rect 6822 3068 6828 3120
rect 6880 3108 6886 3120
rect 23492 3117 23520 3148
rect 24210 3136 24216 3148
rect 24268 3136 24274 3188
rect 24670 3176 24676 3188
rect 24631 3148 24676 3176
rect 24670 3136 24676 3148
rect 24728 3136 24734 3188
rect 24946 3176 24952 3188
rect 24780 3148 24952 3176
rect 21361 3111 21419 3117
rect 6880 3080 9260 3108
rect 6880 3068 6886 3080
rect 6730 3040 6736 3052
rect 6691 3012 6736 3040
rect 6730 3000 6736 3012
rect 6788 3000 6794 3052
rect 7006 3040 7012 3052
rect 6967 3012 7012 3040
rect 7006 3000 7012 3012
rect 7064 3000 7070 3052
rect 8018 3000 8024 3052
rect 8076 3040 8082 3052
rect 9232 3049 9260 3080
rect 21361 3077 21373 3111
rect 21407 3108 21419 3111
rect 23477 3111 23535 3117
rect 21407 3080 22310 3108
rect 21407 3077 21419 3080
rect 21361 3071 21419 3077
rect 23477 3077 23489 3111
rect 23523 3077 23535 3111
rect 23477 3071 23535 3077
rect 8297 3043 8355 3049
rect 8297 3040 8309 3043
rect 8076 3012 8309 3040
rect 8076 3000 8082 3012
rect 8297 3009 8309 3012
rect 8343 3009 8355 3043
rect 8297 3003 8355 3009
rect 9217 3043 9275 3049
rect 9217 3009 9229 3043
rect 9263 3009 9275 3043
rect 9398 3040 9404 3052
rect 9359 3012 9404 3040
rect 9217 3003 9275 3009
rect 9398 3000 9404 3012
rect 9456 3000 9462 3052
rect 20809 3043 20867 3049
rect 20809 3009 20821 3043
rect 20855 3040 20867 3043
rect 20990 3040 20996 3052
rect 20855 3012 20996 3040
rect 20855 3009 20867 3012
rect 20809 3003 20867 3009
rect 20990 3000 20996 3012
rect 21048 3040 21054 3052
rect 21269 3043 21327 3049
rect 21269 3040 21281 3043
rect 21048 3012 21281 3040
rect 21048 3000 21054 3012
rect 21269 3009 21281 3012
rect 21315 3040 21327 3043
rect 22094 3040 22100 3052
rect 21315 3012 22100 3040
rect 21315 3009 21327 3012
rect 21269 3003 21327 3009
rect 22094 3000 22100 3012
rect 22152 3000 22158 3052
rect 23750 3000 23756 3052
rect 23808 3040 23814 3052
rect 24581 3043 24639 3049
rect 23808 3012 23853 3040
rect 23808 3000 23814 3012
rect 24581 3009 24593 3043
rect 24627 3009 24639 3043
rect 24581 3003 24639 3009
rect 3878 2932 3884 2984
rect 3936 2972 3942 2984
rect 20257 2975 20315 2981
rect 3936 2944 5396 2972
rect 3936 2932 3942 2944
rect 5261 2907 5319 2913
rect 5261 2873 5273 2907
rect 5307 2873 5319 2907
rect 5368 2904 5396 2944
rect 20257 2941 20269 2975
rect 20303 2972 20315 2975
rect 21450 2972 21456 2984
rect 20303 2944 21456 2972
rect 20303 2941 20315 2944
rect 20257 2935 20315 2941
rect 21450 2932 21456 2944
rect 21508 2932 21514 2984
rect 21910 2932 21916 2984
rect 21968 2972 21974 2984
rect 22005 2975 22063 2981
rect 22005 2972 22017 2975
rect 21968 2944 22017 2972
rect 21968 2932 21974 2944
rect 22005 2941 22017 2944
rect 22051 2972 22063 2975
rect 24596 2972 24624 3003
rect 24780 2981 24808 3148
rect 24946 3136 24952 3148
rect 25004 3176 25010 3188
rect 27338 3176 27344 3188
rect 25004 3148 26372 3176
rect 27299 3148 27344 3176
rect 25004 3136 25010 3148
rect 26344 3108 26372 3148
rect 27338 3136 27344 3148
rect 27396 3136 27402 3188
rect 27709 3179 27767 3185
rect 27709 3145 27721 3179
rect 27755 3176 27767 3179
rect 27982 3176 27988 3188
rect 27755 3148 27988 3176
rect 27755 3145 27767 3148
rect 27709 3139 27767 3145
rect 27982 3136 27988 3148
rect 28040 3136 28046 3188
rect 28537 3179 28595 3185
rect 28537 3145 28549 3179
rect 28583 3145 28595 3179
rect 28537 3139 28595 3145
rect 27522 3108 27528 3120
rect 26344 3080 27528 3108
rect 27522 3068 27528 3080
rect 27580 3068 27586 3120
rect 27801 3111 27859 3117
rect 27801 3077 27813 3111
rect 27847 3108 27859 3111
rect 28350 3108 28356 3120
rect 27847 3080 28356 3108
rect 27847 3077 27859 3080
rect 27801 3071 27859 3077
rect 28350 3068 28356 3080
rect 28408 3068 28414 3120
rect 25777 3043 25835 3049
rect 25777 3009 25789 3043
rect 25823 3009 25835 3043
rect 25777 3003 25835 3009
rect 22051 2944 24624 2972
rect 24765 2975 24823 2981
rect 22051 2941 22063 2944
rect 22005 2935 22063 2941
rect 24765 2941 24777 2975
rect 24811 2941 24823 2975
rect 25792 2972 25820 3003
rect 25866 3000 25872 3052
rect 25924 3040 25930 3052
rect 26326 3040 26332 3052
rect 25924 3012 26332 3040
rect 25924 3000 25930 3012
rect 26326 3000 26332 3012
rect 26384 3040 26390 3052
rect 26421 3043 26479 3049
rect 26421 3040 26433 3043
rect 26384 3012 26433 3040
rect 26384 3000 26390 3012
rect 26421 3009 26433 3012
rect 26467 3009 26479 3043
rect 28552 3040 28580 3139
rect 28810 3136 28816 3188
rect 28868 3176 28874 3188
rect 28997 3179 29055 3185
rect 28997 3176 29009 3179
rect 28868 3148 29009 3176
rect 28868 3136 28874 3148
rect 28997 3145 29009 3148
rect 29043 3145 29055 3179
rect 30834 3176 30840 3188
rect 30795 3148 30840 3176
rect 28997 3139 29055 3145
rect 30834 3136 30840 3148
rect 30892 3136 30898 3188
rect 33778 3176 33784 3188
rect 30944 3148 31800 3176
rect 33739 3148 33784 3176
rect 28626 3068 28632 3120
rect 28684 3108 28690 3120
rect 28902 3108 28908 3120
rect 28684 3080 28908 3108
rect 28684 3068 28690 3080
rect 28902 3068 28908 3080
rect 28960 3068 28966 3120
rect 29822 3108 29828 3120
rect 29783 3080 29828 3108
rect 29822 3068 29828 3080
rect 29880 3068 29886 3120
rect 30098 3068 30104 3120
rect 30156 3108 30162 3120
rect 30282 3108 30288 3120
rect 30156 3080 30288 3108
rect 30156 3068 30162 3080
rect 30282 3068 30288 3080
rect 30340 3108 30346 3120
rect 30745 3111 30803 3117
rect 30745 3108 30757 3111
rect 30340 3080 30757 3108
rect 30340 3068 30346 3080
rect 30745 3077 30757 3080
rect 30791 3077 30803 3111
rect 30745 3071 30803 3077
rect 30944 3040 30972 3148
rect 31478 3108 31484 3120
rect 31439 3080 31484 3108
rect 31478 3068 31484 3080
rect 31536 3068 31542 3120
rect 31662 3108 31668 3120
rect 31623 3080 31668 3108
rect 31662 3068 31668 3080
rect 31720 3068 31726 3120
rect 26421 3003 26479 3009
rect 26528 3012 28580 3040
rect 30116 3012 30972 3040
rect 26528 2972 26556 3012
rect 25792 2944 26556 2972
rect 24765 2935 24823 2941
rect 27614 2932 27620 2984
rect 27672 2972 27678 2984
rect 30116 2981 30144 3012
rect 27893 2975 27951 2981
rect 27893 2972 27905 2975
rect 27672 2944 27905 2972
rect 27672 2932 27678 2944
rect 27893 2941 27905 2944
rect 27939 2972 27951 2975
rect 29089 2975 29147 2981
rect 29089 2972 29101 2975
rect 27939 2944 29101 2972
rect 27939 2941 27951 2944
rect 27893 2935 27951 2941
rect 29089 2941 29101 2944
rect 29135 2972 29147 2975
rect 30101 2975 30159 2981
rect 30101 2972 30113 2975
rect 29135 2944 30113 2972
rect 29135 2941 29147 2944
rect 29089 2935 29147 2941
rect 30101 2941 30113 2944
rect 30147 2941 30159 2975
rect 31772 2972 31800 3148
rect 33778 3136 33784 3148
rect 33836 3136 33842 3188
rect 34146 3176 34152 3188
rect 34107 3148 34152 3176
rect 34146 3136 34152 3148
rect 34204 3136 34210 3188
rect 34241 3179 34299 3185
rect 34241 3145 34253 3179
rect 34287 3176 34299 3179
rect 34422 3176 34428 3188
rect 34287 3148 34428 3176
rect 34287 3145 34299 3148
rect 34241 3139 34299 3145
rect 32401 3111 32459 3117
rect 32401 3077 32413 3111
rect 32447 3108 32459 3111
rect 34256 3108 34284 3139
rect 34422 3136 34428 3148
rect 34480 3136 34486 3188
rect 37458 3176 37464 3188
rect 37419 3148 37464 3176
rect 37458 3136 37464 3148
rect 37516 3136 37522 3188
rect 37921 3179 37979 3185
rect 37921 3145 37933 3179
rect 37967 3176 37979 3179
rect 38102 3176 38108 3188
rect 37967 3148 38108 3176
rect 37967 3145 37979 3148
rect 37921 3139 37979 3145
rect 38102 3136 38108 3148
rect 38160 3136 38166 3188
rect 45005 3179 45063 3185
rect 45005 3176 45017 3179
rect 38212 3148 45017 3176
rect 38212 3120 38240 3148
rect 45005 3145 45017 3148
rect 45051 3176 45063 3179
rect 46842 3176 46848 3188
rect 45051 3148 46848 3176
rect 45051 3145 45063 3148
rect 45005 3139 45063 3145
rect 46842 3136 46848 3148
rect 46900 3176 46906 3188
rect 54018 3176 54024 3188
rect 46900 3148 47808 3176
rect 46900 3136 46906 3148
rect 32447 3080 34284 3108
rect 36909 3111 36967 3117
rect 32447 3077 32459 3080
rect 32401 3071 32459 3077
rect 36909 3077 36921 3111
rect 36955 3108 36967 3111
rect 38194 3108 38200 3120
rect 36955 3080 38200 3108
rect 36955 3077 36967 3080
rect 36909 3071 36967 3077
rect 38194 3068 38200 3080
rect 38252 3068 38258 3120
rect 39206 3108 39212 3120
rect 39167 3080 39212 3108
rect 39206 3068 39212 3080
rect 39264 3068 39270 3120
rect 39942 3068 39948 3120
rect 40000 3068 40006 3120
rect 41506 3068 41512 3120
rect 41564 3108 41570 3120
rect 41601 3111 41659 3117
rect 41601 3108 41613 3111
rect 41564 3080 41613 3108
rect 41564 3068 41570 3080
rect 41601 3077 41613 3080
rect 41647 3077 41659 3111
rect 41601 3071 41659 3077
rect 41693 3111 41751 3117
rect 41693 3077 41705 3111
rect 41739 3108 41751 3111
rect 43346 3108 43352 3120
rect 41739 3080 43352 3108
rect 41739 3077 41751 3080
rect 41693 3071 41751 3077
rect 43346 3068 43352 3080
rect 43404 3068 43410 3120
rect 45925 3111 45983 3117
rect 45925 3077 45937 3111
rect 45971 3108 45983 3111
rect 46014 3108 46020 3120
rect 45971 3080 46020 3108
rect 45971 3077 45983 3080
rect 45925 3071 45983 3077
rect 46014 3068 46020 3080
rect 46072 3068 46078 3120
rect 47780 3117 47808 3148
rect 49528 3148 54024 3176
rect 49528 3117 49556 3148
rect 54018 3136 54024 3148
rect 54076 3176 54082 3188
rect 57330 3176 57336 3188
rect 54076 3148 54340 3176
rect 57291 3148 57336 3176
rect 54076 3136 54082 3148
rect 47765 3111 47823 3117
rect 47765 3077 47777 3111
rect 47811 3077 47823 3111
rect 47765 3071 47823 3077
rect 49513 3111 49571 3117
rect 49513 3077 49525 3111
rect 49559 3077 49571 3111
rect 50890 3108 50896 3120
rect 50851 3080 50896 3108
rect 49513 3071 49571 3077
rect 50890 3068 50896 3080
rect 50948 3068 50954 3120
rect 51626 3068 51632 3120
rect 51684 3068 51690 3120
rect 53282 3108 53288 3120
rect 53243 3080 53288 3108
rect 53282 3068 53288 3080
rect 53340 3068 53346 3120
rect 53377 3111 53435 3117
rect 53377 3077 53389 3111
rect 53423 3108 53435 3111
rect 53834 3108 53840 3120
rect 53423 3080 53840 3108
rect 53423 3077 53435 3080
rect 53377 3071 53435 3077
rect 53834 3068 53840 3080
rect 53892 3068 53898 3120
rect 32766 3000 32772 3052
rect 32824 3040 32830 3052
rect 32861 3043 32919 3049
rect 32861 3040 32873 3043
rect 32824 3012 32873 3040
rect 32824 3000 32830 3012
rect 32861 3009 32873 3012
rect 32907 3009 32919 3043
rect 37829 3043 37887 3049
rect 32861 3003 32919 3009
rect 32968 3012 35894 3040
rect 32968 2972 32996 3012
rect 31772 2944 32996 2972
rect 33137 2975 33195 2981
rect 30101 2935 30159 2941
rect 33137 2941 33149 2975
rect 33183 2972 33195 2975
rect 33686 2972 33692 2984
rect 33183 2944 33692 2972
rect 33183 2941 33195 2944
rect 33137 2935 33195 2941
rect 33686 2932 33692 2944
rect 33744 2932 33750 2984
rect 34440 2981 34468 3012
rect 34425 2975 34483 2981
rect 34425 2941 34437 2975
rect 34471 2941 34483 2975
rect 34425 2935 34483 2941
rect 34790 2932 34796 2984
rect 34848 2972 34854 2984
rect 35161 2975 35219 2981
rect 35161 2972 35173 2975
rect 34848 2944 35173 2972
rect 34848 2932 34854 2944
rect 35161 2941 35173 2944
rect 35207 2941 35219 2975
rect 35866 2972 35894 3012
rect 37829 3009 37841 3043
rect 37875 3040 37887 3043
rect 37875 3012 38516 3040
rect 37875 3009 37887 3012
rect 37829 3003 37887 3009
rect 35986 2972 35992 2984
rect 35866 2944 35992 2972
rect 35161 2935 35219 2941
rect 35986 2932 35992 2944
rect 36044 2972 36050 2984
rect 36906 2972 36912 2984
rect 36044 2944 36912 2972
rect 36044 2932 36050 2944
rect 36906 2932 36912 2944
rect 36964 2972 36970 2984
rect 38013 2975 38071 2981
rect 38013 2972 38025 2975
rect 36964 2944 38025 2972
rect 36964 2932 36970 2944
rect 38013 2941 38025 2944
rect 38059 2941 38071 2975
rect 38488 2972 38516 3012
rect 38562 3000 38568 3052
rect 38620 3040 38626 3052
rect 38933 3043 38991 3049
rect 38933 3040 38945 3043
rect 38620 3012 38945 3040
rect 38620 3000 38626 3012
rect 38933 3009 38945 3012
rect 38979 3009 38991 3043
rect 42518 3040 42524 3052
rect 38933 3003 38991 3009
rect 41432 3012 42524 3040
rect 41432 2984 41460 3012
rect 42518 3000 42524 3012
rect 42576 3000 42582 3052
rect 42610 3000 42616 3052
rect 42668 3040 42674 3052
rect 42705 3043 42763 3049
rect 42705 3040 42717 3043
rect 42668 3012 42717 3040
rect 42668 3000 42674 3012
rect 42705 3009 42717 3012
rect 42751 3040 42763 3043
rect 43717 3043 43775 3049
rect 43717 3040 43729 3043
rect 42751 3012 43729 3040
rect 42751 3009 42763 3012
rect 42705 3003 42763 3009
rect 43717 3009 43729 3012
rect 43763 3009 43775 3043
rect 43717 3003 43775 3009
rect 45462 3000 45468 3052
rect 45520 3040 45526 3052
rect 46109 3043 46167 3049
rect 46109 3040 46121 3043
rect 45520 3012 46121 3040
rect 45520 3000 45526 3012
rect 46109 3009 46121 3012
rect 46155 3009 46167 3043
rect 46109 3003 46167 3009
rect 46753 3043 46811 3049
rect 46753 3009 46765 3043
rect 46799 3009 46811 3043
rect 46753 3003 46811 3009
rect 39206 2972 39212 2984
rect 38488 2944 39212 2972
rect 38013 2935 38071 2941
rect 39206 2932 39212 2944
rect 39264 2932 39270 2984
rect 41414 2932 41420 2984
rect 41472 2972 41478 2984
rect 46768 2972 46796 3003
rect 49326 3000 49332 3052
rect 49384 3040 49390 3052
rect 50157 3043 50215 3049
rect 50157 3040 50169 3043
rect 49384 3012 50169 3040
rect 49384 3000 49390 3012
rect 50157 3009 50169 3012
rect 50203 3009 50215 3043
rect 50614 3040 50620 3052
rect 50575 3012 50620 3040
rect 50157 3003 50215 3009
rect 50614 3000 50620 3012
rect 50672 3000 50678 3052
rect 54312 3049 54340 3148
rect 57330 3136 57336 3148
rect 57388 3136 57394 3188
rect 58710 3136 58716 3188
rect 58768 3176 58774 3188
rect 65150 3176 65156 3188
rect 58768 3148 65156 3176
rect 58768 3136 58774 3148
rect 54570 3108 54576 3120
rect 54531 3080 54576 3108
rect 54570 3068 54576 3080
rect 54628 3068 54634 3120
rect 55214 3068 55220 3120
rect 55272 3068 55278 3120
rect 57425 3111 57483 3117
rect 57425 3077 57437 3111
rect 57471 3108 57483 3111
rect 57698 3108 57704 3120
rect 57471 3080 57704 3108
rect 57471 3077 57483 3080
rect 57425 3071 57483 3077
rect 57698 3068 57704 3080
rect 57756 3108 57762 3120
rect 58066 3108 58072 3120
rect 57756 3080 58072 3108
rect 57756 3068 57762 3080
rect 58066 3068 58072 3080
rect 58124 3068 58130 3120
rect 58529 3111 58587 3117
rect 58529 3077 58541 3111
rect 58575 3108 58587 3111
rect 58986 3108 58992 3120
rect 58575 3080 58992 3108
rect 58575 3077 58587 3080
rect 58529 3071 58587 3077
rect 58986 3068 58992 3080
rect 59044 3068 59050 3120
rect 54297 3043 54355 3049
rect 54297 3009 54309 3043
rect 54343 3009 54355 3043
rect 54297 3003 54355 3009
rect 41472 2944 41517 2972
rect 41984 2944 46796 2972
rect 52365 2975 52423 2981
rect 41472 2932 41478 2944
rect 41690 2904 41696 2916
rect 5368 2876 22094 2904
rect 5261 2867 5319 2873
rect 4709 2839 4767 2845
rect 4709 2805 4721 2839
rect 4755 2836 4767 2839
rect 5276 2836 5304 2867
rect 5350 2836 5356 2848
rect 4755 2808 5356 2836
rect 4755 2805 4767 2808
rect 4709 2799 4767 2805
rect 5350 2796 5356 2808
rect 5408 2796 5414 2848
rect 14918 2796 14924 2848
rect 14976 2836 14982 2848
rect 15013 2839 15071 2845
rect 15013 2836 15025 2839
rect 14976 2808 15025 2836
rect 14976 2796 14982 2808
rect 15013 2805 15025 2808
rect 15059 2805 15071 2839
rect 15013 2799 15071 2805
rect 20622 2796 20628 2848
rect 20680 2836 20686 2848
rect 21818 2836 21824 2848
rect 20680 2808 21824 2836
rect 20680 2796 20686 2808
rect 21818 2796 21824 2808
rect 21876 2796 21882 2848
rect 22066 2836 22094 2876
rect 23676 2876 35894 2904
rect 23676 2836 23704 2876
rect 22066 2808 23704 2836
rect 25961 2839 26019 2845
rect 25961 2805 25973 2839
rect 26007 2836 26019 2839
rect 26326 2836 26332 2848
rect 26007 2808 26332 2836
rect 26007 2805 26019 2808
rect 25961 2799 26019 2805
rect 26326 2796 26332 2808
rect 26384 2796 26390 2848
rect 26513 2839 26571 2845
rect 26513 2805 26525 2839
rect 26559 2836 26571 2839
rect 27890 2836 27896 2848
rect 26559 2808 27896 2836
rect 26559 2805 26571 2808
rect 26513 2799 26571 2805
rect 27890 2796 27896 2808
rect 27948 2796 27954 2848
rect 35866 2836 35894 2876
rect 40604 2876 41696 2904
rect 40604 2836 40632 2876
rect 41690 2864 41696 2876
rect 41748 2864 41754 2916
rect 35866 2808 40632 2836
rect 40678 2796 40684 2848
rect 40736 2836 40742 2848
rect 41984 2836 42012 2944
rect 52365 2941 52377 2975
rect 52411 2972 52423 2975
rect 52454 2972 52460 2984
rect 52411 2944 52460 2972
rect 52411 2941 52423 2944
rect 52365 2935 52423 2941
rect 52454 2932 52460 2944
rect 52512 2932 52518 2984
rect 53561 2975 53619 2981
rect 53561 2941 53573 2975
rect 53607 2972 53619 2975
rect 54202 2972 54208 2984
rect 53607 2944 54208 2972
rect 53607 2941 53619 2944
rect 53561 2935 53619 2941
rect 54202 2932 54208 2944
rect 54260 2932 54266 2984
rect 52178 2864 52184 2916
rect 52236 2904 52242 2916
rect 52917 2907 52975 2913
rect 52917 2904 52929 2907
rect 52236 2876 52929 2904
rect 52236 2864 52242 2876
rect 52917 2873 52929 2876
rect 52963 2873 52975 2907
rect 52917 2867 52975 2873
rect 40736 2808 42012 2836
rect 42061 2839 42119 2845
rect 40736 2796 40742 2808
rect 42061 2805 42073 2839
rect 42107 2836 42119 2839
rect 42150 2836 42156 2848
rect 42107 2808 42156 2836
rect 42107 2805 42119 2808
rect 42061 2799 42119 2805
rect 42150 2796 42156 2808
rect 42208 2796 42214 2848
rect 42518 2796 42524 2848
rect 42576 2836 42582 2848
rect 43165 2839 43223 2845
rect 43165 2836 43177 2839
rect 42576 2808 43177 2836
rect 42576 2796 42582 2808
rect 43165 2805 43177 2808
rect 43211 2805 43223 2839
rect 43165 2799 43223 2805
rect 46658 2796 46664 2848
rect 46716 2836 46722 2848
rect 46937 2839 46995 2845
rect 46937 2836 46949 2839
rect 46716 2808 46949 2836
rect 46716 2796 46722 2808
rect 46937 2805 46949 2808
rect 46983 2805 46995 2839
rect 50062 2836 50068 2848
rect 50023 2808 50068 2836
rect 46937 2799 46995 2805
rect 50062 2796 50068 2808
rect 50120 2796 50126 2848
rect 54312 2836 54340 3003
rect 56502 3000 56508 3052
rect 56560 3040 56566 3052
rect 56597 3043 56655 3049
rect 56597 3040 56609 3043
rect 56560 3012 56609 3040
rect 56560 3000 56566 3012
rect 56597 3009 56609 3012
rect 56643 3009 56655 3043
rect 56597 3003 56655 3009
rect 58437 3043 58495 3049
rect 58437 3009 58449 3043
rect 58483 3040 58495 3043
rect 59630 3040 59636 3052
rect 58483 3012 59636 3040
rect 58483 3009 58495 3012
rect 58437 3003 58495 3009
rect 59630 3000 59636 3012
rect 59688 3000 59694 3052
rect 59740 3049 59768 3148
rect 65150 3136 65156 3148
rect 65208 3176 65214 3188
rect 65208 3148 65288 3176
rect 65208 3136 65214 3148
rect 59998 3108 60004 3120
rect 59959 3080 60004 3108
rect 59998 3068 60004 3080
rect 60056 3068 60062 3120
rect 61378 3108 61384 3120
rect 61226 3080 61384 3108
rect 61378 3068 61384 3080
rect 61436 3068 61442 3120
rect 62114 3068 62120 3120
rect 62172 3108 62178 3120
rect 62209 3111 62267 3117
rect 62209 3108 62221 3111
rect 62172 3080 62221 3108
rect 62172 3068 62178 3080
rect 62209 3077 62221 3080
rect 62255 3077 62267 3111
rect 62209 3071 62267 3077
rect 63681 3111 63739 3117
rect 63681 3077 63693 3111
rect 63727 3108 63739 3111
rect 64046 3108 64052 3120
rect 63727 3080 64052 3108
rect 63727 3077 63739 3080
rect 63681 3071 63739 3077
rect 64046 3068 64052 3080
rect 64104 3068 64110 3120
rect 64322 3068 64328 3120
rect 64380 3108 64386 3120
rect 64598 3108 64604 3120
rect 64380 3080 64604 3108
rect 64380 3068 64386 3080
rect 64598 3068 64604 3080
rect 64656 3068 64662 3120
rect 64782 3108 64788 3120
rect 64743 3080 64788 3108
rect 64782 3068 64788 3080
rect 64840 3068 64846 3120
rect 59725 3043 59783 3049
rect 59725 3009 59737 3043
rect 59771 3009 59783 3043
rect 59725 3003 59783 3009
rect 61838 3000 61844 3052
rect 61896 3040 61902 3052
rect 61933 3043 61991 3049
rect 61933 3040 61945 3043
rect 61896 3012 61945 3040
rect 61896 3000 61902 3012
rect 61933 3009 61945 3012
rect 61979 3009 61991 3043
rect 63586 3040 63592 3052
rect 63499 3012 63592 3040
rect 61933 3003 61991 3009
rect 63586 3000 63592 3012
rect 63644 3040 63650 3052
rect 65260 3049 65288 3148
rect 66162 3136 66168 3188
rect 66220 3176 66226 3188
rect 68925 3179 68983 3185
rect 66220 3148 68876 3176
rect 66220 3136 66226 3148
rect 65518 3108 65524 3120
rect 65479 3080 65524 3108
rect 65518 3068 65524 3080
rect 65576 3068 65582 3120
rect 67266 3108 67272 3120
rect 66746 3080 67272 3108
rect 67266 3068 67272 3080
rect 67324 3068 67330 3120
rect 68848 3108 68876 3148
rect 68925 3145 68937 3179
rect 68971 3176 68983 3179
rect 69290 3176 69296 3188
rect 68971 3148 69296 3176
rect 68971 3145 68983 3148
rect 68925 3139 68983 3145
rect 69290 3136 69296 3148
rect 69348 3136 69354 3188
rect 69658 3136 69664 3188
rect 69716 3176 69722 3188
rect 71869 3179 71927 3185
rect 71869 3176 71881 3179
rect 69716 3148 71881 3176
rect 69716 3136 69722 3148
rect 71869 3145 71881 3148
rect 71915 3176 71927 3179
rect 72510 3176 72516 3188
rect 71915 3148 72516 3176
rect 71915 3145 71927 3148
rect 71869 3139 71927 3145
rect 72510 3136 72516 3148
rect 72568 3136 72574 3188
rect 73706 3176 73712 3188
rect 73667 3148 73712 3176
rect 73706 3136 73712 3148
rect 73764 3136 73770 3188
rect 77202 3176 77208 3188
rect 77163 3148 77208 3176
rect 77202 3136 77208 3148
rect 77260 3136 77266 3188
rect 78033 3179 78091 3185
rect 78033 3145 78045 3179
rect 78079 3176 78091 3179
rect 79778 3176 79784 3188
rect 78079 3148 79784 3176
rect 78079 3145 78091 3148
rect 78033 3139 78091 3145
rect 79778 3136 79784 3148
rect 79836 3136 79842 3188
rect 81710 3176 81716 3188
rect 81671 3148 81716 3176
rect 81710 3136 81716 3148
rect 81768 3136 81774 3188
rect 82173 3179 82231 3185
rect 82173 3145 82185 3179
rect 82219 3176 82231 3179
rect 82354 3176 82360 3188
rect 82219 3148 82360 3176
rect 82219 3145 82231 3148
rect 82173 3139 82231 3145
rect 82354 3136 82360 3148
rect 82412 3136 82418 3188
rect 83001 3179 83059 3185
rect 83001 3145 83013 3179
rect 83047 3176 83059 3179
rect 83182 3176 83188 3188
rect 83047 3148 83188 3176
rect 83047 3145 83059 3148
rect 83001 3139 83059 3145
rect 83182 3136 83188 3148
rect 83240 3136 83246 3188
rect 83366 3136 83372 3188
rect 83424 3176 83430 3188
rect 84102 3176 84108 3188
rect 83424 3148 84108 3176
rect 83424 3136 83430 3148
rect 84102 3136 84108 3148
rect 84160 3176 84166 3188
rect 125502 3176 125508 3188
rect 84160 3148 125508 3176
rect 84160 3136 84166 3148
rect 125502 3136 125508 3148
rect 125560 3136 125566 3188
rect 145926 3176 145932 3188
rect 145887 3148 145932 3176
rect 145926 3136 145932 3148
rect 145984 3136 145990 3188
rect 69842 3108 69848 3120
rect 68848 3080 69848 3108
rect 69842 3068 69848 3080
rect 69900 3068 69906 3120
rect 70394 3108 70400 3120
rect 70355 3080 70400 3108
rect 70394 3068 70400 3080
rect 70452 3068 70458 3120
rect 70486 3068 70492 3120
rect 70544 3108 70550 3120
rect 78677 3111 78735 3117
rect 78677 3108 78689 3111
rect 70544 3080 70886 3108
rect 77312 3080 78689 3108
rect 70544 3068 70550 3080
rect 65245 3043 65303 3049
rect 63644 3012 65012 3040
rect 63644 3000 63650 3012
rect 58618 2972 58624 2984
rect 58579 2944 58624 2972
rect 58618 2932 58624 2944
rect 58676 2932 58682 2984
rect 61470 2972 61476 2984
rect 61431 2944 61476 2972
rect 61470 2932 61476 2944
rect 61528 2932 61534 2984
rect 63862 2972 63868 2984
rect 63823 2944 63868 2972
rect 63862 2932 63868 2944
rect 63920 2932 63926 2984
rect 58069 2907 58127 2913
rect 58069 2873 58081 2907
rect 58115 2904 58127 2907
rect 58158 2904 58164 2916
rect 58115 2876 58164 2904
rect 58115 2873 58127 2876
rect 58069 2867 58127 2873
rect 58158 2864 58164 2876
rect 58216 2864 58222 2916
rect 62022 2864 62028 2916
rect 62080 2904 62086 2916
rect 63221 2907 63279 2913
rect 63221 2904 63233 2907
rect 62080 2876 63233 2904
rect 62080 2864 62086 2876
rect 63221 2873 63233 2876
rect 63267 2873 63279 2907
rect 63221 2867 63279 2873
rect 55674 2836 55680 2848
rect 54312 2808 55680 2836
rect 55674 2796 55680 2808
rect 55732 2796 55738 2848
rect 56042 2836 56048 2848
rect 56003 2808 56048 2836
rect 56042 2796 56048 2808
rect 56100 2796 56106 2848
rect 56686 2836 56692 2848
rect 56647 2808 56692 2836
rect 56686 2796 56692 2808
rect 56744 2796 56750 2848
rect 64984 2836 65012 3012
rect 65245 3009 65257 3043
rect 65291 3009 65303 3043
rect 65245 3003 65303 3009
rect 66806 3000 66812 3052
rect 66864 3040 66870 3052
rect 67545 3043 67603 3049
rect 67545 3040 67557 3043
rect 66864 3012 67557 3040
rect 66864 3000 66870 3012
rect 67545 3009 67557 3012
rect 67591 3009 67603 3043
rect 67545 3003 67603 3009
rect 68002 3000 68008 3052
rect 68060 3040 68066 3052
rect 68830 3040 68836 3052
rect 68060 3012 68836 3040
rect 68060 3000 68066 3012
rect 68830 3000 68836 3012
rect 68888 3000 68894 3052
rect 69477 3043 69535 3049
rect 69477 3009 69489 3043
rect 69523 3040 69535 3043
rect 69750 3040 69756 3052
rect 69523 3012 69756 3040
rect 69523 3009 69535 3012
rect 69477 3003 69535 3009
rect 69750 3000 69756 3012
rect 69808 3000 69814 3052
rect 70121 3043 70179 3049
rect 70121 3009 70133 3043
rect 70167 3009 70179 3043
rect 72418 3040 72424 3052
rect 72379 3012 72424 3040
rect 70121 3003 70179 3009
rect 65058 2932 65064 2984
rect 65116 2972 65122 2984
rect 69934 2972 69940 2984
rect 65116 2944 69940 2972
rect 65116 2932 65122 2944
rect 69934 2932 69940 2944
rect 69992 2932 69998 2984
rect 70136 2916 70164 3003
rect 72418 3000 72424 3012
rect 72476 3000 72482 3052
rect 72878 3000 72884 3052
rect 72936 3040 72942 3052
rect 73617 3043 73675 3049
rect 73617 3040 73629 3043
rect 72936 3012 73629 3040
rect 72936 3000 72942 3012
rect 73617 3009 73629 3012
rect 73663 3009 73675 3043
rect 74442 3040 74448 3052
rect 74403 3012 74448 3040
rect 73617 3003 73675 3009
rect 74442 3000 74448 3012
rect 74500 3000 74506 3052
rect 75086 3040 75092 3052
rect 75047 3012 75092 3040
rect 75086 3000 75092 3012
rect 75144 3000 75150 3052
rect 75730 3040 75736 3052
rect 75691 3012 75736 3040
rect 75730 3000 75736 3012
rect 75788 3000 75794 3052
rect 77018 3000 77024 3052
rect 77076 3040 77082 3052
rect 77312 3049 77340 3080
rect 78677 3077 78689 3080
rect 78723 3077 78735 3111
rect 82814 3108 82820 3120
rect 80730 3080 82820 3108
rect 78677 3071 78735 3077
rect 82814 3068 82820 3080
rect 82872 3068 82878 3120
rect 84565 3111 84623 3117
rect 84565 3108 84577 3111
rect 82924 3080 84577 3108
rect 77297 3043 77355 3049
rect 77297 3040 77309 3043
rect 77076 3012 77309 3040
rect 77076 3000 77082 3012
rect 77297 3009 77309 3012
rect 77343 3009 77355 3043
rect 77297 3003 77355 3009
rect 77849 3043 77907 3049
rect 77849 3009 77861 3043
rect 77895 3009 77907 3043
rect 77849 3003 77907 3009
rect 81253 3043 81311 3049
rect 81253 3009 81265 3043
rect 81299 3040 81311 3043
rect 82081 3043 82139 3049
rect 82081 3040 82093 3043
rect 81299 3012 82093 3040
rect 81299 3009 81311 3012
rect 81253 3003 81311 3009
rect 82081 3009 82093 3012
rect 82127 3040 82139 3043
rect 82924 3040 82952 3080
rect 84565 3077 84577 3080
rect 84611 3108 84623 3111
rect 137278 3108 137284 3120
rect 84611 3080 137284 3108
rect 84611 3077 84623 3080
rect 84565 3071 84623 3077
rect 137278 3068 137284 3080
rect 137336 3068 137342 3120
rect 82127 3012 82952 3040
rect 83093 3043 83151 3049
rect 82127 3009 82139 3012
rect 82081 3003 82139 3009
rect 83093 3009 83105 3043
rect 83139 3040 83151 3043
rect 83274 3040 83280 3052
rect 83139 3012 83280 3040
rect 83139 3009 83151 3012
rect 83093 3003 83151 3009
rect 74074 2932 74080 2984
rect 74132 2972 74138 2984
rect 75104 2972 75132 3000
rect 74132 2944 75132 2972
rect 74132 2932 74138 2944
rect 76190 2932 76196 2984
rect 76248 2972 76254 2984
rect 77864 2972 77892 3003
rect 83274 3000 83280 3012
rect 83332 3000 83338 3052
rect 84013 3043 84071 3049
rect 84013 3009 84025 3043
rect 84059 3040 84071 3043
rect 84194 3040 84200 3052
rect 84059 3012 84200 3040
rect 84059 3009 84071 3012
rect 84013 3003 84071 3009
rect 84194 3000 84200 3012
rect 84252 3040 84258 3052
rect 84930 3040 84936 3052
rect 84252 3012 84936 3040
rect 84252 3000 84258 3012
rect 84930 3000 84936 3012
rect 84988 3040 84994 3052
rect 85390 3040 85396 3052
rect 84988 3012 85396 3040
rect 84988 3000 84994 3012
rect 85390 3000 85396 3012
rect 85448 3040 85454 3052
rect 86129 3043 86187 3049
rect 86129 3040 86141 3043
rect 85448 3012 86141 3040
rect 85448 3000 85454 3012
rect 86129 3009 86141 3012
rect 86175 3009 86187 3043
rect 104526 3040 104532 3052
rect 104487 3012 104532 3040
rect 86129 3003 86187 3009
rect 104526 3000 104532 3012
rect 104584 3000 104590 3052
rect 76248 2944 77892 2972
rect 76248 2932 76254 2944
rect 78674 2932 78680 2984
rect 78732 2972 78738 2984
rect 79134 2972 79140 2984
rect 78732 2944 79140 2972
rect 78732 2932 78738 2944
rect 79134 2932 79140 2944
rect 79192 2972 79198 2984
rect 79229 2975 79287 2981
rect 79229 2972 79241 2975
rect 79192 2944 79241 2972
rect 79192 2932 79198 2944
rect 79229 2941 79241 2944
rect 79275 2941 79287 2975
rect 79229 2935 79287 2941
rect 79505 2975 79563 2981
rect 79505 2941 79517 2975
rect 79551 2972 79563 2975
rect 80238 2972 80244 2984
rect 79551 2944 80244 2972
rect 79551 2941 79563 2944
rect 79505 2935 79563 2941
rect 80238 2932 80244 2944
rect 80296 2932 80302 2984
rect 81986 2932 81992 2984
rect 82044 2972 82050 2984
rect 82265 2975 82323 2981
rect 82265 2972 82277 2975
rect 82044 2944 82277 2972
rect 82044 2932 82050 2944
rect 82265 2941 82277 2944
rect 82311 2941 82323 2975
rect 82265 2935 82323 2941
rect 83642 2932 83648 2984
rect 83700 2972 83706 2984
rect 85025 2975 85083 2981
rect 85025 2972 85037 2975
rect 83700 2944 85037 2972
rect 83700 2932 83706 2944
rect 85025 2941 85037 2944
rect 85071 2941 85083 2975
rect 85025 2935 85083 2941
rect 70026 2904 70032 2916
rect 66548 2876 70032 2904
rect 66548 2836 66576 2876
rect 70026 2864 70032 2876
rect 70084 2864 70090 2916
rect 70118 2864 70124 2916
rect 70176 2864 70182 2916
rect 71498 2864 71504 2916
rect 71556 2904 71562 2916
rect 72605 2907 72663 2913
rect 72605 2904 72617 2907
rect 71556 2876 72617 2904
rect 71556 2864 71562 2876
rect 72605 2873 72617 2876
rect 72651 2873 72663 2907
rect 72605 2867 72663 2873
rect 75181 2907 75239 2913
rect 75181 2873 75193 2907
rect 75227 2904 75239 2907
rect 76834 2904 76840 2916
rect 75227 2876 76840 2904
rect 75227 2873 75239 2876
rect 75181 2867 75239 2873
rect 76834 2864 76840 2876
rect 76892 2864 76898 2916
rect 84838 2904 84844 2916
rect 83108 2876 84844 2904
rect 64984 2808 66576 2836
rect 66993 2839 67051 2845
rect 66993 2805 67005 2839
rect 67039 2836 67051 2839
rect 67266 2836 67272 2848
rect 67039 2808 67272 2836
rect 67039 2805 67051 2808
rect 66993 2799 67051 2805
rect 67266 2796 67272 2808
rect 67324 2796 67330 2848
rect 67358 2796 67364 2848
rect 67416 2836 67422 2848
rect 67729 2839 67787 2845
rect 67729 2836 67741 2839
rect 67416 2808 67741 2836
rect 67416 2796 67422 2808
rect 67729 2805 67741 2808
rect 67775 2805 67787 2839
rect 67729 2799 67787 2805
rect 69661 2839 69719 2845
rect 69661 2805 69673 2839
rect 69707 2836 69719 2839
rect 71130 2836 71136 2848
rect 69707 2808 71136 2836
rect 69707 2805 69719 2808
rect 69661 2799 69719 2805
rect 71130 2796 71136 2808
rect 71188 2796 71194 2848
rect 73798 2796 73804 2848
rect 73856 2836 73862 2848
rect 74261 2839 74319 2845
rect 74261 2836 74273 2839
rect 73856 2808 74273 2836
rect 73856 2796 73862 2808
rect 74261 2805 74273 2808
rect 74307 2805 74319 2839
rect 74261 2799 74319 2805
rect 75638 2796 75644 2848
rect 75696 2836 75702 2848
rect 75917 2839 75975 2845
rect 75917 2836 75929 2839
rect 75696 2808 75929 2836
rect 75696 2796 75702 2808
rect 75917 2805 75929 2808
rect 75963 2805 75975 2839
rect 76466 2836 76472 2848
rect 76427 2808 76472 2836
rect 75917 2799 75975 2805
rect 76466 2796 76472 2808
rect 76524 2796 76530 2848
rect 76558 2796 76564 2848
rect 76616 2836 76622 2848
rect 83108 2836 83136 2876
rect 84838 2864 84844 2876
rect 84896 2864 84902 2916
rect 76616 2808 83136 2836
rect 76616 2796 76622 2808
rect 83182 2796 83188 2848
rect 83240 2836 83246 2848
rect 83921 2839 83979 2845
rect 83921 2836 83933 2839
rect 83240 2808 83933 2836
rect 83240 2796 83246 2808
rect 83921 2805 83933 2808
rect 83967 2805 83979 2839
rect 85666 2836 85672 2848
rect 85627 2808 85672 2836
rect 83921 2799 83979 2805
rect 85666 2796 85672 2808
rect 85724 2796 85730 2848
rect 97718 2836 97724 2848
rect 97679 2808 97724 2836
rect 97718 2796 97724 2808
rect 97776 2796 97782 2848
rect 101858 2836 101864 2848
rect 101819 2808 101864 2836
rect 101858 2796 101864 2808
rect 101916 2796 101922 2848
rect 110233 2839 110291 2845
rect 110233 2805 110245 2839
rect 110279 2836 110291 2839
rect 110414 2836 110420 2848
rect 110279 2808 110420 2836
rect 110279 2805 110291 2808
rect 110233 2799 110291 2805
rect 110414 2796 110420 2808
rect 110472 2796 110478 2848
rect 118418 2836 118424 2848
rect 118379 2808 118424 2836
rect 118418 2796 118424 2808
rect 118476 2796 118482 2848
rect 122558 2836 122564 2848
rect 122519 2808 122564 2836
rect 122558 2796 122564 2808
rect 122616 2796 122622 2848
rect 125321 2839 125379 2845
rect 125321 2805 125333 2839
rect 125367 2836 125379 2839
rect 125410 2836 125416 2848
rect 125367 2808 125416 2836
rect 125367 2805 125379 2808
rect 125321 2799 125379 2805
rect 125410 2796 125416 2808
rect 125468 2796 125474 2848
rect 130838 2836 130844 2848
rect 130799 2808 130844 2836
rect 130838 2796 130844 2808
rect 130896 2796 130902 2848
rect 143258 2836 143264 2848
rect 143219 2808 143264 2836
rect 143258 2796 143264 2808
rect 143316 2796 143322 2848
rect 1104 2746 148856 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 65654 2746
rect 65706 2694 65718 2746
rect 65770 2694 65782 2746
rect 65834 2694 65846 2746
rect 65898 2694 65910 2746
rect 65962 2694 96374 2746
rect 96426 2694 96438 2746
rect 96490 2694 96502 2746
rect 96554 2694 96566 2746
rect 96618 2694 96630 2746
rect 96682 2694 127094 2746
rect 127146 2694 127158 2746
rect 127210 2694 127222 2746
rect 127274 2694 127286 2746
rect 127338 2694 127350 2746
rect 127402 2694 148856 2746
rect 1104 2672 148856 2694
rect 4249 2635 4307 2641
rect 4249 2601 4261 2635
rect 4295 2632 4307 2635
rect 4614 2632 4620 2644
rect 4295 2604 4620 2632
rect 4295 2601 4307 2604
rect 4249 2595 4307 2601
rect 2869 2431 2927 2437
rect 2869 2397 2881 2431
rect 2915 2428 2927 2431
rect 4264 2428 4292 2595
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 9398 2592 9404 2644
rect 9456 2632 9462 2644
rect 9493 2635 9551 2641
rect 9493 2632 9505 2635
rect 9456 2604 9505 2632
rect 9456 2592 9462 2604
rect 9493 2601 9505 2604
rect 9539 2601 9551 2635
rect 14458 2632 14464 2644
rect 14419 2604 14464 2632
rect 9493 2595 9551 2601
rect 14458 2592 14464 2604
rect 14516 2592 14522 2644
rect 15378 2632 15384 2644
rect 15339 2604 15384 2632
rect 15378 2592 15384 2604
rect 15436 2592 15442 2644
rect 21266 2632 21272 2644
rect 21227 2604 21272 2632
rect 21266 2592 21272 2604
rect 21324 2592 21330 2644
rect 24762 2632 24768 2644
rect 24723 2604 24768 2632
rect 24762 2592 24768 2604
rect 24820 2592 24826 2644
rect 25682 2632 25688 2644
rect 25643 2604 25688 2632
rect 25682 2592 25688 2604
rect 25740 2592 25746 2644
rect 26510 2632 26516 2644
rect 26471 2604 26516 2632
rect 26510 2592 26516 2604
rect 26568 2592 26574 2644
rect 28902 2632 28908 2644
rect 28863 2604 28908 2632
rect 28902 2592 28908 2604
rect 28960 2592 28966 2644
rect 34057 2635 34115 2641
rect 34057 2601 34069 2635
rect 34103 2632 34115 2635
rect 34146 2632 34152 2644
rect 34103 2604 34152 2632
rect 34103 2601 34115 2604
rect 34057 2595 34115 2601
rect 34146 2592 34152 2604
rect 34204 2592 34210 2644
rect 36633 2635 36691 2641
rect 36633 2601 36645 2635
rect 36679 2632 36691 2635
rect 37090 2632 37096 2644
rect 36679 2604 37096 2632
rect 36679 2601 36691 2604
rect 36633 2595 36691 2601
rect 37090 2592 37096 2604
rect 37148 2592 37154 2644
rect 39206 2632 39212 2644
rect 39167 2604 39212 2632
rect 39206 2592 39212 2604
rect 39264 2592 39270 2644
rect 40034 2632 40040 2644
rect 39995 2604 40040 2632
rect 40034 2592 40040 2604
rect 40092 2592 40098 2644
rect 41325 2635 41383 2641
rect 41325 2601 41337 2635
rect 41371 2632 41383 2635
rect 41506 2632 41512 2644
rect 41371 2604 41512 2632
rect 41371 2601 41383 2604
rect 41325 2595 41383 2601
rect 41506 2592 41512 2604
rect 41564 2592 41570 2644
rect 44174 2592 44180 2644
rect 44232 2632 44238 2644
rect 44361 2635 44419 2641
rect 44361 2632 44373 2635
rect 44232 2604 44373 2632
rect 44232 2592 44238 2604
rect 44361 2601 44373 2604
rect 44407 2601 44419 2635
rect 47210 2632 47216 2644
rect 47171 2604 47216 2632
rect 44361 2595 44419 2601
rect 47210 2592 47216 2604
rect 47268 2592 47274 2644
rect 49510 2632 49516 2644
rect 49471 2604 49516 2632
rect 49510 2592 49516 2604
rect 49568 2592 49574 2644
rect 50614 2632 50620 2644
rect 50527 2604 50620 2632
rect 50614 2592 50620 2604
rect 50672 2632 50678 2644
rect 60826 2632 60832 2644
rect 50672 2604 60832 2632
rect 50672 2592 50678 2604
rect 60826 2592 60832 2604
rect 60884 2632 60890 2644
rect 62669 2635 62727 2641
rect 60884 2604 60964 2632
rect 60884 2592 60890 2604
rect 19705 2567 19763 2573
rect 19705 2533 19717 2567
rect 19751 2564 19763 2567
rect 19978 2564 19984 2576
rect 19751 2536 19984 2564
rect 19751 2533 19763 2536
rect 19705 2527 19763 2533
rect 19978 2524 19984 2536
rect 20036 2524 20042 2576
rect 20714 2564 20720 2576
rect 20675 2536 20720 2564
rect 20714 2524 20720 2536
rect 20772 2524 20778 2576
rect 39224 2564 39252 2592
rect 23860 2536 27292 2564
rect 39224 2536 41828 2564
rect 23860 2508 23888 2536
rect 5997 2499 6055 2505
rect 5997 2465 6009 2499
rect 6043 2496 6055 2499
rect 6362 2496 6368 2508
rect 6043 2468 6368 2496
rect 6043 2465 6055 2468
rect 5997 2459 6055 2465
rect 6362 2456 6368 2468
rect 6420 2496 6426 2508
rect 6549 2499 6607 2505
rect 6549 2496 6561 2499
rect 6420 2468 6561 2496
rect 6420 2456 6426 2468
rect 6549 2465 6561 2468
rect 6595 2496 6607 2499
rect 9214 2496 9220 2508
rect 6595 2468 9220 2496
rect 6595 2465 6607 2468
rect 6549 2459 6607 2465
rect 9214 2456 9220 2468
rect 9272 2496 9278 2508
rect 22005 2499 22063 2505
rect 22005 2496 22017 2499
rect 9272 2468 22017 2496
rect 9272 2456 9278 2468
rect 22005 2465 22017 2468
rect 22051 2496 22063 2499
rect 23842 2496 23848 2508
rect 22051 2468 23848 2496
rect 22051 2465 22063 2468
rect 22005 2459 22063 2465
rect 23842 2456 23848 2468
rect 23900 2456 23906 2508
rect 26234 2456 26240 2508
rect 26292 2496 26298 2508
rect 27157 2499 27215 2505
rect 27157 2496 27169 2499
rect 26292 2468 27169 2496
rect 26292 2456 26298 2468
rect 27157 2465 27169 2468
rect 27203 2465 27215 2499
rect 27264 2496 27292 2536
rect 29917 2499 29975 2505
rect 29917 2496 29929 2499
rect 27264 2468 29929 2496
rect 27157 2459 27215 2465
rect 29917 2465 29929 2468
rect 29963 2496 29975 2499
rect 32306 2496 32312 2508
rect 29963 2468 32312 2496
rect 29963 2465 29975 2468
rect 29917 2459 29975 2465
rect 32306 2456 32312 2468
rect 32364 2496 32370 2508
rect 34790 2496 34796 2508
rect 32364 2468 34796 2496
rect 32364 2456 32370 2468
rect 34790 2456 34796 2468
rect 34848 2496 34854 2508
rect 34885 2499 34943 2505
rect 34885 2496 34897 2499
rect 34848 2468 34897 2496
rect 34848 2456 34854 2468
rect 34885 2465 34897 2468
rect 34931 2465 34943 2499
rect 34885 2459 34943 2465
rect 37461 2499 37519 2505
rect 37461 2465 37473 2499
rect 37507 2496 37519 2499
rect 38470 2496 38476 2508
rect 37507 2468 38476 2496
rect 37507 2465 37519 2468
rect 37461 2459 37519 2465
rect 38470 2456 38476 2468
rect 38528 2456 38534 2508
rect 40589 2499 40647 2505
rect 40589 2465 40601 2499
rect 40635 2496 40647 2499
rect 41414 2496 41420 2508
rect 40635 2468 41420 2496
rect 40635 2465 40647 2468
rect 40589 2459 40647 2465
rect 41414 2456 41420 2468
rect 41472 2456 41478 2508
rect 2915 2400 4292 2428
rect 2915 2397 2927 2400
rect 2869 2391 2927 2397
rect 7926 2388 7932 2440
rect 7984 2388 7990 2440
rect 9398 2388 9404 2440
rect 9456 2428 9462 2440
rect 9677 2431 9735 2437
rect 9677 2428 9689 2431
rect 9456 2400 9689 2428
rect 9456 2388 9462 2400
rect 9677 2397 9689 2400
rect 9723 2428 9735 2431
rect 10137 2431 10195 2437
rect 10137 2428 10149 2431
rect 9723 2400 10149 2428
rect 9723 2397 9735 2400
rect 9677 2391 9735 2397
rect 10137 2397 10149 2400
rect 10183 2397 10195 2431
rect 10137 2391 10195 2397
rect 12529 2431 12587 2437
rect 12529 2397 12541 2431
rect 12575 2428 12587 2431
rect 12575 2400 14596 2428
rect 12575 2397 12587 2400
rect 12529 2391 12587 2397
rect 5626 2360 5632 2372
rect 5290 2332 5632 2360
rect 5626 2320 5632 2332
rect 5684 2320 5690 2372
rect 5721 2363 5779 2369
rect 5721 2329 5733 2363
rect 5767 2329 5779 2363
rect 6822 2360 6828 2372
rect 6783 2332 6828 2360
rect 5721 2323 5779 2329
rect 2498 2252 2504 2304
rect 2556 2292 2562 2304
rect 2685 2295 2743 2301
rect 2685 2292 2697 2295
rect 2556 2264 2697 2292
rect 2556 2252 2562 2264
rect 2685 2261 2697 2264
rect 2731 2261 2743 2295
rect 2685 2255 2743 2261
rect 3421 2295 3479 2301
rect 3421 2261 3433 2295
rect 3467 2292 3479 2295
rect 5350 2292 5356 2304
rect 3467 2264 5356 2292
rect 3467 2261 3479 2264
rect 3421 2255 3479 2261
rect 5350 2252 5356 2264
rect 5408 2292 5414 2304
rect 5736 2292 5764 2323
rect 6822 2320 6828 2332
rect 6880 2320 6886 2372
rect 8570 2360 8576 2372
rect 8531 2332 8576 2360
rect 8570 2320 8576 2332
rect 8628 2320 8634 2372
rect 14369 2363 14427 2369
rect 14369 2360 14381 2363
rect 13648 2332 14381 2360
rect 8588 2292 8616 2320
rect 5408 2264 8616 2292
rect 5408 2252 5414 2264
rect 12158 2252 12164 2304
rect 12216 2292 12222 2304
rect 12345 2295 12403 2301
rect 12345 2292 12357 2295
rect 12216 2264 12357 2292
rect 12216 2252 12222 2264
rect 12345 2261 12357 2264
rect 12391 2261 12403 2295
rect 12345 2255 12403 2261
rect 13538 2252 13544 2304
rect 13596 2292 13602 2304
rect 13648 2301 13676 2332
rect 14369 2329 14381 2332
rect 14415 2329 14427 2363
rect 14568 2360 14596 2400
rect 14918 2388 14924 2440
rect 14976 2428 14982 2440
rect 15197 2431 15255 2437
rect 15197 2428 15209 2431
rect 14976 2400 15209 2428
rect 14976 2388 14982 2400
rect 15197 2397 15209 2400
rect 15243 2397 15255 2431
rect 15197 2391 15255 2397
rect 18049 2431 18107 2437
rect 18049 2397 18061 2431
rect 18095 2428 18107 2431
rect 20622 2428 20628 2440
rect 18095 2400 20628 2428
rect 18095 2397 18107 2400
rect 18049 2391 18107 2397
rect 20622 2388 20628 2400
rect 20680 2388 20686 2440
rect 21450 2428 21456 2440
rect 21363 2400 21456 2428
rect 21450 2388 21456 2400
rect 21508 2428 21514 2440
rect 21818 2428 21824 2440
rect 21508 2400 21824 2428
rect 21508 2388 21514 2400
rect 21818 2388 21824 2400
rect 21876 2388 21882 2440
rect 26326 2388 26332 2440
rect 26384 2428 26390 2440
rect 30282 2428 30288 2440
rect 26384 2400 26556 2428
rect 30243 2400 30288 2428
rect 26384 2388 26390 2400
rect 19426 2360 19432 2372
rect 14568 2332 19432 2360
rect 14369 2323 14427 2329
rect 19426 2320 19432 2332
rect 19484 2320 19490 2372
rect 19521 2363 19579 2369
rect 19521 2329 19533 2363
rect 19567 2329 19579 2363
rect 19521 2323 19579 2329
rect 13633 2295 13691 2301
rect 13633 2292 13645 2295
rect 13596 2264 13645 2292
rect 13596 2252 13602 2264
rect 13633 2261 13645 2264
rect 13679 2261 13691 2295
rect 13633 2255 13691 2261
rect 17678 2252 17684 2304
rect 17736 2292 17742 2304
rect 17865 2295 17923 2301
rect 17865 2292 17877 2295
rect 17736 2264 17877 2292
rect 17736 2252 17742 2264
rect 17865 2261 17877 2264
rect 17911 2261 17923 2295
rect 17865 2255 17923 2261
rect 18877 2295 18935 2301
rect 18877 2261 18889 2295
rect 18923 2292 18935 2295
rect 19058 2292 19064 2304
rect 18923 2264 19064 2292
rect 18923 2261 18935 2264
rect 18877 2255 18935 2261
rect 19058 2252 19064 2264
rect 19116 2292 19122 2304
rect 19536 2292 19564 2323
rect 19610 2320 19616 2372
rect 19668 2320 19674 2372
rect 20438 2320 20444 2372
rect 20496 2360 20502 2372
rect 20533 2363 20591 2369
rect 20533 2360 20545 2363
rect 20496 2332 20545 2360
rect 20496 2320 20502 2332
rect 20533 2329 20545 2332
rect 20579 2329 20591 2363
rect 22278 2360 22284 2372
rect 22239 2332 22284 2360
rect 20533 2323 20591 2329
rect 22278 2320 22284 2332
rect 22336 2320 22342 2372
rect 22738 2320 22744 2372
rect 22796 2320 22802 2372
rect 24854 2360 24860 2372
rect 24815 2332 24860 2360
rect 24854 2320 24860 2332
rect 24912 2320 24918 2372
rect 25777 2363 25835 2369
rect 25777 2329 25789 2363
rect 25823 2360 25835 2363
rect 25958 2360 25964 2372
rect 25823 2332 25964 2360
rect 25823 2329 25835 2332
rect 25777 2323 25835 2329
rect 25958 2320 25964 2332
rect 26016 2320 26022 2372
rect 26418 2360 26424 2372
rect 26331 2332 26424 2360
rect 26418 2320 26424 2332
rect 26476 2320 26482 2372
rect 26528 2360 26556 2400
rect 30282 2388 30288 2400
rect 30340 2388 30346 2440
rect 31754 2428 31760 2440
rect 31715 2400 31760 2428
rect 31754 2388 31760 2400
rect 31812 2388 31818 2440
rect 40405 2431 40463 2437
rect 40405 2397 40417 2431
rect 40451 2428 40463 2431
rect 40678 2428 40684 2440
rect 40451 2400 40684 2428
rect 40451 2397 40463 2400
rect 40405 2391 40463 2397
rect 40678 2388 40684 2400
rect 40736 2388 40742 2440
rect 41800 2437 41828 2536
rect 42610 2496 42616 2508
rect 42571 2468 42616 2496
rect 42610 2456 42616 2468
rect 42668 2496 42674 2508
rect 45465 2499 45523 2505
rect 45465 2496 45477 2499
rect 42668 2468 45477 2496
rect 42668 2456 42674 2468
rect 45465 2465 45477 2468
rect 45511 2465 45523 2499
rect 45465 2459 45523 2465
rect 45741 2499 45799 2505
rect 45741 2465 45753 2499
rect 45787 2496 45799 2499
rect 46290 2496 46296 2508
rect 45787 2468 46296 2496
rect 45787 2465 45799 2468
rect 45741 2459 45799 2465
rect 46290 2456 46296 2468
rect 46348 2456 46354 2508
rect 47762 2496 47768 2508
rect 47723 2468 47768 2496
rect 47762 2456 47768 2468
rect 47820 2456 47826 2508
rect 50632 2505 50660 2592
rect 52365 2567 52423 2573
rect 52365 2533 52377 2567
rect 52411 2564 52423 2567
rect 53282 2564 53288 2576
rect 52411 2536 53288 2564
rect 52411 2533 52423 2536
rect 52365 2527 52423 2533
rect 53282 2524 53288 2536
rect 53340 2524 53346 2576
rect 53561 2567 53619 2573
rect 53561 2533 53573 2567
rect 53607 2564 53619 2567
rect 54938 2564 54944 2576
rect 53607 2536 54944 2564
rect 53607 2533 53619 2536
rect 53561 2527 53619 2533
rect 54938 2524 54944 2536
rect 54996 2524 55002 2576
rect 50617 2499 50675 2505
rect 50617 2465 50629 2499
rect 50663 2465 50675 2499
rect 50617 2459 50675 2465
rect 50893 2499 50951 2505
rect 50893 2465 50905 2499
rect 50939 2496 50951 2499
rect 51534 2496 51540 2508
rect 50939 2468 51540 2496
rect 50939 2465 50951 2468
rect 50893 2459 50951 2465
rect 51534 2456 51540 2468
rect 51592 2456 51598 2508
rect 51902 2456 51908 2508
rect 51960 2496 51966 2508
rect 54202 2496 54208 2508
rect 51960 2468 53420 2496
rect 54115 2468 54208 2496
rect 51960 2456 51966 2468
rect 53392 2437 53420 2468
rect 54202 2456 54208 2468
rect 54260 2496 54266 2508
rect 55122 2496 55128 2508
rect 54260 2468 55128 2496
rect 54260 2456 54266 2468
rect 55122 2456 55128 2468
rect 55180 2456 55186 2508
rect 55674 2496 55680 2508
rect 55587 2468 55680 2496
rect 55674 2456 55680 2468
rect 55732 2496 55738 2508
rect 58069 2499 58127 2505
rect 58069 2496 58081 2499
rect 55732 2468 58081 2496
rect 55732 2456 55738 2468
rect 58069 2465 58081 2468
rect 58115 2496 58127 2499
rect 58710 2496 58716 2508
rect 58115 2468 58716 2496
rect 58115 2465 58127 2468
rect 58069 2459 58127 2465
rect 58710 2456 58716 2468
rect 58768 2456 58774 2508
rect 60936 2505 60964 2604
rect 62669 2601 62681 2635
rect 62715 2632 62727 2635
rect 63586 2632 63592 2644
rect 62715 2604 63592 2632
rect 62715 2601 62727 2604
rect 62669 2595 62727 2601
rect 63586 2592 63592 2604
rect 63644 2592 63650 2644
rect 64969 2635 65027 2641
rect 64969 2601 64981 2635
rect 65015 2632 65027 2635
rect 65058 2632 65064 2644
rect 65015 2604 65064 2632
rect 65015 2601 65027 2604
rect 64969 2595 65027 2601
rect 65058 2592 65064 2604
rect 65116 2592 65122 2644
rect 69014 2632 69020 2644
rect 68975 2604 69020 2632
rect 69014 2592 69020 2604
rect 69072 2592 69078 2644
rect 69106 2592 69112 2644
rect 69164 2632 69170 2644
rect 70118 2632 70124 2644
rect 69164 2604 70124 2632
rect 69164 2592 69170 2604
rect 70118 2592 70124 2604
rect 70176 2632 70182 2644
rect 70946 2632 70952 2644
rect 70176 2604 70952 2632
rect 70176 2592 70182 2604
rect 70946 2592 70952 2604
rect 71004 2632 71010 2644
rect 71004 2604 81296 2632
rect 71004 2592 71010 2604
rect 68830 2524 68836 2576
rect 68888 2564 68894 2576
rect 69661 2567 69719 2573
rect 68888 2536 69612 2564
rect 68888 2524 68894 2536
rect 60921 2499 60979 2505
rect 60921 2465 60933 2499
rect 60967 2496 60979 2499
rect 63221 2499 63279 2505
rect 63221 2496 63233 2499
rect 60967 2468 63233 2496
rect 60967 2465 60979 2468
rect 60921 2459 60979 2465
rect 63221 2465 63233 2468
rect 63267 2496 63279 2499
rect 65797 2499 65855 2505
rect 65797 2496 65809 2499
rect 63267 2468 65809 2496
rect 63267 2465 63279 2468
rect 63221 2459 63279 2465
rect 65797 2465 65809 2468
rect 65843 2496 65855 2499
rect 69106 2496 69112 2508
rect 65843 2468 69112 2496
rect 65843 2465 65855 2468
rect 65797 2459 65855 2465
rect 69106 2456 69112 2468
rect 69164 2456 69170 2508
rect 41785 2431 41843 2437
rect 41785 2397 41797 2431
rect 41831 2397 41843 2431
rect 41785 2391 41843 2397
rect 53377 2431 53435 2437
rect 53377 2397 53389 2431
rect 53423 2397 53435 2431
rect 53377 2391 53435 2397
rect 54294 2388 54300 2440
rect 54352 2428 54358 2440
rect 54481 2431 54539 2437
rect 54481 2428 54493 2431
rect 54352 2400 54493 2428
rect 54352 2388 54358 2400
rect 54481 2397 54493 2400
rect 54527 2397 54539 2431
rect 54481 2391 54539 2397
rect 62298 2388 62304 2440
rect 62356 2388 62362 2440
rect 69584 2437 69612 2536
rect 69661 2533 69673 2567
rect 69707 2564 69719 2567
rect 70486 2564 70492 2576
rect 69707 2536 70492 2564
rect 69707 2533 69719 2536
rect 69661 2527 69719 2533
rect 70486 2524 70492 2536
rect 70544 2524 70550 2576
rect 70946 2456 70952 2508
rect 71004 2496 71010 2508
rect 73522 2496 73528 2508
rect 71004 2468 71049 2496
rect 73483 2468 73528 2496
rect 71004 2456 71010 2468
rect 73522 2456 73528 2468
rect 73580 2496 73586 2508
rect 76101 2499 76159 2505
rect 76101 2496 76113 2499
rect 73580 2468 76113 2496
rect 73580 2456 73586 2468
rect 76101 2465 76113 2468
rect 76147 2496 76159 2499
rect 76466 2496 76472 2508
rect 76147 2468 76472 2496
rect 76147 2465 76159 2468
rect 76101 2459 76159 2465
rect 76466 2456 76472 2468
rect 76524 2496 76530 2508
rect 78674 2496 78680 2508
rect 76524 2468 78680 2496
rect 76524 2456 76530 2468
rect 78674 2456 78680 2468
rect 78732 2456 78738 2508
rect 78953 2499 79011 2505
rect 78953 2465 78965 2499
rect 78999 2496 79011 2499
rect 80238 2496 80244 2508
rect 78999 2468 80244 2496
rect 78999 2465 79011 2468
rect 78953 2459 79011 2465
rect 80238 2456 80244 2468
rect 80296 2456 80302 2508
rect 81268 2505 81296 2604
rect 81342 2592 81348 2644
rect 81400 2632 81406 2644
rect 85482 2632 85488 2644
rect 81400 2604 84516 2632
rect 85443 2604 85488 2632
rect 81400 2592 81406 2604
rect 82906 2524 82912 2576
rect 82964 2564 82970 2576
rect 84102 2564 84108 2576
rect 82964 2536 84108 2564
rect 82964 2524 82970 2536
rect 84102 2524 84108 2536
rect 84160 2524 84166 2576
rect 81253 2499 81311 2505
rect 81253 2465 81265 2499
rect 81299 2496 81311 2499
rect 84194 2496 84200 2508
rect 81299 2468 84200 2496
rect 81299 2465 81311 2468
rect 81253 2459 81311 2465
rect 84194 2456 84200 2468
rect 84252 2456 84258 2508
rect 69569 2431 69627 2437
rect 67468 2400 69060 2428
rect 27433 2363 27491 2369
rect 27433 2360 27445 2363
rect 26528 2332 27445 2360
rect 27433 2329 27445 2332
rect 27479 2329 27491 2363
rect 27433 2323 27491 2329
rect 27890 2320 27896 2372
rect 27948 2320 27954 2372
rect 30742 2320 30748 2372
rect 30800 2320 30806 2372
rect 32585 2363 32643 2369
rect 32585 2329 32597 2363
rect 32631 2329 32643 2363
rect 32585 2323 32643 2329
rect 19116 2264 19564 2292
rect 19628 2292 19656 2320
rect 23106 2292 23112 2304
rect 19628 2264 23112 2292
rect 19116 2252 19122 2264
rect 23106 2252 23112 2264
rect 23164 2292 23170 2304
rect 23753 2295 23811 2301
rect 23753 2292 23765 2295
rect 23164 2264 23765 2292
rect 23164 2252 23170 2264
rect 23753 2261 23765 2264
rect 23799 2261 23811 2295
rect 26436 2292 26464 2320
rect 27338 2292 27344 2304
rect 26436 2264 27344 2292
rect 23753 2255 23811 2261
rect 27338 2252 27344 2264
rect 27396 2252 27402 2304
rect 32600 2292 32628 2323
rect 33318 2320 33324 2372
rect 33376 2320 33382 2372
rect 34698 2320 34704 2372
rect 34756 2360 34762 2372
rect 35161 2363 35219 2369
rect 35161 2360 35173 2363
rect 34756 2332 35173 2360
rect 34756 2320 34762 2332
rect 35161 2329 35173 2332
rect 35207 2329 35219 2363
rect 35161 2323 35219 2329
rect 35894 2320 35900 2372
rect 35952 2320 35958 2372
rect 37734 2360 37740 2372
rect 37695 2332 37740 2360
rect 37734 2320 37740 2332
rect 37792 2320 37798 2372
rect 38746 2320 38752 2372
rect 38804 2320 38810 2372
rect 40497 2363 40555 2369
rect 40497 2329 40509 2363
rect 40543 2360 40555 2363
rect 40586 2360 40592 2372
rect 40543 2332 40592 2360
rect 40543 2329 40555 2332
rect 40497 2323 40555 2329
rect 40586 2320 40592 2332
rect 40644 2320 40650 2372
rect 42886 2360 42892 2372
rect 42847 2332 42892 2360
rect 42886 2320 42892 2332
rect 42944 2320 42950 2372
rect 45278 2360 45284 2372
rect 44114 2332 45284 2360
rect 45278 2320 45284 2332
rect 45336 2320 45342 2372
rect 46198 2320 46204 2372
rect 46256 2320 46262 2372
rect 47670 2320 47676 2372
rect 47728 2360 47734 2372
rect 48041 2363 48099 2369
rect 48041 2360 48053 2363
rect 47728 2332 48053 2360
rect 47728 2320 47734 2332
rect 48041 2329 48053 2332
rect 48087 2329 48099 2363
rect 50062 2360 50068 2372
rect 49266 2332 50068 2360
rect 48041 2323 48099 2329
rect 50062 2320 50068 2332
rect 50120 2320 50126 2372
rect 52270 2360 52276 2372
rect 52118 2332 52276 2360
rect 52270 2320 52276 2332
rect 52328 2320 52334 2372
rect 55953 2363 56011 2369
rect 55953 2329 55965 2363
rect 55999 2329 56011 2363
rect 55953 2323 56011 2329
rect 33870 2292 33876 2304
rect 32600 2264 33876 2292
rect 33870 2252 33876 2264
rect 33928 2252 33934 2304
rect 41969 2295 42027 2301
rect 41969 2261 41981 2295
rect 42015 2292 42027 2295
rect 42518 2292 42524 2304
rect 42015 2264 42524 2292
rect 42015 2261 42027 2264
rect 41969 2255 42027 2261
rect 42518 2252 42524 2264
rect 42576 2252 42582 2304
rect 55968 2292 55996 2323
rect 56686 2320 56692 2372
rect 56744 2320 56750 2372
rect 58342 2360 58348 2372
rect 58303 2332 58348 2360
rect 58342 2320 58348 2332
rect 58400 2320 58406 2372
rect 59354 2320 59360 2372
rect 59412 2320 59418 2372
rect 61194 2360 61200 2372
rect 61155 2332 61200 2360
rect 61194 2320 61200 2332
rect 61252 2320 61258 2372
rect 63494 2360 63500 2372
rect 63455 2332 63500 2360
rect 63494 2320 63500 2332
rect 63552 2320 63558 2372
rect 63954 2320 63960 2372
rect 64012 2320 64018 2372
rect 65242 2320 65248 2372
rect 65300 2360 65306 2372
rect 66073 2363 66131 2369
rect 66073 2360 66085 2363
rect 65300 2332 66085 2360
rect 65300 2320 65306 2332
rect 66073 2329 66085 2332
rect 66119 2329 66131 2363
rect 66073 2323 66131 2329
rect 66530 2320 66536 2372
rect 66588 2320 66594 2372
rect 56594 2292 56600 2304
rect 55968 2264 56600 2292
rect 56594 2252 56600 2264
rect 56652 2252 56658 2304
rect 57422 2292 57428 2304
rect 57383 2264 57428 2292
rect 57422 2252 57428 2264
rect 57480 2252 57486 2304
rect 59814 2292 59820 2304
rect 59775 2264 59820 2292
rect 59814 2252 59820 2264
rect 59872 2252 59878 2304
rect 61470 2252 61476 2304
rect 61528 2292 61534 2304
rect 67468 2292 67496 2400
rect 68922 2360 68928 2372
rect 68883 2332 68928 2360
rect 68922 2320 68928 2332
rect 68980 2320 68986 2372
rect 69032 2360 69060 2400
rect 69569 2397 69581 2431
rect 69615 2428 69627 2431
rect 70213 2431 70271 2437
rect 70213 2428 70225 2431
rect 69615 2400 70225 2428
rect 69615 2397 69627 2400
rect 69569 2391 69627 2397
rect 70213 2397 70225 2400
rect 70259 2397 70271 2431
rect 70213 2391 70271 2397
rect 75549 2431 75607 2437
rect 75549 2397 75561 2431
rect 75595 2428 75607 2431
rect 75822 2428 75828 2440
rect 75595 2400 75828 2428
rect 75595 2397 75607 2400
rect 75549 2391 75607 2397
rect 75822 2388 75828 2400
rect 75880 2388 75886 2440
rect 80790 2428 80796 2440
rect 80086 2400 80796 2428
rect 80790 2388 80796 2400
rect 80848 2388 80854 2440
rect 82814 2388 82820 2440
rect 82872 2428 82878 2440
rect 84289 2431 84347 2437
rect 82872 2400 84194 2428
rect 82872 2388 82878 2400
rect 69032 2332 71084 2360
rect 61528 2264 67496 2292
rect 61528 2252 61534 2264
rect 67542 2252 67548 2304
rect 67600 2292 67606 2304
rect 70305 2295 70363 2301
rect 67600 2264 67645 2292
rect 67600 2252 67606 2264
rect 70305 2261 70317 2295
rect 70351 2292 70363 2295
rect 70946 2292 70952 2304
rect 70351 2264 70952 2292
rect 70351 2261 70363 2264
rect 70305 2255 70363 2261
rect 70946 2252 70952 2264
rect 71004 2252 71010 2304
rect 71056 2292 71084 2332
rect 71130 2320 71136 2372
rect 71188 2360 71194 2372
rect 71225 2363 71283 2369
rect 71225 2360 71237 2363
rect 71188 2332 71237 2360
rect 71188 2320 71194 2332
rect 71225 2329 71237 2332
rect 71271 2329 71283 2363
rect 71225 2323 71283 2329
rect 71682 2320 71688 2372
rect 71740 2320 71746 2372
rect 73798 2360 73804 2372
rect 72528 2332 73660 2360
rect 73759 2332 73804 2360
rect 72528 2292 72556 2332
rect 72694 2292 72700 2304
rect 71056 2264 72556 2292
rect 72655 2264 72700 2292
rect 72694 2252 72700 2264
rect 72752 2252 72758 2304
rect 73632 2292 73660 2332
rect 73798 2320 73804 2332
rect 73856 2320 73862 2372
rect 74534 2320 74540 2372
rect 74592 2320 74598 2372
rect 76374 2360 76380 2372
rect 76335 2332 76380 2360
rect 76374 2320 76380 2332
rect 76432 2320 76438 2372
rect 76834 2320 76840 2372
rect 76892 2320 76898 2372
rect 78122 2360 78128 2372
rect 78083 2332 78128 2360
rect 78122 2320 78128 2332
rect 78180 2320 78186 2372
rect 80701 2363 80759 2369
rect 80701 2329 80713 2363
rect 80747 2360 80759 2363
rect 81529 2363 81587 2369
rect 80747 2332 81480 2360
rect 80747 2329 80759 2332
rect 80701 2323 80759 2329
rect 81342 2292 81348 2304
rect 73632 2264 81348 2292
rect 81342 2252 81348 2264
rect 81400 2252 81406 2304
rect 81452 2292 81480 2332
rect 81529 2329 81541 2363
rect 81575 2360 81587 2363
rect 81618 2360 81624 2372
rect 81575 2332 81624 2360
rect 81575 2329 81587 2332
rect 81529 2323 81587 2329
rect 81618 2320 81624 2332
rect 81676 2320 81682 2372
rect 83090 2360 83096 2372
rect 82754 2332 83096 2360
rect 83090 2320 83096 2332
rect 83148 2320 83154 2372
rect 84166 2360 84194 2400
rect 84289 2397 84301 2431
rect 84335 2428 84347 2431
rect 84488 2428 84516 2604
rect 85482 2592 85488 2604
rect 85540 2592 85546 2644
rect 89714 2632 89720 2644
rect 89675 2604 89720 2632
rect 89714 2592 89720 2604
rect 89772 2592 89778 2644
rect 94314 2632 94320 2644
rect 94275 2604 94320 2632
rect 94314 2592 94320 2604
rect 94372 2592 94378 2644
rect 97810 2592 97816 2644
rect 97868 2632 97874 2644
rect 97997 2635 98055 2641
rect 97997 2632 98009 2635
rect 97868 2604 98009 2632
rect 97868 2592 97874 2604
rect 97997 2601 98009 2604
rect 98043 2601 98055 2635
rect 102134 2632 102140 2644
rect 102095 2604 102140 2632
rect 97997 2595 98055 2601
rect 102134 2592 102140 2604
rect 102192 2592 102198 2644
rect 106274 2632 106280 2644
rect 106235 2604 106280 2632
rect 106274 2592 106280 2604
rect 106332 2592 106338 2644
rect 110506 2632 110512 2644
rect 110467 2604 110512 2632
rect 110506 2592 110512 2604
rect 110564 2592 110570 2644
rect 114830 2592 114836 2644
rect 114888 2632 114894 2644
rect 114925 2635 114983 2641
rect 114925 2632 114937 2635
rect 114888 2604 114937 2632
rect 114888 2592 114894 2604
rect 114925 2601 114937 2604
rect 114971 2601 114983 2635
rect 118694 2632 118700 2644
rect 118655 2604 118700 2632
rect 114925 2595 114983 2601
rect 118694 2592 118700 2604
rect 118752 2592 118758 2644
rect 122834 2592 122840 2644
rect 122892 2632 122898 2644
rect 126974 2632 126980 2644
rect 122892 2604 122937 2632
rect 126935 2604 126980 2632
rect 122892 2592 122898 2604
rect 126974 2592 126980 2604
rect 127032 2592 127038 2644
rect 131114 2632 131120 2644
rect 131075 2604 131120 2632
rect 131114 2592 131120 2604
rect 131172 2592 131178 2644
rect 137278 2632 137284 2644
rect 137239 2604 137284 2632
rect 137278 2592 137284 2604
rect 137336 2592 137342 2644
rect 139397 2635 139455 2641
rect 139397 2601 139409 2635
rect 139443 2632 139455 2635
rect 141326 2632 141332 2644
rect 139443 2604 141332 2632
rect 139443 2601 139455 2604
rect 139397 2595 139455 2601
rect 141326 2592 141332 2604
rect 141384 2592 141390 2644
rect 143534 2632 143540 2644
rect 143495 2604 143540 2632
rect 143534 2592 143540 2604
rect 143592 2592 143598 2644
rect 147306 2632 147312 2644
rect 147267 2604 147312 2632
rect 147306 2592 147312 2604
rect 147364 2592 147370 2644
rect 108758 2524 108764 2576
rect 108816 2564 108822 2576
rect 109773 2567 109831 2573
rect 109773 2564 109785 2567
rect 108816 2536 109785 2564
rect 108816 2524 108822 2536
rect 109773 2533 109785 2536
rect 109819 2533 109831 2567
rect 109773 2527 109831 2533
rect 117222 2524 117228 2576
rect 117280 2564 117286 2576
rect 129553 2567 129611 2573
rect 129553 2564 129565 2567
rect 117280 2536 129565 2564
rect 117280 2524 117286 2536
rect 129553 2533 129565 2536
rect 129599 2533 129611 2567
rect 129553 2527 129611 2533
rect 135533 2567 135591 2573
rect 135533 2533 135545 2567
rect 135579 2564 135591 2567
rect 139486 2564 139492 2576
rect 135579 2536 139492 2564
rect 135579 2533 135591 2536
rect 135533 2527 135591 2533
rect 86497 2499 86555 2505
rect 86497 2496 86509 2499
rect 84764 2468 86509 2496
rect 84764 2428 84792 2468
rect 86497 2465 86509 2468
rect 86543 2465 86555 2499
rect 86497 2459 86555 2465
rect 108298 2456 108304 2508
rect 108356 2496 108362 2508
rect 120721 2499 120779 2505
rect 120721 2496 120733 2499
rect 108356 2468 120733 2496
rect 108356 2456 108362 2468
rect 120721 2465 120733 2468
rect 120767 2465 120779 2499
rect 120721 2459 120779 2465
rect 84930 2428 84936 2440
rect 84335 2400 84792 2428
rect 84891 2400 84936 2428
rect 84335 2397 84347 2400
rect 84289 2391 84347 2397
rect 84930 2388 84936 2400
rect 84988 2388 84994 2440
rect 88153 2431 88211 2437
rect 88153 2428 88165 2431
rect 87616 2400 88165 2428
rect 84841 2363 84899 2369
rect 84841 2360 84853 2363
rect 84166 2332 84853 2360
rect 84841 2329 84853 2332
rect 84887 2329 84899 2363
rect 84841 2323 84899 2329
rect 85298 2320 85304 2372
rect 85356 2360 85362 2372
rect 85577 2363 85635 2369
rect 85577 2360 85589 2363
rect 85356 2332 85589 2360
rect 85356 2320 85362 2332
rect 85577 2329 85589 2332
rect 85623 2360 85635 2363
rect 86957 2363 87015 2369
rect 86957 2360 86969 2363
rect 85623 2332 86969 2360
rect 85623 2329 85635 2332
rect 85577 2323 85635 2329
rect 86957 2329 86969 2332
rect 87003 2329 87015 2363
rect 86957 2323 87015 2329
rect 87616 2304 87644 2400
rect 88153 2397 88165 2400
rect 88199 2397 88211 2431
rect 92293 2431 92351 2437
rect 92293 2428 92305 2431
rect 88153 2391 88211 2397
rect 91756 2400 92305 2428
rect 89073 2363 89131 2369
rect 89073 2329 89085 2363
rect 89119 2360 89131 2363
rect 89438 2360 89444 2372
rect 89119 2332 89444 2360
rect 89119 2329 89131 2332
rect 89073 2323 89131 2329
rect 89438 2320 89444 2332
rect 89496 2360 89502 2372
rect 89625 2363 89683 2369
rect 89625 2360 89637 2363
rect 89496 2332 89637 2360
rect 89496 2320 89502 2332
rect 89625 2329 89637 2332
rect 89671 2329 89683 2363
rect 89625 2323 89683 2329
rect 91756 2304 91784 2400
rect 92293 2397 92305 2400
rect 92339 2397 92351 2431
rect 96709 2431 96767 2437
rect 96709 2428 96721 2431
rect 92293 2391 92351 2397
rect 96080 2400 96721 2428
rect 94225 2363 94283 2369
rect 94225 2360 94237 2363
rect 93826 2332 94237 2360
rect 82814 2292 82820 2304
rect 81452 2264 82820 2292
rect 82814 2252 82820 2264
rect 82872 2252 82878 2304
rect 82998 2292 83004 2304
rect 82959 2264 83004 2292
rect 82998 2252 83004 2264
rect 83056 2252 83062 2304
rect 83918 2252 83924 2304
rect 83976 2292 83982 2304
rect 84105 2295 84163 2301
rect 84105 2292 84117 2295
rect 83976 2264 84117 2292
rect 83976 2252 83982 2264
rect 84105 2261 84117 2264
rect 84151 2261 84163 2295
rect 84105 2255 84163 2261
rect 84194 2252 84200 2304
rect 84252 2292 84258 2304
rect 85666 2292 85672 2304
rect 84252 2264 85672 2292
rect 84252 2252 84258 2264
rect 85666 2252 85672 2264
rect 85724 2252 85730 2304
rect 87598 2292 87604 2304
rect 87559 2264 87604 2292
rect 87598 2252 87604 2264
rect 87656 2252 87662 2304
rect 88058 2252 88064 2304
rect 88116 2292 88122 2304
rect 88337 2295 88395 2301
rect 88337 2292 88349 2295
rect 88116 2264 88349 2292
rect 88116 2252 88122 2264
rect 88337 2261 88349 2264
rect 88383 2261 88395 2295
rect 91738 2292 91744 2304
rect 91699 2264 91744 2292
rect 88337 2255 88395 2261
rect 91738 2252 91744 2264
rect 91796 2252 91802 2304
rect 92198 2252 92204 2304
rect 92256 2292 92262 2304
rect 92477 2295 92535 2301
rect 92477 2292 92489 2295
rect 92256 2264 92489 2292
rect 92256 2252 92262 2264
rect 92477 2261 92489 2264
rect 92523 2261 92535 2295
rect 93578 2292 93584 2304
rect 93539 2264 93584 2292
rect 92477 2255 92535 2261
rect 93578 2252 93584 2264
rect 93636 2292 93642 2304
rect 93826 2292 93854 2332
rect 94225 2329 94237 2332
rect 94271 2329 94283 2363
rect 94225 2323 94283 2329
rect 96080 2304 96108 2400
rect 96709 2397 96721 2400
rect 96755 2397 96767 2431
rect 100573 2431 100631 2437
rect 100573 2428 100585 2431
rect 96709 2391 96767 2397
rect 100036 2400 100585 2428
rect 97718 2320 97724 2372
rect 97776 2360 97782 2372
rect 97905 2363 97963 2369
rect 97905 2360 97917 2363
rect 97776 2332 97917 2360
rect 97776 2320 97782 2332
rect 97905 2329 97917 2332
rect 97951 2329 97963 2363
rect 97905 2323 97963 2329
rect 100036 2304 100064 2400
rect 100573 2397 100585 2400
rect 100619 2397 100631 2431
rect 100573 2391 100631 2397
rect 104526 2388 104532 2440
rect 104584 2428 104590 2440
rect 104713 2431 104771 2437
rect 104713 2428 104725 2431
rect 104584 2400 104725 2428
rect 104584 2388 104590 2400
rect 104713 2397 104725 2400
rect 104759 2397 104771 2431
rect 109589 2431 109647 2437
rect 109589 2428 109601 2431
rect 104713 2391 104771 2397
rect 109052 2400 109601 2428
rect 101858 2320 101864 2372
rect 101916 2360 101922 2372
rect 102045 2363 102103 2369
rect 102045 2360 102057 2363
rect 101916 2332 102057 2360
rect 101916 2320 101922 2332
rect 102045 2329 102057 2332
rect 102091 2329 102103 2363
rect 102045 2323 102103 2329
rect 105633 2363 105691 2369
rect 105633 2329 105645 2363
rect 105679 2360 105691 2363
rect 105998 2360 106004 2372
rect 105679 2332 106004 2360
rect 105679 2329 105691 2332
rect 105633 2323 105691 2329
rect 105998 2320 106004 2332
rect 106056 2360 106062 2372
rect 106185 2363 106243 2369
rect 106185 2360 106197 2363
rect 106056 2332 106197 2360
rect 106056 2320 106062 2332
rect 106185 2329 106197 2332
rect 106231 2329 106243 2363
rect 106185 2323 106243 2329
rect 109052 2304 109080 2400
rect 109589 2397 109601 2400
rect 109635 2397 109647 2431
rect 112993 2431 113051 2437
rect 112993 2428 113005 2431
rect 109589 2391 109647 2397
rect 112456 2400 113005 2428
rect 110414 2360 110420 2372
rect 110375 2332 110420 2360
rect 110414 2320 110420 2332
rect 110472 2320 110478 2372
rect 112456 2304 112484 2400
rect 112993 2397 113005 2400
rect 113039 2397 113051 2431
rect 117317 2431 117375 2437
rect 117317 2428 117329 2431
rect 112993 2391 113051 2397
rect 116688 2400 117329 2428
rect 114833 2363 114891 2369
rect 114833 2329 114845 2363
rect 114879 2329 114891 2363
rect 114833 2323 114891 2329
rect 96062 2292 96068 2304
rect 93636 2264 93854 2292
rect 96023 2264 96068 2292
rect 93636 2252 93642 2264
rect 96062 2252 96068 2264
rect 96120 2252 96126 2304
rect 96338 2252 96344 2304
rect 96396 2292 96402 2304
rect 96893 2295 96951 2301
rect 96893 2292 96905 2295
rect 96396 2264 96905 2292
rect 96396 2252 96402 2264
rect 96893 2261 96905 2264
rect 96939 2261 96951 2295
rect 100018 2292 100024 2304
rect 99979 2264 100024 2292
rect 96893 2255 96951 2261
rect 100018 2252 100024 2264
rect 100076 2252 100082 2304
rect 100478 2252 100484 2304
rect 100536 2292 100542 2304
rect 100757 2295 100815 2301
rect 100757 2292 100769 2295
rect 100536 2264 100769 2292
rect 100536 2252 100542 2264
rect 100757 2261 100769 2264
rect 100803 2261 100815 2295
rect 100757 2255 100815 2261
rect 104618 2252 104624 2304
rect 104676 2292 104682 2304
rect 104897 2295 104955 2301
rect 104897 2292 104909 2295
rect 104676 2264 104909 2292
rect 104676 2252 104682 2264
rect 104897 2261 104909 2264
rect 104943 2261 104955 2295
rect 109034 2292 109040 2304
rect 108995 2264 109040 2292
rect 104897 2255 104955 2261
rect 109034 2252 109040 2264
rect 109092 2252 109098 2304
rect 112438 2292 112444 2304
rect 112399 2264 112444 2292
rect 112438 2252 112444 2264
rect 112496 2252 112502 2304
rect 112898 2252 112904 2304
rect 112956 2292 112962 2304
rect 113177 2295 113235 2301
rect 113177 2292 113189 2295
rect 112956 2264 113189 2292
rect 112956 2252 112962 2264
rect 113177 2261 113189 2264
rect 113223 2261 113235 2295
rect 113177 2255 113235 2261
rect 114189 2295 114247 2301
rect 114189 2261 114201 2295
rect 114235 2292 114247 2295
rect 114278 2292 114284 2304
rect 114235 2264 114284 2292
rect 114235 2261 114247 2264
rect 114189 2255 114247 2261
rect 114278 2252 114284 2264
rect 114336 2292 114342 2304
rect 114848 2292 114876 2323
rect 116688 2304 116716 2400
rect 117317 2397 117329 2400
rect 117363 2397 117375 2431
rect 120736 2428 120764 2459
rect 121273 2431 121331 2437
rect 121273 2428 121285 2431
rect 120736 2400 121285 2428
rect 117317 2391 117375 2397
rect 121273 2397 121285 2400
rect 121319 2397 121331 2431
rect 125410 2428 125416 2440
rect 125371 2400 125416 2428
rect 121273 2391 121331 2397
rect 125410 2388 125416 2400
rect 125468 2388 125474 2440
rect 125502 2388 125508 2440
rect 125560 2428 125566 2440
rect 129568 2428 129596 2527
rect 139486 2524 139492 2536
rect 139544 2524 139550 2576
rect 130197 2431 130255 2437
rect 130197 2428 130209 2431
rect 125560 2400 127664 2428
rect 129568 2400 130209 2428
rect 125560 2388 125566 2400
rect 118418 2320 118424 2372
rect 118476 2360 118482 2372
rect 118605 2363 118663 2369
rect 118605 2360 118617 2363
rect 118476 2332 118617 2360
rect 118476 2320 118482 2332
rect 118605 2329 118617 2332
rect 118651 2329 118663 2363
rect 118605 2323 118663 2329
rect 122558 2320 122564 2372
rect 122616 2360 122622 2372
rect 122745 2363 122803 2369
rect 122745 2360 122757 2363
rect 122616 2332 122757 2360
rect 122616 2320 122622 2332
rect 122745 2329 122757 2332
rect 122791 2329 122803 2363
rect 122745 2323 122803 2329
rect 126333 2363 126391 2369
rect 126333 2329 126345 2363
rect 126379 2360 126391 2363
rect 126698 2360 126704 2372
rect 126379 2332 126704 2360
rect 126379 2329 126391 2332
rect 126333 2323 126391 2329
rect 126698 2320 126704 2332
rect 126756 2360 126762 2372
rect 126885 2363 126943 2369
rect 126885 2360 126897 2363
rect 126756 2332 126897 2360
rect 126756 2320 126762 2332
rect 126885 2329 126897 2332
rect 126931 2329 126943 2363
rect 127636 2360 127664 2400
rect 130197 2397 130209 2400
rect 130243 2397 130255 2431
rect 133141 2431 133199 2437
rect 133141 2428 133153 2431
rect 130197 2391 130255 2397
rect 130304 2400 133153 2428
rect 130304 2360 130332 2400
rect 133141 2397 133153 2400
rect 133187 2428 133199 2431
rect 133693 2431 133751 2437
rect 133693 2428 133705 2431
rect 133187 2400 133705 2428
rect 133187 2397 133199 2400
rect 133141 2391 133199 2397
rect 133693 2397 133705 2400
rect 133739 2397 133751 2431
rect 135349 2431 135407 2437
rect 135349 2428 135361 2431
rect 133693 2391 133751 2397
rect 134996 2400 135361 2428
rect 127636 2332 130332 2360
rect 126885 2323 126943 2329
rect 130838 2320 130844 2372
rect 130896 2360 130902 2372
rect 131025 2363 131083 2369
rect 131025 2360 131037 2363
rect 130896 2332 131037 2360
rect 130896 2320 130902 2332
rect 131025 2329 131037 2332
rect 131071 2329 131083 2363
rect 131025 2323 131083 2329
rect 134996 2304 135024 2400
rect 135349 2397 135361 2400
rect 135395 2397 135407 2431
rect 135349 2391 135407 2397
rect 137278 2388 137284 2440
rect 137336 2428 137342 2440
rect 137925 2431 137983 2437
rect 137925 2428 137937 2431
rect 137336 2400 137937 2428
rect 137336 2388 137342 2400
rect 137925 2397 137937 2400
rect 137971 2397 137983 2431
rect 137925 2391 137983 2397
rect 138753 2431 138811 2437
rect 138753 2397 138765 2431
rect 138799 2428 138811 2431
rect 139118 2428 139124 2440
rect 138799 2400 139124 2428
rect 138799 2397 138811 2400
rect 138753 2391 138811 2397
rect 139118 2388 139124 2400
rect 139176 2428 139182 2440
rect 139213 2431 139271 2437
rect 139213 2428 139225 2431
rect 139176 2400 139225 2428
rect 139176 2388 139182 2400
rect 139213 2397 139225 2400
rect 139259 2397 139271 2431
rect 141973 2431 142031 2437
rect 141973 2428 141985 2431
rect 139213 2391 139271 2397
rect 141436 2400 141985 2428
rect 141436 2304 141464 2400
rect 141973 2397 141985 2400
rect 142019 2397 142031 2431
rect 141973 2391 142031 2397
rect 145926 2388 145932 2440
rect 145984 2428 145990 2440
rect 146113 2431 146171 2437
rect 146113 2428 146125 2431
rect 145984 2400 146125 2428
rect 145984 2388 145990 2400
rect 146113 2397 146125 2400
rect 146159 2397 146171 2431
rect 146113 2391 146171 2397
rect 143258 2320 143264 2372
rect 143316 2360 143322 2372
rect 143445 2363 143503 2369
rect 143445 2360 143457 2363
rect 143316 2332 143457 2360
rect 143316 2320 143322 2332
rect 143445 2329 143457 2332
rect 143491 2329 143503 2363
rect 143445 2323 143503 2329
rect 147398 2320 147404 2372
rect 147456 2360 147462 2372
rect 147585 2363 147643 2369
rect 147585 2360 147597 2363
rect 147456 2332 147597 2360
rect 147456 2320 147462 2332
rect 147585 2329 147597 2332
rect 147631 2360 147643 2363
rect 148229 2363 148287 2369
rect 148229 2360 148241 2363
rect 147631 2332 148241 2360
rect 147631 2329 147643 2332
rect 147585 2323 147643 2329
rect 148229 2329 148241 2332
rect 148275 2329 148287 2363
rect 148229 2323 148287 2329
rect 116670 2292 116676 2304
rect 114336 2264 114876 2292
rect 116631 2264 116676 2292
rect 114336 2252 114342 2264
rect 116670 2252 116676 2264
rect 116728 2252 116734 2304
rect 117038 2252 117044 2304
rect 117096 2292 117102 2304
rect 117501 2295 117559 2301
rect 117501 2292 117513 2295
rect 117096 2264 117513 2292
rect 117096 2252 117102 2264
rect 117501 2261 117513 2264
rect 117547 2261 117559 2295
rect 117501 2255 117559 2261
rect 121178 2252 121184 2304
rect 121236 2292 121242 2304
rect 121457 2295 121515 2301
rect 121457 2292 121469 2295
rect 121236 2264 121469 2292
rect 121236 2252 121242 2264
rect 121457 2261 121469 2264
rect 121503 2261 121515 2295
rect 121457 2255 121515 2261
rect 125318 2252 125324 2304
rect 125376 2292 125382 2304
rect 125597 2295 125655 2301
rect 125597 2292 125609 2295
rect 125376 2264 125609 2292
rect 125376 2252 125382 2264
rect 125597 2261 125609 2264
rect 125643 2261 125655 2295
rect 125597 2255 125655 2261
rect 129642 2252 129648 2304
rect 129700 2292 129706 2304
rect 130381 2295 130439 2301
rect 130381 2292 130393 2295
rect 129700 2264 130393 2292
rect 129700 2252 129706 2264
rect 130381 2261 130393 2264
rect 130427 2261 130439 2295
rect 130381 2255 130439 2261
rect 133598 2252 133604 2304
rect 133656 2292 133662 2304
rect 133877 2295 133935 2301
rect 133877 2292 133889 2295
rect 133656 2264 133889 2292
rect 133656 2252 133662 2264
rect 133877 2261 133889 2264
rect 133923 2261 133935 2295
rect 133877 2255 133935 2261
rect 134797 2295 134855 2301
rect 134797 2261 134809 2295
rect 134843 2292 134855 2295
rect 134978 2292 134984 2304
rect 134843 2264 134984 2292
rect 134843 2261 134855 2264
rect 134797 2255 134855 2261
rect 134978 2252 134984 2264
rect 135036 2252 135042 2304
rect 137738 2252 137744 2304
rect 137796 2292 137802 2304
rect 138109 2295 138167 2301
rect 138109 2292 138121 2295
rect 137796 2264 138121 2292
rect 137796 2252 137802 2264
rect 138109 2261 138121 2264
rect 138155 2261 138167 2295
rect 141418 2292 141424 2304
rect 141379 2264 141424 2292
rect 138109 2255 138167 2261
rect 141418 2252 141424 2264
rect 141476 2252 141482 2304
rect 141878 2252 141884 2304
rect 141936 2292 141942 2304
rect 142157 2295 142215 2301
rect 142157 2292 142169 2295
rect 141936 2264 142169 2292
rect 141936 2252 141942 2264
rect 142157 2261 142169 2264
rect 142203 2261 142215 2295
rect 142157 2255 142215 2261
rect 146018 2252 146024 2304
rect 146076 2292 146082 2304
rect 146297 2295 146355 2301
rect 146297 2292 146309 2295
rect 146076 2264 146309 2292
rect 146076 2252 146082 2264
rect 146297 2261 146309 2264
rect 146343 2261 146355 2295
rect 146297 2255 146355 2261
rect 1104 2202 148856 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 81014 2202
rect 81066 2150 81078 2202
rect 81130 2150 81142 2202
rect 81194 2150 81206 2202
rect 81258 2150 81270 2202
rect 81322 2150 111734 2202
rect 111786 2150 111798 2202
rect 111850 2150 111862 2202
rect 111914 2150 111926 2202
rect 111978 2150 111990 2202
rect 112042 2150 142454 2202
rect 142506 2150 142518 2202
rect 142570 2150 142582 2202
rect 142634 2150 142646 2202
rect 142698 2150 142710 2202
rect 142762 2150 148856 2202
rect 1104 2128 148856 2150
rect 8570 2048 8576 2100
rect 8628 2088 8634 2100
rect 23290 2088 23296 2100
rect 8628 2060 23296 2088
rect 8628 2048 8634 2060
rect 23290 2048 23296 2060
rect 23348 2048 23354 2100
rect 57422 2048 57428 2100
rect 57480 2088 57486 2100
rect 96062 2088 96068 2100
rect 57480 2060 96068 2088
rect 57480 2048 57486 2060
rect 96062 2048 96068 2060
rect 96120 2048 96126 2100
rect 56042 1980 56048 2032
rect 56100 2020 56106 2032
rect 91738 2020 91744 2032
rect 56100 1992 91744 2020
rect 56100 1980 56106 1992
rect 91738 1980 91744 1992
rect 91796 1980 91802 2032
rect 64874 1912 64880 1964
rect 64932 1952 64938 1964
rect 67542 1952 67548 1964
rect 64932 1924 67548 1952
rect 64932 1912 64938 1924
rect 67542 1912 67548 1924
rect 67600 1952 67606 1964
rect 100018 1952 100024 1964
rect 67600 1924 100024 1952
rect 67600 1912 67606 1924
rect 100018 1912 100024 1924
rect 100076 1912 100082 1964
rect 70946 1844 70952 1896
rect 71004 1884 71010 1896
rect 71682 1884 71688 1896
rect 71004 1856 71688 1884
rect 71004 1844 71010 1856
rect 71682 1844 71688 1856
rect 71740 1844 71746 1896
rect 81158 1844 81164 1896
rect 81216 1884 81222 1896
rect 83274 1884 83280 1896
rect 81216 1856 83280 1884
rect 81216 1844 81222 1856
rect 83274 1844 83280 1856
rect 83332 1844 83338 1896
rect 72694 1776 72700 1828
rect 72752 1816 72758 1828
rect 116670 1816 116676 1828
rect 72752 1788 116676 1816
rect 72752 1776 72758 1788
rect 116670 1776 116676 1788
rect 116728 1776 116734 1828
rect 71222 1708 71228 1760
rect 71280 1748 71286 1760
rect 109034 1748 109040 1760
rect 71280 1720 109040 1748
rect 71280 1708 71286 1720
rect 109034 1708 109040 1720
rect 109092 1708 109098 1760
rect 78122 1640 78128 1692
rect 78180 1680 78186 1692
rect 141418 1680 141424 1692
rect 78180 1652 141424 1680
rect 78180 1640 78186 1652
rect 141418 1640 141424 1652
rect 141476 1640 141482 1692
rect 59814 1572 59820 1624
rect 59872 1612 59878 1624
rect 87598 1612 87604 1624
rect 59872 1584 87604 1612
rect 59872 1572 59878 1584
rect 87598 1572 87604 1584
rect 87656 1572 87662 1624
rect 82998 1504 83004 1556
rect 83056 1544 83062 1556
rect 125410 1544 125416 1556
rect 83056 1516 125416 1544
rect 83056 1504 83062 1516
rect 125410 1504 125416 1516
rect 125468 1504 125474 1556
rect 81434 1436 81440 1488
rect 81492 1476 81498 1488
rect 112438 1476 112444 1488
rect 81492 1448 112444 1476
rect 81492 1436 81498 1448
rect 112438 1436 112444 1448
rect 112496 1436 112502 1488
<< via1 >>
rect 42616 39312 42668 39364
rect 73620 39312 73672 39364
rect 39396 39244 39448 39296
rect 68652 39244 68704 39296
rect 46296 39176 46348 39228
rect 84936 39244 84988 39296
rect 22192 39108 22244 39160
rect 83832 39176 83884 39228
rect 75184 39108 75236 39160
rect 85304 39108 85356 39160
rect 63500 39040 63552 39092
rect 118056 39040 118108 39092
rect 43996 38972 44048 39024
rect 82084 38972 82136 39024
rect 46940 38904 46992 38956
rect 89812 38904 89864 38956
rect 49792 38836 49844 38888
rect 93032 38836 93084 38888
rect 95056 38836 95108 38888
rect 123116 38836 123168 38888
rect 35532 38768 35584 38820
rect 94228 38768 94280 38820
rect 54944 38700 54996 38752
rect 105268 38700 105320 38752
rect 59912 38632 59964 38684
rect 113732 38632 113784 38684
rect 60096 38564 60148 38616
rect 117872 38564 117924 38616
rect 61292 38496 61344 38548
rect 120080 38496 120132 38548
rect 62856 38428 62908 38480
rect 122564 38428 122616 38480
rect 53196 38360 53248 38412
rect 112996 38360 113048 38412
rect 64696 38292 64748 38344
rect 126520 38292 126572 38344
rect 48044 38224 48096 38276
rect 111248 38224 111300 38276
rect 58532 38156 58584 38208
rect 121460 38156 121512 38208
rect 66536 38088 66588 38140
rect 130292 38088 130344 38140
rect 58716 38020 58768 38072
rect 125876 38020 125928 38072
rect 51172 37952 51224 38004
rect 97540 37952 97592 38004
rect 54300 37884 54352 37936
rect 101956 37884 102008 37936
rect 33600 37816 33652 37868
rect 75184 37816 75236 37868
rect 75920 37816 75972 37868
rect 79324 37816 79376 37868
rect 80244 37816 80296 37868
rect 83188 37816 83240 37868
rect 99472 37816 99524 37868
rect 124956 37816 125008 37868
rect 45376 37748 45428 37800
rect 62672 37748 62724 37800
rect 64420 37748 64472 37800
rect 116216 37748 116268 37800
rect 40040 37680 40092 37732
rect 67548 37680 67600 37732
rect 68376 37680 68428 37732
rect 120632 37680 120684 37732
rect 19432 37612 19484 37664
rect 25136 37612 25188 37664
rect 29092 37612 29144 37664
rect 31024 37612 31076 37664
rect 33416 37612 33468 37664
rect 53564 37612 53616 37664
rect 55220 37612 55272 37664
rect 56140 37612 56192 37664
rect 110236 37612 110288 37664
rect 119896 37612 119948 37664
rect 126428 37612 126480 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 65654 37510 65706 37562
rect 65718 37510 65770 37562
rect 65782 37510 65834 37562
rect 65846 37510 65898 37562
rect 65910 37510 65962 37562
rect 96374 37510 96426 37562
rect 96438 37510 96490 37562
rect 96502 37510 96554 37562
rect 96566 37510 96618 37562
rect 96630 37510 96682 37562
rect 127094 37510 127146 37562
rect 127158 37510 127210 37562
rect 127222 37510 127274 37562
rect 127286 37510 127338 37562
rect 127350 37510 127402 37562
rect 2780 37451 2832 37460
rect 2780 37417 2789 37451
rect 2789 37417 2823 37451
rect 2823 37417 2832 37451
rect 2780 37408 2832 37417
rect 4528 37340 4580 37392
rect 4896 37247 4948 37256
rect 4896 37213 4905 37247
rect 4905 37213 4939 37247
rect 4939 37213 4948 37247
rect 4896 37204 4948 37213
rect 4620 37068 4672 37120
rect 5540 37068 5592 37120
rect 6920 37204 6972 37256
rect 8208 37204 8260 37256
rect 8576 37247 8628 37256
rect 8576 37213 8585 37247
rect 8585 37213 8619 37247
rect 8619 37213 8628 37247
rect 8576 37204 8628 37213
rect 9772 37204 9824 37256
rect 10048 37204 10100 37256
rect 12256 37247 12308 37256
rect 12256 37213 12265 37247
rect 12265 37213 12299 37247
rect 12299 37213 12308 37247
rect 12256 37204 12308 37213
rect 13176 37247 13228 37256
rect 13176 37213 13185 37247
rect 13185 37213 13219 37247
rect 13219 37213 13228 37247
rect 13176 37204 13228 37213
rect 15936 37247 15988 37256
rect 15936 37213 15945 37247
rect 15945 37213 15979 37247
rect 15979 37213 15988 37247
rect 15936 37204 15988 37213
rect 17316 37204 17368 37256
rect 17408 37204 17460 37256
rect 19064 37204 19116 37256
rect 19708 37247 19760 37256
rect 19708 37213 19717 37247
rect 19717 37213 19751 37247
rect 19751 37213 19760 37247
rect 19708 37204 19760 37213
rect 20628 37204 20680 37256
rect 20720 37204 20772 37256
rect 22284 37204 22336 37256
rect 29092 37340 29144 37392
rect 29644 37340 29696 37392
rect 31024 37408 31076 37460
rect 45376 37451 45428 37460
rect 45376 37417 45385 37451
rect 45385 37417 45419 37451
rect 45419 37417 45428 37451
rect 45376 37408 45428 37417
rect 47860 37408 47912 37460
rect 51724 37408 51776 37460
rect 55220 37408 55272 37460
rect 57520 37408 57572 37460
rect 58164 37408 58216 37460
rect 62396 37408 62448 37460
rect 72332 37408 72384 37460
rect 58348 37340 58400 37392
rect 59820 37383 59872 37392
rect 59820 37349 59829 37383
rect 59829 37349 59863 37383
rect 59863 37349 59872 37383
rect 59820 37340 59872 37349
rect 61108 37340 61160 37392
rect 22468 37204 22520 37256
rect 23296 37247 23348 37256
rect 23296 37213 23305 37247
rect 23305 37213 23339 37247
rect 23339 37213 23348 37247
rect 23296 37204 23348 37213
rect 23388 37204 23440 37256
rect 25136 37272 25188 37324
rect 27988 37315 28040 37324
rect 24676 37204 24728 37256
rect 7288 37068 7340 37120
rect 8300 37068 8352 37120
rect 9128 37068 9180 37120
rect 10324 37111 10376 37120
rect 10324 37077 10333 37111
rect 10333 37077 10367 37111
rect 10367 37077 10376 37111
rect 10324 37068 10376 37077
rect 10968 37111 11020 37120
rect 10968 37077 10977 37111
rect 10977 37077 11011 37111
rect 11011 37077 11020 37111
rect 10968 37068 11020 37077
rect 11888 37068 11940 37120
rect 12808 37068 12860 37120
rect 14648 37068 14700 37120
rect 21548 37136 21600 37188
rect 15476 37068 15528 37120
rect 15568 37068 15620 37120
rect 16580 37068 16632 37120
rect 17776 37111 17828 37120
rect 17776 37077 17785 37111
rect 17785 37077 17819 37111
rect 17819 37077 17828 37111
rect 17776 37068 17828 37077
rect 18328 37068 18380 37120
rect 19340 37068 19392 37120
rect 20168 37068 20220 37120
rect 21364 37111 21416 37120
rect 21364 37077 21373 37111
rect 21373 37077 21407 37111
rect 21407 37077 21416 37111
rect 21364 37068 21416 37077
rect 22100 37068 22152 37120
rect 22928 37068 22980 37120
rect 23940 37136 23992 37188
rect 25872 37204 25924 37256
rect 25044 37136 25096 37188
rect 25504 37136 25556 37188
rect 25964 37136 26016 37188
rect 24032 37068 24084 37120
rect 25136 37111 25188 37120
rect 25136 37077 25145 37111
rect 25145 37077 25179 37111
rect 25179 37077 25188 37111
rect 25136 37068 25188 37077
rect 25320 37068 25372 37120
rect 27988 37281 27997 37315
rect 27997 37281 28031 37315
rect 28031 37281 28040 37315
rect 27988 37272 28040 37281
rect 30012 37315 30064 37324
rect 27344 37247 27396 37256
rect 26516 37111 26568 37120
rect 26516 37077 26525 37111
rect 26525 37077 26559 37111
rect 26559 37077 26568 37111
rect 26516 37068 26568 37077
rect 27344 37213 27353 37247
rect 27353 37213 27387 37247
rect 27387 37213 27396 37247
rect 27344 37204 27396 37213
rect 30012 37281 30021 37315
rect 30021 37281 30055 37315
rect 30055 37281 30064 37315
rect 30012 37272 30064 37281
rect 33600 37315 33652 37324
rect 33600 37281 33609 37315
rect 33609 37281 33643 37315
rect 33643 37281 33652 37315
rect 33600 37272 33652 37281
rect 37556 37272 37608 37324
rect 40868 37272 40920 37324
rect 46204 37315 46256 37324
rect 28724 37204 28776 37256
rect 28908 37204 28960 37256
rect 27252 37136 27304 37188
rect 31300 37204 31352 37256
rect 34336 37247 34388 37256
rect 28172 37111 28224 37120
rect 28172 37077 28181 37111
rect 28181 37077 28215 37111
rect 28215 37077 28224 37111
rect 28172 37068 28224 37077
rect 28632 37068 28684 37120
rect 29368 37136 29420 37188
rect 29828 37179 29880 37188
rect 29828 37145 29837 37179
rect 29837 37145 29871 37179
rect 29871 37145 29880 37179
rect 29828 37136 29880 37145
rect 30748 37136 30800 37188
rect 31760 37136 31812 37188
rect 31116 37068 31168 37120
rect 31208 37068 31260 37120
rect 31484 37068 31536 37120
rect 34336 37213 34345 37247
rect 34345 37213 34379 37247
rect 34379 37213 34388 37247
rect 34336 37204 34388 37213
rect 34704 37204 34756 37256
rect 39396 37247 39448 37256
rect 39396 37213 39405 37247
rect 39405 37213 39439 37247
rect 39439 37213 39448 37247
rect 39396 37204 39448 37213
rect 40040 37247 40092 37256
rect 40040 37213 40049 37247
rect 40049 37213 40083 37247
rect 40083 37213 40092 37247
rect 40040 37204 40092 37213
rect 40132 37204 40184 37256
rect 42708 37204 42760 37256
rect 42800 37204 42852 37256
rect 46204 37281 46213 37315
rect 46213 37281 46247 37315
rect 46247 37281 46256 37315
rect 46204 37272 46256 37281
rect 32956 37136 33008 37188
rect 33600 37136 33652 37188
rect 35532 37179 35584 37188
rect 35532 37145 35541 37179
rect 35541 37145 35575 37179
rect 35575 37145 35584 37179
rect 35532 37136 35584 37145
rect 35716 37136 35768 37188
rect 32496 37111 32548 37120
rect 32496 37077 32505 37111
rect 32505 37077 32539 37111
rect 32539 37077 32548 37111
rect 32496 37068 32548 37077
rect 34428 37068 34480 37120
rect 34796 37068 34848 37120
rect 36084 37068 36136 37120
rect 36544 37111 36596 37120
rect 36544 37077 36553 37111
rect 36553 37077 36587 37111
rect 36587 37077 36596 37111
rect 36544 37068 36596 37077
rect 36636 37111 36688 37120
rect 36636 37077 36645 37111
rect 36645 37077 36679 37111
rect 36679 37077 36688 37111
rect 36636 37068 36688 37077
rect 38200 37068 38252 37120
rect 38476 37068 38528 37120
rect 38660 37068 38712 37120
rect 40408 37068 40460 37120
rect 40592 37068 40644 37120
rect 41236 37111 41288 37120
rect 41236 37077 41245 37111
rect 41245 37077 41279 37111
rect 41279 37077 41288 37111
rect 41236 37068 41288 37077
rect 41512 37068 41564 37120
rect 43812 37136 43864 37188
rect 45376 37204 45428 37256
rect 45652 37136 45704 37188
rect 45836 37136 45888 37188
rect 46940 37247 46992 37256
rect 46940 37213 46949 37247
rect 46949 37213 46983 37247
rect 46983 37213 46992 37247
rect 47860 37272 47912 37324
rect 48136 37315 48188 37324
rect 48136 37281 48145 37315
rect 48145 37281 48179 37315
rect 48179 37281 48188 37315
rect 48136 37272 48188 37281
rect 51724 37315 51776 37324
rect 46940 37204 46992 37213
rect 43444 37068 43496 37120
rect 43720 37068 43772 37120
rect 48504 37204 48556 37256
rect 49792 37247 49844 37256
rect 49792 37213 49801 37247
rect 49801 37213 49835 37247
rect 49835 37213 49844 37247
rect 49792 37204 49844 37213
rect 51172 37247 51224 37256
rect 51172 37213 51181 37247
rect 51181 37213 51215 37247
rect 51215 37213 51224 37247
rect 51724 37281 51733 37315
rect 51733 37281 51767 37315
rect 51767 37281 51776 37315
rect 51724 37272 51776 37281
rect 58256 37272 58308 37324
rect 58624 37315 58676 37324
rect 58624 37281 58633 37315
rect 58633 37281 58667 37315
rect 58667 37281 58676 37315
rect 58624 37272 58676 37281
rect 61292 37315 61344 37324
rect 61292 37281 61301 37315
rect 61301 37281 61335 37315
rect 61335 37281 61344 37315
rect 61292 37272 61344 37281
rect 61384 37272 61436 37324
rect 65064 37340 65116 37392
rect 66260 37340 66312 37392
rect 67548 37383 67600 37392
rect 65156 37272 65208 37324
rect 65432 37272 65484 37324
rect 67548 37349 67557 37383
rect 67557 37349 67591 37383
rect 67591 37349 67600 37383
rect 67548 37340 67600 37349
rect 67824 37340 67876 37392
rect 79140 37340 79192 37392
rect 79324 37408 79376 37460
rect 81348 37408 81400 37460
rect 81624 37340 81676 37392
rect 70860 37272 70912 37324
rect 51172 37204 51224 37213
rect 54944 37247 54996 37256
rect 54944 37213 54953 37247
rect 54953 37213 54987 37247
rect 54987 37213 54996 37247
rect 54944 37204 54996 37213
rect 56140 37204 56192 37256
rect 56692 37204 56744 37256
rect 58348 37204 58400 37256
rect 53564 37136 53616 37188
rect 55588 37136 55640 37188
rect 55680 37136 55732 37188
rect 59820 37136 59872 37188
rect 47768 37068 47820 37120
rect 48964 37068 49016 37120
rect 49608 37111 49660 37120
rect 49608 37077 49617 37111
rect 49617 37077 49651 37111
rect 49651 37077 49660 37111
rect 49608 37068 49660 37077
rect 51448 37068 51500 37120
rect 51540 37068 51592 37120
rect 52368 37111 52420 37120
rect 52368 37077 52377 37111
rect 52377 37077 52411 37111
rect 52411 37077 52420 37111
rect 52368 37068 52420 37077
rect 53196 37111 53248 37120
rect 53196 37077 53205 37111
rect 53205 37077 53239 37111
rect 53239 37077 53248 37111
rect 53196 37068 53248 37077
rect 53656 37111 53708 37120
rect 53656 37077 53665 37111
rect 53665 37077 53699 37111
rect 53699 37077 53708 37111
rect 53656 37068 53708 37077
rect 55128 37068 55180 37120
rect 56508 37068 56560 37120
rect 56784 37111 56836 37120
rect 56784 37077 56793 37111
rect 56793 37077 56827 37111
rect 56827 37077 56836 37111
rect 56784 37068 56836 37077
rect 57152 37111 57204 37120
rect 57152 37077 57161 37111
rect 57161 37077 57195 37111
rect 57195 37077 57204 37111
rect 57152 37068 57204 37077
rect 57520 37068 57572 37120
rect 57980 37068 58032 37120
rect 58624 37068 58676 37120
rect 58716 37068 58768 37120
rect 60740 37068 60792 37120
rect 61016 37204 61068 37256
rect 61752 37204 61804 37256
rect 63500 37247 63552 37256
rect 63500 37213 63509 37247
rect 63509 37213 63543 37247
rect 63543 37213 63552 37247
rect 63500 37204 63552 37213
rect 64144 37204 64196 37256
rect 64788 37247 64840 37256
rect 64788 37213 64797 37247
rect 64797 37213 64831 37247
rect 64831 37213 64840 37247
rect 64788 37204 64840 37213
rect 64880 37204 64932 37256
rect 65524 37204 65576 37256
rect 62396 37179 62448 37188
rect 62396 37145 62405 37179
rect 62405 37145 62439 37179
rect 62439 37145 62448 37179
rect 62396 37136 62448 37145
rect 62580 37136 62632 37188
rect 66260 37179 66312 37188
rect 63592 37111 63644 37120
rect 63592 37077 63601 37111
rect 63601 37077 63635 37111
rect 63635 37077 63644 37111
rect 63592 37068 63644 37077
rect 64052 37068 64104 37120
rect 65984 37068 66036 37120
rect 66260 37145 66269 37179
rect 66269 37145 66303 37179
rect 66303 37145 66312 37179
rect 66260 37136 66312 37145
rect 67272 37204 67324 37256
rect 67732 37179 67784 37188
rect 66812 37111 66864 37120
rect 66812 37077 66831 37111
rect 66831 37077 66864 37111
rect 67732 37145 67741 37179
rect 67741 37145 67775 37179
rect 67775 37145 67784 37179
rect 67732 37136 67784 37145
rect 68560 37179 68612 37188
rect 68560 37145 68569 37179
rect 68569 37145 68603 37179
rect 68603 37145 68612 37179
rect 68560 37136 68612 37145
rect 70492 37204 70544 37256
rect 72516 37204 72568 37256
rect 74540 37204 74592 37256
rect 75828 37272 75880 37324
rect 76196 37272 76248 37324
rect 77024 37315 77076 37324
rect 77024 37281 77033 37315
rect 77033 37281 77067 37315
rect 77067 37281 77076 37315
rect 79508 37315 79560 37324
rect 77024 37272 77076 37281
rect 71136 37136 71188 37188
rect 71596 37136 71648 37188
rect 73620 37179 73672 37188
rect 73620 37145 73629 37179
rect 73629 37145 73663 37179
rect 73663 37145 73672 37179
rect 73620 37136 73672 37145
rect 73804 37179 73856 37188
rect 73804 37145 73813 37179
rect 73813 37145 73847 37179
rect 73847 37145 73856 37179
rect 73804 37136 73856 37145
rect 69020 37111 69072 37120
rect 66812 37068 66864 37077
rect 69020 37077 69039 37111
rect 69039 37077 69072 37111
rect 69020 37068 69072 37077
rect 69848 37068 69900 37120
rect 71320 37111 71372 37120
rect 71320 37077 71329 37111
rect 71329 37077 71363 37111
rect 71363 37077 71372 37111
rect 71320 37068 71372 37077
rect 71504 37068 71556 37120
rect 71780 37068 71832 37120
rect 73528 37068 73580 37120
rect 74724 37204 74776 37256
rect 75092 37136 75144 37188
rect 75552 37136 75604 37188
rect 77392 37204 77444 37256
rect 79508 37281 79517 37315
rect 79517 37281 79551 37315
rect 79551 37281 79560 37315
rect 79508 37272 79560 37281
rect 80796 37272 80848 37324
rect 81348 37272 81400 37324
rect 75736 37068 75788 37120
rect 76472 37111 76524 37120
rect 76472 37077 76505 37111
rect 76505 37077 76524 37111
rect 76472 37068 76524 37077
rect 77116 37068 77168 37120
rect 77300 37068 77352 37120
rect 79048 37111 79100 37120
rect 79048 37077 79057 37111
rect 79057 37077 79091 37111
rect 79091 37077 79100 37111
rect 79048 37068 79100 37077
rect 80428 37247 80480 37256
rect 80428 37213 80437 37247
rect 80437 37213 80471 37247
rect 80471 37213 80480 37247
rect 82728 37272 82780 37324
rect 89720 37408 89772 37460
rect 89812 37451 89864 37460
rect 89812 37417 89821 37451
rect 89821 37417 89855 37451
rect 89855 37417 89864 37451
rect 94228 37451 94280 37460
rect 89812 37408 89864 37417
rect 94228 37417 94237 37451
rect 94237 37417 94271 37451
rect 94271 37417 94280 37451
rect 94228 37408 94280 37417
rect 95056 37451 95108 37460
rect 95056 37417 95065 37451
rect 95065 37417 95099 37451
rect 95099 37417 95108 37451
rect 95056 37408 95108 37417
rect 97540 37451 97592 37460
rect 97540 37417 97549 37451
rect 97549 37417 97583 37451
rect 97583 37417 97592 37451
rect 97540 37408 97592 37417
rect 99472 37451 99524 37460
rect 99472 37417 99481 37451
rect 99481 37417 99515 37451
rect 99515 37417 99524 37451
rect 99472 37408 99524 37417
rect 101956 37451 102008 37460
rect 101956 37417 101965 37451
rect 101965 37417 101999 37451
rect 101999 37417 102008 37451
rect 101956 37408 102008 37417
rect 119896 37408 119948 37460
rect 120080 37451 120132 37460
rect 120080 37417 120089 37451
rect 120089 37417 120123 37451
rect 120123 37417 120132 37451
rect 120080 37408 120132 37417
rect 120448 37408 120500 37460
rect 122564 37451 122616 37460
rect 122564 37417 122573 37451
rect 122573 37417 122607 37451
rect 122607 37417 122616 37451
rect 122564 37408 122616 37417
rect 125876 37408 125928 37460
rect 83188 37340 83240 37392
rect 80428 37204 80480 37213
rect 82636 37204 82688 37256
rect 82820 37247 82872 37256
rect 82820 37213 82829 37247
rect 82829 37213 82863 37247
rect 82863 37213 82872 37247
rect 82820 37204 82872 37213
rect 83096 37272 83148 37324
rect 84200 37272 84252 37324
rect 89720 37272 89772 37324
rect 99472 37272 99524 37324
rect 102048 37272 102100 37324
rect 105912 37315 105964 37324
rect 105912 37281 105921 37315
rect 105921 37281 105955 37315
rect 105955 37281 105964 37315
rect 105912 37272 105964 37281
rect 110236 37272 110288 37324
rect 116216 37315 116268 37324
rect 116216 37281 116225 37315
rect 116225 37281 116259 37315
rect 116259 37281 116268 37315
rect 116216 37272 116268 37281
rect 118056 37315 118108 37324
rect 118056 37281 118065 37315
rect 118065 37281 118099 37315
rect 118099 37281 118108 37315
rect 118056 37272 118108 37281
rect 120632 37315 120684 37324
rect 120632 37281 120641 37315
rect 120641 37281 120675 37315
rect 120675 37281 120684 37315
rect 120632 37272 120684 37281
rect 123484 37272 123536 37324
rect 84844 37247 84896 37256
rect 84844 37213 84853 37247
rect 84853 37213 84887 37247
rect 84887 37213 84896 37247
rect 84844 37204 84896 37213
rect 85304 37247 85356 37256
rect 85304 37213 85313 37247
rect 85313 37213 85347 37247
rect 85347 37213 85356 37247
rect 85304 37204 85356 37213
rect 86776 37204 86828 37256
rect 86960 37204 87012 37256
rect 87512 37204 87564 37256
rect 88064 37204 88116 37256
rect 89628 37204 89680 37256
rect 90088 37204 90140 37256
rect 90732 37247 90784 37256
rect 90732 37213 90741 37247
rect 90741 37213 90775 37247
rect 90775 37213 90784 37247
rect 90732 37204 90784 37213
rect 91560 37247 91612 37256
rect 91560 37213 91569 37247
rect 91569 37213 91603 37247
rect 91603 37213 91612 37247
rect 91560 37204 91612 37213
rect 92112 37204 92164 37256
rect 92940 37204 92992 37256
rect 93860 37204 93912 37256
rect 96160 37204 96212 37256
rect 96712 37204 96764 37256
rect 98460 37247 98512 37256
rect 98460 37213 98469 37247
rect 98469 37213 98503 37247
rect 98503 37213 98512 37247
rect 98460 37204 98512 37213
rect 99288 37204 99340 37256
rect 99840 37204 99892 37256
rect 100576 37204 100628 37256
rect 81440 37136 81492 37188
rect 82268 37136 82320 37188
rect 83924 37179 83976 37188
rect 83924 37145 83933 37179
rect 83933 37145 83967 37179
rect 83967 37145 83976 37179
rect 83924 37136 83976 37145
rect 84568 37136 84620 37188
rect 80796 37068 80848 37120
rect 81808 37068 81860 37120
rect 82452 37111 82504 37120
rect 82452 37077 82461 37111
rect 82461 37077 82495 37111
rect 82495 37077 82504 37111
rect 82452 37068 82504 37077
rect 83096 37068 83148 37120
rect 84660 37111 84712 37120
rect 84660 37077 84669 37111
rect 84669 37077 84703 37111
rect 84703 37077 84712 37111
rect 84660 37068 84712 37077
rect 90364 37136 90416 37188
rect 97816 37136 97868 37188
rect 98736 37136 98788 37188
rect 99380 37179 99432 37188
rect 99380 37145 99389 37179
rect 99389 37145 99423 37179
rect 99423 37145 99432 37179
rect 99380 37136 99432 37145
rect 102784 37204 102836 37256
rect 102876 37247 102928 37256
rect 102876 37213 102885 37247
rect 102885 37213 102919 37247
rect 102919 37213 102928 37247
rect 104440 37247 104492 37256
rect 102876 37204 102928 37213
rect 104440 37213 104449 37247
rect 104449 37213 104483 37247
rect 104483 37213 104492 37247
rect 104440 37204 104492 37213
rect 104900 37204 104952 37256
rect 85580 37068 85632 37120
rect 87236 37111 87288 37120
rect 87236 37077 87245 37111
rect 87245 37077 87279 37111
rect 87279 37077 87288 37111
rect 87236 37068 87288 37077
rect 87328 37068 87380 37120
rect 88340 37068 88392 37120
rect 89260 37068 89312 37120
rect 91100 37068 91152 37120
rect 91928 37068 91980 37120
rect 92848 37068 92900 37120
rect 94320 37068 94372 37120
rect 95240 37068 95292 37120
rect 96804 37111 96856 37120
rect 96804 37077 96813 37111
rect 96813 37077 96847 37111
rect 96847 37077 96856 37111
rect 96804 37068 96856 37077
rect 98000 37068 98052 37120
rect 98552 37068 98604 37120
rect 102140 37136 102192 37188
rect 103428 37179 103480 37188
rect 103428 37145 103437 37179
rect 103437 37145 103471 37179
rect 103471 37145 103480 37179
rect 103428 37136 103480 37145
rect 100208 37111 100260 37120
rect 100208 37077 100217 37111
rect 100217 37077 100251 37111
rect 100251 37077 100260 37111
rect 100208 37068 100260 37077
rect 100760 37068 100812 37120
rect 102692 37111 102744 37120
rect 102692 37077 102701 37111
rect 102701 37077 102735 37111
rect 102735 37077 102744 37111
rect 102692 37068 102744 37077
rect 102784 37068 102836 37120
rect 106648 37204 106700 37256
rect 107292 37247 107344 37256
rect 107292 37213 107301 37247
rect 107301 37213 107335 37247
rect 107335 37213 107344 37247
rect 107292 37204 107344 37213
rect 107752 37247 107804 37256
rect 107752 37213 107761 37247
rect 107761 37213 107795 37247
rect 107795 37213 107804 37247
rect 107752 37204 107804 37213
rect 108488 37204 108540 37256
rect 109592 37247 109644 37256
rect 109592 37213 109601 37247
rect 109601 37213 109635 37247
rect 109635 37213 109644 37247
rect 109592 37204 109644 37213
rect 110696 37204 110748 37256
rect 112168 37247 112220 37256
rect 112168 37213 112177 37247
rect 112177 37213 112211 37247
rect 112211 37213 112220 37247
rect 112168 37204 112220 37213
rect 112260 37204 112312 37256
rect 112720 37204 112772 37256
rect 113456 37204 113508 37256
rect 114008 37204 114060 37256
rect 114836 37204 114888 37256
rect 115480 37247 115532 37256
rect 115480 37213 115489 37247
rect 115489 37213 115523 37247
rect 115523 37213 115532 37247
rect 115480 37204 115532 37213
rect 115940 37204 115992 37256
rect 116124 37204 116176 37256
rect 117136 37204 117188 37256
rect 103888 37068 103940 37120
rect 105360 37111 105412 37120
rect 105360 37077 105369 37111
rect 105369 37077 105403 37111
rect 105403 37077 105412 37111
rect 105360 37068 105412 37077
rect 106556 37068 106608 37120
rect 107108 37111 107160 37120
rect 107108 37077 107117 37111
rect 107117 37077 107151 37111
rect 107151 37077 107160 37111
rect 107108 37068 107160 37077
rect 107660 37068 107712 37120
rect 108764 37111 108816 37120
rect 108764 37077 108773 37111
rect 108773 37077 108807 37111
rect 108807 37077 108816 37111
rect 108764 37068 108816 37077
rect 109408 37068 109460 37120
rect 110420 37068 110472 37120
rect 117688 37136 117740 37188
rect 119160 37204 119212 37256
rect 119528 37204 119580 37256
rect 119896 37247 119948 37256
rect 119896 37213 119905 37247
rect 119905 37213 119939 37247
rect 119939 37213 119948 37247
rect 119896 37204 119948 37213
rect 120816 37179 120868 37188
rect 120816 37145 120825 37179
rect 120825 37145 120859 37179
rect 120859 37145 120868 37179
rect 120816 37136 120868 37145
rect 121736 37204 121788 37256
rect 122932 37204 122984 37256
rect 123116 37204 123168 37256
rect 123300 37204 123352 37256
rect 124404 37204 124456 37256
rect 124956 37204 125008 37256
rect 125140 37204 125192 37256
rect 125600 37204 125652 37256
rect 126428 37204 126480 37256
rect 126980 37204 127032 37256
rect 127716 37204 127768 37256
rect 128452 37204 128504 37256
rect 128728 37204 128780 37256
rect 129556 37204 129608 37256
rect 131120 37204 131172 37256
rect 131672 37247 131724 37256
rect 131672 37213 131681 37247
rect 131681 37213 131715 37247
rect 131715 37213 131724 37247
rect 131672 37204 131724 37213
rect 132500 37204 132552 37256
rect 133236 37204 133288 37256
rect 133512 37247 133564 37256
rect 133512 37213 133521 37247
rect 133521 37213 133555 37247
rect 133555 37213 133564 37247
rect 133512 37204 133564 37213
rect 134248 37204 134300 37256
rect 134432 37204 134484 37256
rect 135996 37204 136048 37256
rect 138020 37204 138072 37256
rect 138940 37247 138992 37256
rect 138940 37213 138949 37247
rect 138949 37213 138983 37247
rect 138983 37213 138992 37247
rect 138940 37204 138992 37213
rect 111248 37111 111300 37120
rect 111248 37077 111257 37111
rect 111257 37077 111291 37111
rect 111291 37077 111300 37111
rect 111248 37068 111300 37077
rect 111800 37068 111852 37120
rect 112996 37068 113048 37120
rect 113180 37068 113232 37120
rect 114560 37068 114612 37120
rect 115020 37068 115072 37120
rect 117320 37068 117372 37120
rect 118700 37068 118752 37120
rect 122840 37068 122892 37120
rect 124036 37111 124088 37120
rect 124036 37077 124045 37111
rect 124045 37077 124079 37111
rect 124079 37077 124088 37111
rect 124036 37068 124088 37077
rect 124220 37068 124272 37120
rect 126060 37068 126112 37120
rect 127808 37111 127860 37120
rect 127808 37077 127817 37111
rect 127817 37077 127851 37111
rect 127851 37077 127860 37111
rect 127808 37068 127860 37077
rect 128360 37068 128412 37120
rect 129280 37111 129332 37120
rect 129280 37077 129289 37111
rect 129289 37077 129323 37111
rect 129323 37077 129332 37111
rect 129280 37068 129332 37077
rect 129740 37068 129792 37120
rect 130476 37068 130528 37120
rect 131488 37068 131540 37120
rect 132868 37111 132920 37120
rect 132868 37077 132877 37111
rect 132877 37077 132911 37111
rect 132911 37077 132920 37111
rect 132868 37068 132920 37077
rect 133328 37068 133380 37120
rect 134524 37111 134576 37120
rect 134524 37077 134533 37111
rect 134533 37077 134567 37111
rect 134567 37077 134576 37111
rect 134524 37068 134576 37077
rect 135536 37111 135588 37120
rect 135536 37077 135545 37111
rect 135545 37077 135579 37111
rect 135579 37077 135588 37111
rect 135536 37068 135588 37077
rect 136088 37136 136140 37188
rect 137008 37068 137060 37120
rect 138848 37068 138900 37120
rect 139492 37068 139544 37120
rect 139768 37204 139820 37256
rect 140504 37247 140556 37256
rect 140504 37213 140513 37247
rect 140513 37213 140547 37247
rect 140547 37213 140556 37247
rect 140504 37204 140556 37213
rect 141608 37204 141660 37256
rect 142252 37247 142304 37256
rect 142252 37213 142261 37247
rect 142261 37213 142295 37247
rect 142295 37213 142304 37247
rect 142252 37204 142304 37213
rect 143080 37247 143132 37256
rect 143080 37213 143089 37247
rect 143089 37213 143123 37247
rect 143123 37213 143132 37247
rect 143080 37204 143132 37213
rect 143540 37204 143592 37256
rect 144552 37247 144604 37256
rect 144552 37213 144561 37247
rect 144561 37213 144595 37247
rect 144595 37213 144604 37247
rect 144552 37204 144604 37213
rect 145288 37204 145340 37256
rect 146300 37204 146352 37256
rect 147128 37204 147180 37256
rect 140688 37111 140740 37120
rect 140688 37077 140697 37111
rect 140697 37077 140731 37111
rect 140731 37077 140740 37111
rect 140688 37068 140740 37077
rect 140780 37068 140832 37120
rect 142160 37136 142212 37188
rect 142528 37068 142580 37120
rect 144000 37111 144052 37120
rect 144000 37077 144009 37111
rect 144009 37077 144043 37111
rect 144043 37077 144052 37111
rect 144000 37068 144052 37077
rect 144368 37068 144420 37120
rect 146208 37068 146260 37120
rect 147404 37111 147456 37120
rect 147404 37077 147413 37111
rect 147413 37077 147447 37111
rect 147447 37077 147456 37111
rect 147404 37068 147456 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 81014 36966 81066 37018
rect 81078 36966 81130 37018
rect 81142 36966 81194 37018
rect 81206 36966 81258 37018
rect 81270 36966 81322 37018
rect 111734 36966 111786 37018
rect 111798 36966 111850 37018
rect 111862 36966 111914 37018
rect 111926 36966 111978 37018
rect 111990 36966 112042 37018
rect 142454 36966 142506 37018
rect 142518 36966 142570 37018
rect 142582 36966 142634 37018
rect 142646 36966 142698 37018
rect 142710 36966 142762 37018
rect 3608 36864 3660 36916
rect 4528 36907 4580 36916
rect 4528 36873 4537 36907
rect 4537 36873 4571 36907
rect 4571 36873 4580 36907
rect 4528 36864 4580 36873
rect 8208 36907 8260 36916
rect 8208 36873 8217 36907
rect 8217 36873 8251 36907
rect 8251 36873 8260 36907
rect 8208 36864 8260 36873
rect 9772 36907 9824 36916
rect 9772 36873 9781 36907
rect 9781 36873 9815 36907
rect 9815 36873 9824 36907
rect 9772 36864 9824 36873
rect 12256 36864 12308 36916
rect 16580 36864 16632 36916
rect 17316 36907 17368 36916
rect 17316 36873 17325 36907
rect 17325 36873 17359 36907
rect 17359 36873 17368 36907
rect 17316 36864 17368 36873
rect 19064 36907 19116 36916
rect 19064 36873 19073 36907
rect 19073 36873 19107 36907
rect 19107 36873 19116 36907
rect 19064 36864 19116 36873
rect 19156 36864 19208 36916
rect 20444 36864 20496 36916
rect 20628 36907 20680 36916
rect 20628 36873 20637 36907
rect 20637 36873 20671 36907
rect 20671 36873 20680 36907
rect 20628 36864 20680 36873
rect 28356 36907 28408 36916
rect 28356 36873 28365 36907
rect 28365 36873 28399 36907
rect 28399 36873 28408 36907
rect 28356 36864 28408 36873
rect 28448 36864 28500 36916
rect 4896 36796 4948 36848
rect 6368 36728 6420 36780
rect 8392 36771 8444 36780
rect 8392 36737 8401 36771
rect 8401 36737 8435 36771
rect 8435 36737 8444 36771
rect 8392 36728 8444 36737
rect 10508 36728 10560 36780
rect 13176 36796 13228 36848
rect 21548 36796 21600 36848
rect 13820 36771 13872 36780
rect 13820 36737 13829 36771
rect 13829 36737 13863 36771
rect 13863 36737 13872 36771
rect 13820 36728 13872 36737
rect 17960 36728 18012 36780
rect 18052 36728 18104 36780
rect 19156 36728 19208 36780
rect 12900 36592 12952 36644
rect 18052 36592 18104 36644
rect 8392 36524 8444 36576
rect 9588 36524 9640 36576
rect 10508 36567 10560 36576
rect 10508 36533 10517 36567
rect 10517 36533 10551 36567
rect 10551 36533 10560 36567
rect 10508 36524 10560 36533
rect 15936 36524 15988 36576
rect 17684 36524 17736 36576
rect 17960 36567 18012 36576
rect 17960 36533 17969 36567
rect 17969 36533 18003 36567
rect 18003 36533 18012 36567
rect 17960 36524 18012 36533
rect 19524 36660 19576 36712
rect 20720 36728 20772 36780
rect 20168 36660 20220 36712
rect 21272 36728 21324 36780
rect 23940 36796 23992 36848
rect 24492 36839 24544 36848
rect 24492 36805 24501 36839
rect 24501 36805 24535 36839
rect 24535 36805 24544 36839
rect 24492 36796 24544 36805
rect 24676 36796 24728 36848
rect 21824 36728 21876 36780
rect 22744 36771 22796 36780
rect 22744 36737 22753 36771
rect 22753 36737 22787 36771
rect 22787 36737 22796 36771
rect 22744 36728 22796 36737
rect 23480 36728 23532 36780
rect 23848 36728 23900 36780
rect 24124 36728 24176 36780
rect 25320 36771 25372 36780
rect 21732 36660 21784 36712
rect 25044 36660 25096 36712
rect 25320 36737 25329 36771
rect 25329 36737 25363 36771
rect 25363 36737 25372 36771
rect 25320 36728 25372 36737
rect 25872 36796 25924 36848
rect 27252 36796 27304 36848
rect 27344 36796 27396 36848
rect 29828 36864 29880 36916
rect 30380 36864 30432 36916
rect 30564 36864 30616 36916
rect 33140 36864 33192 36916
rect 36452 36864 36504 36916
rect 36728 36907 36780 36916
rect 36728 36873 36737 36907
rect 36737 36873 36771 36907
rect 36771 36873 36780 36907
rect 36728 36864 36780 36873
rect 36820 36864 36872 36916
rect 28632 36728 28684 36780
rect 28816 36728 28868 36780
rect 29092 36771 29144 36780
rect 29092 36737 29101 36771
rect 29101 36737 29135 36771
rect 29135 36737 29144 36771
rect 29092 36728 29144 36737
rect 25964 36660 26016 36712
rect 27160 36592 27212 36644
rect 27252 36592 27304 36644
rect 28540 36660 28592 36712
rect 30656 36771 30708 36780
rect 30656 36737 30665 36771
rect 30665 36737 30699 36771
rect 30699 36737 30708 36771
rect 30656 36728 30708 36737
rect 31116 36771 31168 36780
rect 31116 36737 31125 36771
rect 31125 36737 31159 36771
rect 31159 36737 31168 36771
rect 31116 36728 31168 36737
rect 31484 36728 31536 36780
rect 33048 36728 33100 36780
rect 33140 36728 33192 36780
rect 33416 36771 33468 36780
rect 33416 36737 33425 36771
rect 33425 36737 33459 36771
rect 33459 36737 33468 36771
rect 33416 36728 33468 36737
rect 37280 36796 37332 36848
rect 38108 36796 38160 36848
rect 33968 36728 34020 36780
rect 34244 36728 34296 36780
rect 35992 36771 36044 36780
rect 35992 36737 36001 36771
rect 36001 36737 36035 36771
rect 36035 36737 36044 36771
rect 35992 36728 36044 36737
rect 36912 36771 36964 36780
rect 36912 36737 36914 36771
rect 36914 36737 36948 36771
rect 36948 36737 36964 36771
rect 36912 36728 36964 36737
rect 37096 36728 37148 36780
rect 40132 36796 40184 36848
rect 41604 36864 41656 36916
rect 42708 36864 42760 36916
rect 44088 36864 44140 36916
rect 44180 36864 44232 36916
rect 53012 36864 53064 36916
rect 53104 36864 53156 36916
rect 60648 36864 60700 36916
rect 64788 36864 64840 36916
rect 64880 36796 64932 36848
rect 38844 36771 38896 36780
rect 38844 36737 38853 36771
rect 38853 36737 38887 36771
rect 38887 36737 38896 36771
rect 38844 36728 38896 36737
rect 40224 36728 40276 36780
rect 40960 36728 41012 36780
rect 42800 36728 42852 36780
rect 43076 36703 43128 36712
rect 20260 36524 20312 36576
rect 20812 36524 20864 36576
rect 22192 36567 22244 36576
rect 22192 36533 22201 36567
rect 22201 36533 22235 36567
rect 22235 36533 22244 36567
rect 22192 36524 22244 36533
rect 23940 36524 23992 36576
rect 24676 36524 24728 36576
rect 24860 36524 24912 36576
rect 25964 36567 26016 36576
rect 25964 36533 25973 36567
rect 25973 36533 26007 36567
rect 26007 36533 26016 36567
rect 25964 36524 26016 36533
rect 26700 36524 26752 36576
rect 27344 36524 27396 36576
rect 27988 36592 28040 36644
rect 28632 36592 28684 36644
rect 28908 36592 28960 36644
rect 29644 36592 29696 36644
rect 33232 36524 33284 36576
rect 33600 36592 33652 36644
rect 35624 36592 35676 36644
rect 35716 36592 35768 36644
rect 40316 36592 40368 36644
rect 33784 36524 33836 36576
rect 34612 36524 34664 36576
rect 35348 36567 35400 36576
rect 35348 36533 35357 36567
rect 35357 36533 35391 36567
rect 35391 36533 35400 36567
rect 35348 36524 35400 36533
rect 37188 36524 37240 36576
rect 37556 36524 37608 36576
rect 39304 36524 39356 36576
rect 41052 36592 41104 36644
rect 41328 36635 41380 36644
rect 41328 36601 41337 36635
rect 41337 36601 41371 36635
rect 41371 36601 41380 36635
rect 41328 36592 41380 36601
rect 43076 36669 43085 36703
rect 43085 36669 43119 36703
rect 43119 36669 43128 36703
rect 43076 36660 43128 36669
rect 43996 36728 44048 36780
rect 44640 36771 44692 36780
rect 44640 36737 44649 36771
rect 44649 36737 44683 36771
rect 44683 36737 44692 36771
rect 44640 36728 44692 36737
rect 45008 36728 45060 36780
rect 46296 36771 46348 36780
rect 46296 36737 46305 36771
rect 46305 36737 46339 36771
rect 46339 36737 46348 36771
rect 46296 36728 46348 36737
rect 47216 36771 47268 36780
rect 47216 36737 47225 36771
rect 47225 36737 47259 36771
rect 47259 36737 47268 36771
rect 47216 36728 47268 36737
rect 47308 36728 47360 36780
rect 48596 36728 48648 36780
rect 50252 36771 50304 36780
rect 50252 36737 50261 36771
rect 50261 36737 50295 36771
rect 50295 36737 50304 36771
rect 50252 36728 50304 36737
rect 50896 36728 50948 36780
rect 51632 36771 51684 36780
rect 51632 36737 51641 36771
rect 51641 36737 51675 36771
rect 51675 36737 51684 36771
rect 51632 36728 51684 36737
rect 52092 36771 52144 36780
rect 52092 36737 52101 36771
rect 52101 36737 52135 36771
rect 52135 36737 52144 36771
rect 52092 36728 52144 36737
rect 44824 36635 44876 36644
rect 44824 36601 44833 36635
rect 44833 36601 44867 36635
rect 44867 36601 44876 36635
rect 44824 36592 44876 36601
rect 41972 36567 42024 36576
rect 41972 36533 41981 36567
rect 41981 36533 42015 36567
rect 42015 36533 42024 36567
rect 41972 36524 42024 36533
rect 42064 36524 42116 36576
rect 45836 36592 45888 36644
rect 45928 36592 45980 36644
rect 47860 36703 47912 36712
rect 47860 36669 47869 36703
rect 47869 36669 47903 36703
rect 47903 36669 47912 36703
rect 48044 36703 48096 36712
rect 47860 36660 47912 36669
rect 48044 36669 48053 36703
rect 48053 36669 48087 36703
rect 48087 36669 48096 36703
rect 48044 36660 48096 36669
rect 51816 36660 51868 36712
rect 53012 36728 53064 36780
rect 53932 36728 53984 36780
rect 55588 36771 55640 36780
rect 49516 36592 49568 36644
rect 54208 36660 54260 36712
rect 54760 36660 54812 36712
rect 55588 36737 55597 36771
rect 55597 36737 55631 36771
rect 55631 36737 55640 36771
rect 55588 36728 55640 36737
rect 56048 36728 56100 36780
rect 57336 36728 57388 36780
rect 57428 36728 57480 36780
rect 60096 36771 60148 36780
rect 56600 36660 56652 36712
rect 58256 36703 58308 36712
rect 58256 36669 58265 36703
rect 58265 36669 58299 36703
rect 58299 36669 58308 36703
rect 58256 36660 58308 36669
rect 58532 36660 58584 36712
rect 60096 36737 60105 36771
rect 60105 36737 60139 36771
rect 60139 36737 60148 36771
rect 60096 36728 60148 36737
rect 60740 36728 60792 36780
rect 61660 36771 61712 36780
rect 61660 36737 61669 36771
rect 61669 36737 61703 36771
rect 61703 36737 61712 36771
rect 61660 36728 61712 36737
rect 62120 36728 62172 36780
rect 63408 36728 63460 36780
rect 64236 36771 64288 36780
rect 64236 36737 64245 36771
rect 64245 36737 64279 36771
rect 64279 36737 64288 36771
rect 64236 36728 64288 36737
rect 64420 36728 64472 36780
rect 64604 36728 64656 36780
rect 66260 36864 66312 36916
rect 72792 36864 72844 36916
rect 74724 36864 74776 36916
rect 76288 36864 76340 36916
rect 77024 36864 77076 36916
rect 78680 36864 78732 36916
rect 80244 36864 80296 36916
rect 80336 36864 80388 36916
rect 119712 36864 119764 36916
rect 119896 36907 119948 36916
rect 119896 36873 119905 36907
rect 119905 36873 119939 36907
rect 119939 36873 119948 36907
rect 119896 36864 119948 36873
rect 119988 36864 120040 36916
rect 123576 36864 123628 36916
rect 124404 36907 124456 36916
rect 124404 36873 124413 36907
rect 124413 36873 124447 36907
rect 124447 36873 124456 36907
rect 124404 36864 124456 36873
rect 124956 36864 125008 36916
rect 125600 36907 125652 36916
rect 125600 36873 125609 36907
rect 125609 36873 125643 36907
rect 125643 36873 125652 36907
rect 125600 36864 125652 36873
rect 126520 36907 126572 36916
rect 126520 36873 126529 36907
rect 126529 36873 126563 36907
rect 126563 36873 126572 36907
rect 126520 36864 126572 36873
rect 127716 36907 127768 36916
rect 127716 36873 127725 36907
rect 127725 36873 127759 36907
rect 127759 36873 127768 36907
rect 127716 36864 127768 36873
rect 128360 36907 128412 36916
rect 128360 36873 128369 36907
rect 128369 36873 128403 36907
rect 128403 36873 128412 36907
rect 128360 36864 128412 36873
rect 128728 36864 128780 36916
rect 131120 36864 131172 36916
rect 133236 36907 133288 36916
rect 65340 36839 65392 36848
rect 65340 36805 65349 36839
rect 65349 36805 65383 36839
rect 65383 36805 65392 36839
rect 65340 36796 65392 36805
rect 65524 36796 65576 36848
rect 87236 36796 87288 36848
rect 87512 36839 87564 36848
rect 87512 36805 87521 36839
rect 87521 36805 87555 36839
rect 87555 36805 87564 36839
rect 87512 36796 87564 36805
rect 87604 36796 87656 36848
rect 66536 36771 66588 36780
rect 66536 36737 66545 36771
rect 66545 36737 66579 36771
rect 66579 36737 66588 36771
rect 66536 36728 66588 36737
rect 67088 36728 67140 36780
rect 68652 36771 68704 36780
rect 68652 36737 68661 36771
rect 68661 36737 68695 36771
rect 68695 36737 68704 36771
rect 68652 36728 68704 36737
rect 69204 36728 69256 36780
rect 69664 36771 69716 36780
rect 69664 36737 69673 36771
rect 69673 36737 69707 36771
rect 69707 36737 69716 36771
rect 69664 36728 69716 36737
rect 70768 36728 70820 36780
rect 72608 36728 72660 36780
rect 74540 36728 74592 36780
rect 75184 36728 75236 36780
rect 76196 36728 76248 36780
rect 76288 36728 76340 36780
rect 78956 36771 79008 36780
rect 78956 36737 78965 36771
rect 78965 36737 78999 36771
rect 78999 36737 79008 36771
rect 78956 36728 79008 36737
rect 79140 36728 79192 36780
rect 62396 36660 62448 36712
rect 63960 36660 64012 36712
rect 65064 36660 65116 36712
rect 53012 36635 53064 36644
rect 53012 36601 53021 36635
rect 53021 36601 53055 36635
rect 53055 36601 53064 36635
rect 53012 36592 53064 36601
rect 46756 36524 46808 36576
rect 47032 36567 47084 36576
rect 47032 36533 47041 36567
rect 47041 36533 47075 36567
rect 47075 36533 47084 36567
rect 47032 36524 47084 36533
rect 47124 36524 47176 36576
rect 47860 36524 47912 36576
rect 48044 36524 48096 36576
rect 48228 36524 48280 36576
rect 49148 36567 49200 36576
rect 49148 36533 49157 36567
rect 49157 36533 49191 36567
rect 49191 36533 49200 36567
rect 49148 36524 49200 36533
rect 51448 36567 51500 36576
rect 51448 36533 51457 36567
rect 51457 36533 51491 36567
rect 51491 36533 51500 36567
rect 51448 36524 51500 36533
rect 51816 36524 51868 36576
rect 64972 36592 65024 36644
rect 65800 36660 65852 36712
rect 75460 36660 75512 36712
rect 76656 36660 76708 36712
rect 80520 36728 80572 36780
rect 80612 36728 80664 36780
rect 82084 36771 82136 36780
rect 82084 36737 82093 36771
rect 82093 36737 82127 36771
rect 82127 36737 82136 36771
rect 82084 36728 82136 36737
rect 82268 36771 82320 36780
rect 82268 36737 82277 36771
rect 82277 36737 82311 36771
rect 82311 36737 82320 36771
rect 82268 36728 82320 36737
rect 83188 36728 83240 36780
rect 83740 36728 83792 36780
rect 83832 36771 83884 36780
rect 83832 36737 83841 36771
rect 83841 36737 83875 36771
rect 83875 36737 83884 36771
rect 84936 36771 84988 36780
rect 83832 36728 83884 36737
rect 84936 36737 84945 36771
rect 84945 36737 84979 36771
rect 84979 36737 84988 36771
rect 84936 36728 84988 36737
rect 85488 36728 85540 36780
rect 89076 36728 89128 36780
rect 90364 36771 90416 36780
rect 90364 36737 90373 36771
rect 90373 36737 90407 36771
rect 90407 36737 90416 36771
rect 90364 36728 90416 36737
rect 93032 36771 93084 36780
rect 93032 36737 93041 36771
rect 93041 36737 93075 36771
rect 93075 36737 93084 36771
rect 93032 36728 93084 36737
rect 94320 36728 94372 36780
rect 95240 36771 95292 36780
rect 95240 36737 95249 36771
rect 95249 36737 95283 36771
rect 95283 36737 95292 36771
rect 95240 36728 95292 36737
rect 95884 36728 95936 36780
rect 96712 36796 96764 36848
rect 98552 36796 98604 36848
rect 98736 36796 98788 36848
rect 99380 36839 99432 36848
rect 99380 36805 99389 36839
rect 99389 36805 99423 36839
rect 99423 36805 99432 36839
rect 99380 36796 99432 36805
rect 99840 36839 99892 36848
rect 99840 36805 99849 36839
rect 99849 36805 99883 36839
rect 99883 36805 99892 36839
rect 99840 36796 99892 36805
rect 102876 36796 102928 36848
rect 105268 36796 105320 36848
rect 106464 36796 106516 36848
rect 98000 36728 98052 36780
rect 100760 36728 100812 36780
rect 103060 36771 103112 36780
rect 103060 36737 103069 36771
rect 103069 36737 103103 36771
rect 103103 36737 103112 36771
rect 103060 36728 103112 36737
rect 106372 36771 106424 36780
rect 106372 36737 106381 36771
rect 106381 36737 106415 36771
rect 106415 36737 106424 36771
rect 106372 36728 106424 36737
rect 107292 36796 107344 36848
rect 108488 36796 108540 36848
rect 107568 36728 107620 36780
rect 112536 36796 112588 36848
rect 110512 36728 110564 36780
rect 112076 36728 112128 36780
rect 113732 36771 113784 36780
rect 113732 36737 113741 36771
rect 113741 36737 113775 36771
rect 113775 36737 113784 36771
rect 113732 36728 113784 36737
rect 114652 36728 114704 36780
rect 80796 36660 80848 36712
rect 81900 36660 81952 36712
rect 84844 36660 84896 36712
rect 85764 36660 85816 36712
rect 108304 36660 108356 36712
rect 116124 36796 116176 36848
rect 116308 36796 116360 36848
rect 116032 36728 116084 36780
rect 117136 36771 117188 36780
rect 117136 36737 117145 36771
rect 117145 36737 117179 36771
rect 117179 36737 117188 36771
rect 117136 36728 117188 36737
rect 117872 36771 117924 36780
rect 117872 36737 117881 36771
rect 117881 36737 117915 36771
rect 117915 36737 117924 36771
rect 117872 36728 117924 36737
rect 118700 36771 118752 36780
rect 118700 36737 118709 36771
rect 118709 36737 118743 36771
rect 118743 36737 118752 36771
rect 118700 36728 118752 36737
rect 119988 36728 120040 36780
rect 121368 36728 121420 36780
rect 122840 36728 122892 36780
rect 126980 36728 127032 36780
rect 129556 36771 129608 36780
rect 129556 36737 129565 36771
rect 129565 36737 129599 36771
rect 129599 36737 129608 36771
rect 129556 36728 129608 36737
rect 130936 36728 130988 36780
rect 132132 36796 132184 36848
rect 133236 36873 133245 36907
rect 133245 36873 133279 36907
rect 133279 36873 133288 36907
rect 133236 36864 133288 36873
rect 134248 36907 134300 36916
rect 134248 36873 134257 36907
rect 134257 36873 134291 36907
rect 134291 36873 134300 36907
rect 134248 36864 134300 36873
rect 135996 36907 136048 36916
rect 135996 36873 136005 36907
rect 136005 36873 136039 36907
rect 136039 36873 136048 36907
rect 135996 36864 136048 36873
rect 138940 36864 138992 36916
rect 140504 36907 140556 36916
rect 140504 36873 140513 36907
rect 140513 36873 140547 36907
rect 140547 36873 140556 36907
rect 140504 36864 140556 36873
rect 143080 36864 143132 36916
rect 144552 36864 144604 36916
rect 145288 36864 145340 36916
rect 146300 36907 146352 36916
rect 146300 36873 146309 36907
rect 146309 36873 146343 36907
rect 146343 36873 146352 36907
rect 146300 36864 146352 36873
rect 147128 36864 147180 36916
rect 133512 36796 133564 36848
rect 137284 36796 137336 36848
rect 142160 36796 142212 36848
rect 142252 36796 142304 36848
rect 132040 36771 132092 36780
rect 132040 36737 132049 36771
rect 132049 36737 132083 36771
rect 132083 36737 132092 36771
rect 132040 36728 132092 36737
rect 53748 36524 53800 36576
rect 54392 36567 54444 36576
rect 54392 36533 54401 36567
rect 54401 36533 54435 36567
rect 54435 36533 54444 36567
rect 54392 36524 54444 36533
rect 55128 36567 55180 36576
rect 55128 36533 55137 36567
rect 55137 36533 55171 36567
rect 55171 36533 55180 36567
rect 55128 36524 55180 36533
rect 56692 36524 56744 36576
rect 57060 36567 57112 36576
rect 57060 36533 57069 36567
rect 57069 36533 57103 36567
rect 57103 36533 57112 36567
rect 57060 36524 57112 36533
rect 59084 36524 59136 36576
rect 61016 36567 61068 36576
rect 61016 36533 61025 36567
rect 61025 36533 61059 36567
rect 61059 36533 61068 36567
rect 61016 36524 61068 36533
rect 63316 36524 63368 36576
rect 63500 36524 63552 36576
rect 63960 36524 64012 36576
rect 64788 36524 64840 36576
rect 64880 36524 64932 36576
rect 71320 36592 71372 36644
rect 73804 36592 73856 36644
rect 74632 36592 74684 36644
rect 75276 36592 75328 36644
rect 76564 36592 76616 36644
rect 65708 36524 65760 36576
rect 66260 36524 66312 36576
rect 70860 36524 70912 36576
rect 71044 36567 71096 36576
rect 71044 36533 71053 36567
rect 71053 36533 71087 36567
rect 71087 36533 71096 36567
rect 71044 36524 71096 36533
rect 71688 36567 71740 36576
rect 71688 36533 71697 36567
rect 71697 36533 71731 36567
rect 71731 36533 71740 36567
rect 71688 36524 71740 36533
rect 73988 36524 74040 36576
rect 76104 36524 76156 36576
rect 77300 36524 77352 36576
rect 77760 36567 77812 36576
rect 77760 36533 77769 36567
rect 77769 36533 77803 36567
rect 77803 36533 77812 36567
rect 77760 36524 77812 36533
rect 79784 36524 79836 36576
rect 123300 36660 123352 36712
rect 134432 36660 134484 36712
rect 82084 36524 82136 36576
rect 82268 36524 82320 36576
rect 83648 36524 83700 36576
rect 86408 36567 86460 36576
rect 86408 36533 86417 36567
rect 86417 36533 86451 36567
rect 86451 36533 86460 36567
rect 86408 36524 86460 36533
rect 86868 36524 86920 36576
rect 88064 36567 88116 36576
rect 88064 36533 88073 36567
rect 88073 36533 88107 36567
rect 88107 36533 88116 36567
rect 88064 36524 88116 36533
rect 89168 36524 89220 36576
rect 90456 36567 90508 36576
rect 90456 36533 90465 36567
rect 90465 36533 90499 36567
rect 90499 36533 90508 36567
rect 90456 36524 90508 36533
rect 91560 36567 91612 36576
rect 91560 36533 91569 36567
rect 91569 36533 91603 36567
rect 91603 36533 91612 36567
rect 91560 36524 91612 36533
rect 92112 36567 92164 36576
rect 92112 36533 92121 36567
rect 92121 36533 92155 36567
rect 92155 36533 92164 36567
rect 92112 36524 92164 36533
rect 94320 36524 94372 36576
rect 95056 36567 95108 36576
rect 95056 36533 95065 36567
rect 95065 36533 95099 36567
rect 95099 36533 95108 36567
rect 95056 36524 95108 36533
rect 95608 36524 95660 36576
rect 96160 36524 96212 36576
rect 98000 36567 98052 36576
rect 98000 36533 98009 36567
rect 98009 36533 98043 36567
rect 98043 36533 98052 36567
rect 98000 36524 98052 36533
rect 98644 36567 98696 36576
rect 98644 36533 98653 36567
rect 98653 36533 98687 36567
rect 98687 36533 98696 36567
rect 98644 36524 98696 36533
rect 100760 36567 100812 36576
rect 100760 36533 100769 36567
rect 100769 36533 100803 36567
rect 100803 36533 100812 36567
rect 100760 36524 100812 36533
rect 101128 36524 101180 36576
rect 102140 36524 102192 36576
rect 102968 36524 103020 36576
rect 104440 36567 104492 36576
rect 104440 36533 104449 36567
rect 104449 36533 104483 36567
rect 104483 36533 104492 36567
rect 104440 36524 104492 36533
rect 105728 36524 105780 36576
rect 109408 36524 109460 36576
rect 109592 36567 109644 36576
rect 109592 36533 109601 36567
rect 109601 36533 109635 36567
rect 109635 36533 109644 36567
rect 109592 36524 109644 36533
rect 110512 36524 110564 36576
rect 111892 36524 111944 36576
rect 116952 36524 117004 36576
rect 119160 36567 119212 36576
rect 119160 36533 119169 36567
rect 119169 36533 119203 36567
rect 119203 36533 119212 36567
rect 119160 36524 119212 36533
rect 121460 36524 121512 36576
rect 122840 36524 122892 36576
rect 127808 36592 127860 36644
rect 137652 36771 137704 36780
rect 137652 36737 137661 36771
rect 137661 36737 137695 36771
rect 137695 36737 137704 36771
rect 137652 36728 137704 36737
rect 143632 36771 143684 36780
rect 135904 36660 135956 36712
rect 141332 36660 141384 36712
rect 143632 36737 143641 36771
rect 143641 36737 143675 36771
rect 143675 36737 143684 36771
rect 143632 36728 143684 36737
rect 146300 36728 146352 36780
rect 123576 36524 123628 36576
rect 126520 36524 126572 36576
rect 126980 36524 127032 36576
rect 130292 36567 130344 36576
rect 130292 36533 130301 36567
rect 130301 36533 130335 36567
rect 130335 36533 130344 36567
rect 130292 36524 130344 36533
rect 130936 36567 130988 36576
rect 130936 36533 130945 36567
rect 130945 36533 130979 36567
rect 130979 36533 130988 36567
rect 130936 36524 130988 36533
rect 139492 36567 139544 36576
rect 139492 36533 139501 36567
rect 139501 36533 139535 36567
rect 139535 36533 139544 36567
rect 139492 36524 139544 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 65654 36422 65706 36474
rect 65718 36422 65770 36474
rect 65782 36422 65834 36474
rect 65846 36422 65898 36474
rect 65910 36422 65962 36474
rect 96374 36422 96426 36474
rect 96438 36422 96490 36474
rect 96502 36422 96554 36474
rect 96566 36422 96618 36474
rect 96630 36422 96682 36474
rect 127094 36422 127146 36474
rect 127158 36422 127210 36474
rect 127222 36422 127274 36474
rect 127286 36422 127338 36474
rect 127350 36422 127402 36474
rect 10048 36363 10100 36372
rect 10048 36329 10057 36363
rect 10057 36329 10091 36363
rect 10091 36329 10100 36363
rect 10048 36320 10100 36329
rect 17408 36363 17460 36372
rect 17408 36329 17417 36363
rect 17417 36329 17451 36363
rect 17451 36329 17460 36363
rect 17408 36320 17460 36329
rect 17776 36320 17828 36372
rect 22468 36363 22520 36372
rect 10508 36184 10560 36236
rect 14832 36184 14884 36236
rect 10324 36116 10376 36168
rect 21732 36252 21784 36304
rect 22468 36329 22477 36363
rect 22477 36329 22511 36363
rect 22511 36329 22520 36363
rect 22468 36320 22520 36329
rect 23480 36363 23532 36372
rect 23480 36329 23489 36363
rect 23489 36329 23523 36363
rect 23523 36329 23532 36363
rect 23480 36320 23532 36329
rect 24124 36320 24176 36372
rect 24860 36320 24912 36372
rect 25688 36320 25740 36372
rect 27620 36320 27672 36372
rect 29368 36320 29420 36372
rect 30656 36320 30708 36372
rect 32312 36320 32364 36372
rect 33692 36320 33744 36372
rect 33968 36320 34020 36372
rect 25136 36252 25188 36304
rect 25412 36252 25464 36304
rect 26332 36252 26384 36304
rect 36544 36320 36596 36372
rect 39304 36320 39356 36372
rect 39488 36363 39540 36372
rect 39488 36329 39497 36363
rect 39497 36329 39531 36363
rect 39531 36329 39540 36363
rect 39488 36320 39540 36329
rect 17960 36184 18012 36236
rect 15016 36116 15068 36168
rect 6920 36091 6972 36100
rect 6920 36057 6929 36091
rect 6929 36057 6963 36091
rect 6963 36057 6972 36091
rect 6920 36048 6972 36057
rect 14464 36048 14516 36100
rect 15108 36048 15160 36100
rect 15476 36116 15528 36168
rect 19524 36116 19576 36168
rect 20168 36159 20220 36168
rect 20168 36125 20177 36159
rect 20177 36125 20211 36159
rect 20211 36125 20220 36159
rect 20168 36116 20220 36125
rect 21088 36116 21140 36168
rect 21824 36159 21876 36168
rect 19432 36048 19484 36100
rect 20720 36048 20772 36100
rect 21824 36125 21833 36159
rect 21833 36125 21867 36159
rect 21867 36125 21876 36159
rect 21824 36116 21876 36125
rect 23940 36184 23992 36236
rect 34244 36295 34296 36304
rect 34244 36261 34253 36295
rect 34253 36261 34287 36295
rect 34287 36261 34296 36295
rect 34244 36252 34296 36261
rect 36360 36252 36412 36304
rect 37280 36295 37332 36304
rect 25136 36159 25188 36168
rect 25136 36125 25145 36159
rect 25145 36125 25179 36159
rect 25179 36125 25188 36159
rect 25136 36116 25188 36125
rect 34428 36184 34480 36236
rect 34612 36184 34664 36236
rect 37280 36261 37289 36295
rect 37289 36261 37323 36295
rect 37323 36261 37332 36295
rect 37280 36252 37332 36261
rect 42248 36320 42300 36372
rect 42892 36320 42944 36372
rect 36544 36184 36596 36236
rect 39948 36184 40000 36236
rect 26608 36116 26660 36168
rect 27896 36159 27948 36168
rect 27896 36125 27905 36159
rect 27905 36125 27939 36159
rect 27939 36125 27948 36159
rect 27896 36116 27948 36125
rect 8576 35980 8628 36032
rect 14740 35980 14792 36032
rect 14832 35980 14884 36032
rect 20536 35980 20588 36032
rect 21272 35980 21324 36032
rect 25412 36048 25464 36100
rect 26332 36048 26384 36100
rect 30840 36116 30892 36168
rect 32128 36116 32180 36168
rect 34704 36116 34756 36168
rect 35900 36159 35952 36168
rect 35900 36125 35909 36159
rect 35909 36125 35943 36159
rect 35943 36125 35952 36159
rect 35900 36116 35952 36125
rect 37280 36116 37332 36168
rect 37648 36116 37700 36168
rect 39488 36116 39540 36168
rect 41512 36184 41564 36236
rect 47308 36252 47360 36304
rect 41144 36116 41196 36168
rect 42616 36159 42668 36168
rect 42616 36125 42625 36159
rect 42625 36125 42659 36159
rect 42659 36125 42668 36159
rect 42616 36116 42668 36125
rect 44088 36159 44140 36168
rect 26792 35980 26844 36032
rect 28632 36023 28684 36032
rect 28632 35989 28641 36023
rect 28641 35989 28675 36023
rect 28675 35989 28684 36023
rect 28632 35980 28684 35989
rect 29276 35980 29328 36032
rect 32312 35980 32364 36032
rect 33140 36023 33192 36032
rect 33140 35989 33149 36023
rect 33149 35989 33183 36023
rect 33183 35989 33192 36023
rect 33140 35980 33192 35989
rect 33232 35980 33284 36032
rect 35992 35980 36044 36032
rect 36544 36023 36596 36032
rect 36544 35989 36553 36023
rect 36553 35989 36587 36023
rect 36587 35989 36596 36023
rect 36544 35980 36596 35989
rect 40040 35980 40092 36032
rect 41052 36048 41104 36100
rect 44088 36125 44097 36159
rect 44097 36125 44131 36159
rect 44131 36125 44140 36159
rect 44088 36116 44140 36125
rect 42064 35980 42116 36032
rect 44364 36048 44416 36100
rect 44640 36048 44692 36100
rect 47216 36184 47268 36236
rect 48596 36252 48648 36304
rect 51264 36252 51316 36304
rect 53012 36252 53064 36304
rect 53380 36320 53432 36372
rect 54300 36320 54352 36372
rect 54760 36363 54812 36372
rect 54760 36329 54769 36363
rect 54769 36329 54803 36363
rect 54803 36329 54812 36363
rect 54760 36320 54812 36329
rect 56048 36320 56100 36372
rect 56140 36320 56192 36372
rect 58716 36320 58768 36372
rect 58808 36320 58860 36372
rect 59820 36320 59872 36372
rect 61660 36320 61712 36372
rect 62488 36320 62540 36372
rect 64328 36320 64380 36372
rect 64788 36320 64840 36372
rect 66260 36320 66312 36372
rect 67088 36363 67140 36372
rect 67088 36329 67097 36363
rect 67097 36329 67131 36363
rect 67131 36329 67140 36363
rect 67088 36320 67140 36329
rect 68008 36320 68060 36372
rect 70400 36363 70452 36372
rect 70400 36329 70409 36363
rect 70409 36329 70443 36363
rect 70443 36329 70452 36363
rect 70400 36320 70452 36329
rect 55128 36252 55180 36304
rect 46848 36116 46900 36168
rect 48504 36116 48556 36168
rect 48688 36116 48740 36168
rect 48412 36048 48464 36100
rect 50620 36159 50672 36168
rect 50620 36125 50629 36159
rect 50629 36125 50663 36159
rect 50663 36125 50672 36159
rect 50620 36116 50672 36125
rect 52276 36116 52328 36168
rect 53104 36116 53156 36168
rect 54300 36116 54352 36168
rect 57980 36159 58032 36168
rect 49700 36048 49752 36100
rect 50252 36048 50304 36100
rect 52736 36091 52788 36100
rect 52736 36057 52745 36091
rect 52745 36057 52779 36091
rect 52779 36057 52788 36091
rect 52736 36048 52788 36057
rect 52920 36091 52972 36100
rect 52920 36057 52929 36091
rect 52929 36057 52963 36091
rect 52963 36057 52972 36091
rect 52920 36048 52972 36057
rect 44180 35980 44232 36032
rect 45284 36023 45336 36032
rect 45284 35989 45293 36023
rect 45293 35989 45327 36023
rect 45327 35989 45336 36023
rect 45284 35980 45336 35989
rect 50712 35980 50764 36032
rect 51540 36023 51592 36032
rect 51540 35989 51549 36023
rect 51549 35989 51583 36023
rect 51583 35989 51592 36023
rect 51540 35980 51592 35989
rect 53012 35980 53064 36032
rect 57152 36091 57204 36100
rect 57152 36057 57161 36091
rect 57161 36057 57195 36091
rect 57195 36057 57204 36091
rect 57152 36048 57204 36057
rect 57980 36125 57989 36159
rect 57989 36125 58023 36159
rect 58023 36125 58032 36159
rect 57980 36116 58032 36125
rect 58072 36048 58124 36100
rect 58900 36091 58952 36100
rect 58900 36057 58909 36091
rect 58909 36057 58943 36091
rect 58943 36057 58952 36091
rect 58900 36048 58952 36057
rect 59268 36048 59320 36100
rect 59728 36184 59780 36236
rect 62580 36252 62632 36304
rect 63316 36252 63368 36304
rect 67824 36252 67876 36304
rect 72332 36320 72384 36372
rect 72608 36363 72660 36372
rect 72608 36329 72617 36363
rect 72617 36329 72651 36363
rect 72651 36329 72660 36363
rect 72608 36320 72660 36329
rect 74448 36320 74500 36372
rect 75552 36320 75604 36372
rect 76288 36363 76340 36372
rect 76288 36329 76297 36363
rect 76297 36329 76331 36363
rect 76331 36329 76340 36363
rect 76288 36320 76340 36329
rect 70860 36252 70912 36304
rect 71136 36252 71188 36304
rect 79968 36320 80020 36372
rect 80152 36320 80204 36372
rect 80520 36320 80572 36372
rect 89260 36320 89312 36372
rect 90732 36363 90784 36372
rect 90732 36329 90741 36363
rect 90741 36329 90775 36363
rect 90775 36329 90784 36363
rect 90732 36320 90784 36329
rect 93860 36320 93912 36372
rect 102876 36320 102928 36372
rect 103060 36320 103112 36372
rect 103428 36363 103480 36372
rect 103428 36329 103437 36363
rect 103437 36329 103471 36363
rect 103471 36329 103480 36363
rect 103428 36320 103480 36329
rect 104900 36320 104952 36372
rect 106372 36363 106424 36372
rect 106372 36329 106381 36363
rect 106381 36329 106415 36363
rect 106415 36329 106424 36363
rect 106372 36320 106424 36329
rect 106556 36320 106608 36372
rect 107568 36320 107620 36372
rect 107752 36320 107804 36372
rect 110696 36320 110748 36372
rect 112352 36320 112404 36372
rect 115480 36320 115532 36372
rect 117688 36320 117740 36372
rect 119712 36320 119764 36372
rect 123208 36320 123260 36372
rect 123300 36320 123352 36372
rect 135904 36320 135956 36372
rect 136088 36363 136140 36372
rect 136088 36329 136097 36363
rect 136097 36329 136131 36363
rect 136131 36329 136140 36363
rect 136088 36320 136140 36329
rect 138020 36363 138072 36372
rect 138020 36329 138029 36363
rect 138029 36329 138063 36363
rect 138063 36329 138072 36363
rect 138020 36320 138072 36329
rect 143540 36320 143592 36372
rect 59912 36116 59964 36168
rect 64604 36184 64656 36236
rect 67732 36184 67784 36236
rect 60372 36116 60424 36168
rect 61384 36159 61436 36168
rect 61384 36125 61393 36159
rect 61393 36125 61427 36159
rect 61427 36125 61436 36159
rect 61384 36116 61436 36125
rect 62580 36116 62632 36168
rect 62856 36159 62908 36168
rect 62856 36125 62865 36159
rect 62865 36125 62899 36159
rect 62899 36125 62908 36159
rect 62856 36116 62908 36125
rect 64696 36159 64748 36168
rect 64696 36125 64705 36159
rect 64705 36125 64739 36159
rect 64739 36125 64748 36159
rect 64696 36116 64748 36125
rect 65340 36116 65392 36168
rect 68192 36116 68244 36168
rect 68376 36159 68428 36168
rect 68376 36125 68385 36159
rect 68385 36125 68419 36159
rect 68419 36125 68428 36159
rect 68376 36116 68428 36125
rect 68928 36116 68980 36168
rect 71044 36184 71096 36236
rect 80612 36184 80664 36236
rect 81348 36227 81400 36236
rect 81348 36193 81357 36227
rect 81357 36193 81391 36227
rect 81391 36193 81400 36227
rect 81348 36184 81400 36193
rect 61660 36048 61712 36100
rect 62028 36048 62080 36100
rect 63684 36091 63736 36100
rect 63684 36057 63693 36091
rect 63693 36057 63727 36091
rect 63727 36057 63736 36091
rect 63684 36048 63736 36057
rect 63868 36091 63920 36100
rect 63868 36057 63877 36091
rect 63877 36057 63911 36091
rect 63911 36057 63920 36091
rect 63868 36048 63920 36057
rect 56600 35980 56652 36032
rect 65432 36048 65484 36100
rect 66076 36091 66128 36100
rect 64788 35980 64840 36032
rect 66076 36057 66085 36091
rect 66085 36057 66119 36091
rect 66119 36057 66128 36091
rect 66076 36048 66128 36057
rect 66444 35980 66496 36032
rect 73988 36048 74040 36100
rect 74448 36116 74500 36168
rect 74632 36116 74684 36168
rect 76104 36159 76156 36168
rect 75092 36048 75144 36100
rect 76104 36125 76113 36159
rect 76113 36125 76147 36159
rect 76147 36125 76156 36159
rect 76104 36116 76156 36125
rect 77300 36159 77352 36168
rect 77300 36125 77309 36159
rect 77309 36125 77343 36159
rect 77343 36125 77352 36159
rect 77300 36116 77352 36125
rect 80060 36159 80112 36168
rect 80060 36125 80069 36159
rect 80069 36125 80103 36159
rect 80103 36125 80112 36159
rect 80060 36116 80112 36125
rect 80428 36116 80480 36168
rect 82820 36184 82872 36236
rect 83648 36184 83700 36236
rect 86408 36252 86460 36304
rect 119160 36252 119212 36304
rect 120816 36252 120868 36304
rect 126428 36295 126480 36304
rect 81624 36159 81676 36168
rect 81624 36125 81633 36159
rect 81633 36125 81667 36159
rect 81667 36125 81676 36159
rect 81624 36116 81676 36125
rect 81716 36116 81768 36168
rect 82360 36116 82412 36168
rect 87604 36116 87656 36168
rect 78496 36091 78548 36100
rect 78496 36057 78505 36091
rect 78505 36057 78539 36091
rect 78539 36057 78548 36091
rect 78496 36048 78548 36057
rect 95056 36116 95108 36168
rect 75184 36023 75236 36032
rect 75184 35989 75193 36023
rect 75193 35989 75227 36023
rect 75227 35989 75236 36023
rect 75184 35980 75236 35989
rect 75736 35980 75788 36032
rect 92388 36048 92440 36100
rect 99380 36116 99432 36168
rect 99472 36116 99524 36168
rect 105636 36116 105688 36168
rect 106464 36184 106516 36236
rect 108304 36184 108356 36236
rect 116308 36184 116360 36236
rect 120908 36184 120960 36236
rect 124220 36184 124272 36236
rect 126428 36261 126437 36295
rect 126437 36261 126471 36295
rect 126471 36261 126480 36295
rect 126428 36252 126480 36261
rect 126520 36252 126572 36304
rect 132040 36252 132092 36304
rect 132132 36252 132184 36304
rect 137284 36252 137336 36304
rect 139492 36184 139544 36236
rect 112352 36116 112404 36168
rect 112536 36116 112588 36168
rect 143632 36116 143684 36168
rect 95240 36048 95292 36100
rect 98460 36048 98512 36100
rect 98644 36048 98696 36100
rect 146300 36048 146352 36100
rect 147312 36048 147364 36100
rect 78956 35980 79008 36032
rect 79140 36023 79192 36032
rect 79140 35989 79149 36023
rect 79149 35989 79183 36023
rect 79183 35989 79192 36023
rect 79140 35980 79192 35989
rect 81716 35980 81768 36032
rect 81992 36023 82044 36032
rect 81992 35989 82001 36023
rect 82001 35989 82035 36023
rect 82035 35989 82044 36023
rect 81992 35980 82044 35989
rect 83096 36023 83148 36032
rect 83096 35989 83105 36023
rect 83105 35989 83139 36023
rect 83139 35989 83148 36023
rect 83096 35980 83148 35989
rect 83648 36023 83700 36032
rect 83648 35989 83657 36023
rect 83657 35989 83691 36023
rect 83691 35989 83700 36023
rect 83648 35980 83700 35989
rect 83740 35980 83792 36032
rect 84200 35980 84252 36032
rect 84752 36023 84804 36032
rect 84752 35989 84761 36023
rect 84761 35989 84795 36023
rect 84795 35989 84804 36023
rect 84752 35980 84804 35989
rect 85488 35980 85540 36032
rect 89076 36023 89128 36032
rect 89076 35989 89085 36023
rect 89085 35989 89119 36023
rect 89119 35989 89128 36023
rect 89076 35980 89128 35989
rect 89628 36023 89680 36032
rect 89628 35989 89637 36023
rect 89637 35989 89671 36023
rect 89671 35989 89680 36023
rect 89628 35980 89680 35989
rect 89720 35980 89772 36032
rect 90364 35980 90416 36032
rect 92848 36023 92900 36032
rect 92848 35989 92857 36023
rect 92857 35989 92891 36023
rect 92891 35989 92900 36023
rect 92848 35980 92900 35989
rect 94320 35980 94372 36032
rect 95884 36023 95936 36032
rect 95884 35989 95893 36023
rect 95893 35989 95927 36023
rect 95927 35989 95936 36023
rect 95884 35980 95936 35989
rect 97816 36023 97868 36032
rect 97816 35989 97825 36023
rect 97825 35989 97859 36023
rect 97859 35989 97868 36023
rect 97816 35980 97868 35989
rect 98368 36023 98420 36032
rect 98368 35989 98377 36023
rect 98377 35989 98411 36023
rect 98411 35989 98420 36023
rect 98368 35980 98420 35989
rect 99380 35980 99432 36032
rect 100576 36023 100628 36032
rect 100576 35989 100585 36023
rect 100585 35989 100619 36023
rect 100619 35989 100628 36023
rect 100576 35980 100628 35989
rect 105820 35980 105872 36032
rect 110236 35980 110288 36032
rect 112168 36023 112220 36032
rect 112168 35989 112177 36023
rect 112177 35989 112211 36023
rect 112211 35989 112220 36023
rect 112168 35980 112220 35989
rect 112720 36023 112772 36032
rect 112720 35989 112729 36023
rect 112729 35989 112763 36023
rect 112763 35989 112772 36023
rect 112720 35980 112772 35989
rect 113456 36023 113508 36032
rect 113456 35989 113465 36023
rect 113465 35989 113499 36023
rect 113499 35989 113508 36023
rect 113456 35980 113508 35989
rect 114652 35980 114704 36032
rect 114928 35980 114980 36032
rect 116952 35980 117004 36032
rect 120908 35980 120960 36032
rect 121552 36023 121604 36032
rect 121552 35989 121561 36023
rect 121561 35989 121595 36023
rect 121595 35989 121604 36023
rect 121552 35980 121604 35989
rect 123116 36023 123168 36032
rect 123116 35989 123125 36023
rect 123125 35989 123159 36023
rect 123159 35989 123168 36023
rect 123116 35980 123168 35989
rect 123208 35980 123260 36032
rect 130476 35980 130528 36032
rect 130936 35980 130988 36032
rect 137652 35980 137704 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 81014 35878 81066 35930
rect 81078 35878 81130 35930
rect 81142 35878 81194 35930
rect 81206 35878 81258 35930
rect 81270 35878 81322 35930
rect 111734 35878 111786 35930
rect 111798 35878 111850 35930
rect 111862 35878 111914 35930
rect 111926 35878 111978 35930
rect 111990 35878 112042 35930
rect 142454 35878 142506 35930
rect 142518 35878 142570 35930
rect 142582 35878 142634 35930
rect 142646 35878 142698 35930
rect 142710 35878 142762 35930
rect 19984 35776 20036 35828
rect 21088 35819 21140 35828
rect 21088 35785 21097 35819
rect 21097 35785 21131 35819
rect 21131 35785 21140 35819
rect 21088 35776 21140 35785
rect 25136 35776 25188 35828
rect 26608 35819 26660 35828
rect 26608 35785 26617 35819
rect 26617 35785 26651 35819
rect 26651 35785 26660 35819
rect 26608 35776 26660 35785
rect 28540 35819 28592 35828
rect 28540 35785 28549 35819
rect 28549 35785 28583 35819
rect 28583 35785 28592 35819
rect 28540 35776 28592 35785
rect 28632 35776 28684 35828
rect 29276 35776 29328 35828
rect 31944 35776 31996 35828
rect 37464 35776 37516 35828
rect 37648 35819 37700 35828
rect 37648 35785 37657 35819
rect 37657 35785 37691 35819
rect 37691 35785 37700 35819
rect 37648 35776 37700 35785
rect 38660 35819 38712 35828
rect 38660 35785 38669 35819
rect 38669 35785 38703 35819
rect 38703 35785 38712 35819
rect 38660 35776 38712 35785
rect 39396 35776 39448 35828
rect 41236 35776 41288 35828
rect 42524 35776 42576 35828
rect 42616 35776 42668 35828
rect 43168 35776 43220 35828
rect 44088 35776 44140 35828
rect 45008 35776 45060 35828
rect 46296 35776 46348 35828
rect 46940 35776 46992 35828
rect 48688 35776 48740 35828
rect 50620 35776 50672 35828
rect 51724 35776 51776 35828
rect 52276 35819 52328 35828
rect 52276 35785 52285 35819
rect 52285 35785 52319 35819
rect 52319 35785 52328 35819
rect 52276 35776 52328 35785
rect 54944 35776 54996 35828
rect 57980 35776 58032 35828
rect 58624 35776 58676 35828
rect 60096 35776 60148 35828
rect 60372 35819 60424 35828
rect 60372 35785 60381 35819
rect 60381 35785 60415 35819
rect 60415 35785 60424 35819
rect 60372 35776 60424 35785
rect 61292 35776 61344 35828
rect 63408 35776 63460 35828
rect 64420 35776 64472 35828
rect 64696 35776 64748 35828
rect 66536 35776 66588 35828
rect 67272 35819 67324 35828
rect 67272 35785 67281 35819
rect 67281 35785 67315 35819
rect 67315 35785 67324 35819
rect 67272 35776 67324 35785
rect 68376 35776 68428 35828
rect 80888 35776 80940 35828
rect 81348 35776 81400 35828
rect 82360 35819 82412 35828
rect 82360 35785 82369 35819
rect 82369 35785 82403 35819
rect 82403 35785 82412 35819
rect 82360 35776 82412 35785
rect 83832 35819 83884 35828
rect 83832 35785 83841 35819
rect 83841 35785 83875 35819
rect 83875 35785 83884 35819
rect 83832 35776 83884 35785
rect 85304 35776 85356 35828
rect 26792 35708 26844 35760
rect 28908 35708 28960 35760
rect 9588 35640 9640 35692
rect 34244 35708 34296 35760
rect 34336 35708 34388 35760
rect 32956 35640 33008 35692
rect 41236 35640 41288 35692
rect 46756 35708 46808 35760
rect 63592 35708 63644 35760
rect 70492 35708 70544 35760
rect 112076 35708 112128 35760
rect 57428 35640 57480 35692
rect 63868 35640 63920 35692
rect 64788 35640 64840 35692
rect 65248 35640 65300 35692
rect 80428 35683 80480 35692
rect 80428 35649 80437 35683
rect 80437 35649 80471 35683
rect 80471 35649 80480 35683
rect 80428 35640 80480 35649
rect 81900 35640 81952 35692
rect 83096 35640 83148 35692
rect 25136 35572 25188 35624
rect 41144 35572 41196 35624
rect 41420 35572 41472 35624
rect 48412 35572 48464 35624
rect 79508 35572 79560 35624
rect 81348 35572 81400 35624
rect 83648 35572 83700 35624
rect 123484 35572 123536 35624
rect 27896 35504 27948 35556
rect 24584 35436 24636 35488
rect 24860 35436 24912 35488
rect 30840 35436 30892 35488
rect 31300 35504 31352 35556
rect 31944 35504 31996 35556
rect 34704 35504 34756 35556
rect 35808 35547 35860 35556
rect 35808 35513 35817 35547
rect 35817 35513 35851 35547
rect 35851 35513 35860 35547
rect 35808 35504 35860 35513
rect 42524 35504 42576 35556
rect 52092 35504 52144 35556
rect 32956 35436 33008 35488
rect 33140 35479 33192 35488
rect 33140 35445 33149 35479
rect 33149 35445 33183 35479
rect 33183 35445 33192 35479
rect 33140 35436 33192 35445
rect 37280 35436 37332 35488
rect 38108 35479 38160 35488
rect 38108 35445 38117 35479
rect 38117 35445 38151 35479
rect 38151 35445 38160 35479
rect 38108 35436 38160 35445
rect 40224 35436 40276 35488
rect 40960 35436 41012 35488
rect 42800 35436 42852 35488
rect 44364 35436 44416 35488
rect 47124 35479 47176 35488
rect 47124 35445 47133 35479
rect 47133 35445 47167 35479
rect 47167 35445 47176 35479
rect 47124 35436 47176 35445
rect 48136 35479 48188 35488
rect 48136 35445 48145 35479
rect 48145 35445 48179 35479
rect 48179 35445 48188 35479
rect 48136 35436 48188 35445
rect 48596 35479 48648 35488
rect 48596 35445 48605 35479
rect 48605 35445 48639 35479
rect 48639 35445 48648 35479
rect 48596 35436 48648 35445
rect 49700 35436 49752 35488
rect 51632 35436 51684 35488
rect 52736 35436 52788 35488
rect 53104 35479 53156 35488
rect 53104 35445 53113 35479
rect 53113 35445 53147 35479
rect 53147 35445 53156 35479
rect 53104 35436 53156 35445
rect 53932 35436 53984 35488
rect 56600 35436 56652 35488
rect 57336 35436 57388 35488
rect 58900 35436 58952 35488
rect 81440 35504 81492 35556
rect 90456 35504 90508 35556
rect 121552 35504 121604 35556
rect 60740 35436 60792 35488
rect 62028 35436 62080 35488
rect 69204 35479 69256 35488
rect 69204 35445 69213 35479
rect 69213 35445 69247 35479
rect 69247 35445 69256 35479
rect 69204 35436 69256 35445
rect 75092 35479 75144 35488
rect 75092 35445 75101 35479
rect 75101 35445 75135 35479
rect 75135 35445 75144 35479
rect 75092 35436 75144 35445
rect 80060 35436 80112 35488
rect 82912 35479 82964 35488
rect 82912 35445 82921 35479
rect 82921 35445 82955 35479
rect 82955 35445 82964 35479
rect 82912 35436 82964 35445
rect 83924 35436 83976 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 65654 35334 65706 35386
rect 65718 35334 65770 35386
rect 65782 35334 65834 35386
rect 65846 35334 65898 35386
rect 65910 35334 65962 35386
rect 96374 35334 96426 35386
rect 96438 35334 96490 35386
rect 96502 35334 96554 35386
rect 96566 35334 96618 35386
rect 96630 35334 96682 35386
rect 127094 35334 127146 35386
rect 127158 35334 127210 35386
rect 127222 35334 127274 35386
rect 127286 35334 127338 35386
rect 127350 35334 127402 35386
rect 19984 35232 20036 35284
rect 20536 35232 20588 35284
rect 24492 35232 24544 35284
rect 24860 35232 24912 35284
rect 25504 35232 25556 35284
rect 28724 35275 28776 35284
rect 28724 35241 28733 35275
rect 28733 35241 28767 35275
rect 28767 35241 28776 35275
rect 28724 35232 28776 35241
rect 25228 35164 25280 35216
rect 75920 35232 75972 35284
rect 79508 35275 79560 35284
rect 79508 35241 79517 35275
rect 79517 35241 79551 35275
rect 79551 35241 79560 35275
rect 79508 35232 79560 35241
rect 79600 35232 79652 35284
rect 80244 35232 80296 35284
rect 81348 35275 81400 35284
rect 81348 35241 81357 35275
rect 81357 35241 81391 35275
rect 81391 35241 81400 35275
rect 81348 35232 81400 35241
rect 84752 35232 84804 35284
rect 140688 35232 140740 35284
rect 35532 35164 35584 35216
rect 36636 35164 36688 35216
rect 41696 35207 41748 35216
rect 41696 35173 41705 35207
rect 41705 35173 41739 35207
rect 41739 35173 41748 35207
rect 41696 35164 41748 35173
rect 43076 35164 43128 35216
rect 43996 35164 44048 35216
rect 35348 35096 35400 35148
rect 44456 35096 44508 35148
rect 57060 35096 57112 35148
rect 58532 35096 58584 35148
rect 59912 35139 59964 35148
rect 59912 35105 59921 35139
rect 59921 35105 59955 35139
rect 59955 35105 59964 35139
rect 59912 35096 59964 35105
rect 62120 35096 62172 35148
rect 62856 35096 62908 35148
rect 64144 35096 64196 35148
rect 65340 35096 65392 35148
rect 68560 35096 68612 35148
rect 17960 35028 18012 35080
rect 36544 35028 36596 35080
rect 36912 35028 36964 35080
rect 43352 35028 43404 35080
rect 44548 35028 44600 35080
rect 63684 35028 63736 35080
rect 65248 35071 65300 35080
rect 65248 35037 65257 35071
rect 65257 35037 65291 35071
rect 65291 35037 65300 35071
rect 65248 35028 65300 35037
rect 80060 35096 80112 35148
rect 30656 34960 30708 35012
rect 44456 34960 44508 35012
rect 25320 34892 25372 34944
rect 25688 34892 25740 34944
rect 40868 34892 40920 34944
rect 42800 34935 42852 34944
rect 42800 34901 42809 34935
rect 42809 34901 42843 34935
rect 42843 34901 42852 34935
rect 47124 34960 47176 35012
rect 48228 34960 48280 35012
rect 49792 34960 49844 35012
rect 51172 34960 51224 35012
rect 53196 34960 53248 35012
rect 54392 34960 54444 35012
rect 92388 34960 92440 35012
rect 45652 34935 45704 34944
rect 42800 34892 42852 34901
rect 45652 34901 45661 34935
rect 45661 34901 45695 34935
rect 45695 34901 45704 34935
rect 45652 34892 45704 34901
rect 46020 34892 46072 34944
rect 60740 34935 60792 34944
rect 60740 34901 60749 34935
rect 60749 34901 60783 34935
rect 60783 34901 60792 34935
rect 61200 34935 61252 34944
rect 60740 34892 60792 34901
rect 61200 34901 61209 34935
rect 61209 34901 61243 34935
rect 61243 34901 61252 34935
rect 61200 34892 61252 34901
rect 61752 34892 61804 34944
rect 62028 34892 62080 34944
rect 62580 34892 62632 34944
rect 64236 34892 64288 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 81014 34790 81066 34842
rect 81078 34790 81130 34842
rect 81142 34790 81194 34842
rect 81206 34790 81258 34842
rect 81270 34790 81322 34842
rect 111734 34790 111786 34842
rect 111798 34790 111850 34842
rect 111862 34790 111914 34842
rect 111926 34790 111978 34842
rect 111990 34790 112042 34842
rect 142454 34790 142506 34842
rect 142518 34790 142570 34842
rect 142582 34790 142634 34842
rect 142646 34790 142698 34842
rect 142710 34790 142762 34842
rect 29092 34688 29144 34740
rect 47032 34688 47084 34740
rect 59268 34688 59320 34740
rect 102876 34688 102928 34740
rect 43812 34663 43864 34672
rect 43812 34629 43821 34663
rect 43821 34629 43855 34663
rect 43855 34629 43864 34663
rect 43812 34620 43864 34629
rect 24584 34484 24636 34536
rect 24768 34484 24820 34536
rect 69020 34484 69072 34536
rect 69204 34484 69256 34536
rect 57520 34416 57572 34468
rect 124036 34416 124088 34468
rect 83096 34348 83148 34400
rect 144000 34348 144052 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 65654 34246 65706 34298
rect 65718 34246 65770 34298
rect 65782 34246 65834 34298
rect 65846 34246 65898 34298
rect 65910 34246 65962 34298
rect 96374 34246 96426 34298
rect 96438 34246 96490 34298
rect 96502 34246 96554 34298
rect 96566 34246 96618 34298
rect 96630 34246 96682 34298
rect 127094 34246 127146 34298
rect 127158 34246 127210 34298
rect 127222 34246 127274 34298
rect 127286 34246 127338 34298
rect 127350 34246 127402 34298
rect 75828 34144 75880 34196
rect 113456 34144 113508 34196
rect 38844 34076 38896 34128
rect 81900 34076 81952 34128
rect 81992 34076 82044 34128
rect 83832 34076 83884 34128
rect 61016 34008 61068 34060
rect 107752 34008 107804 34060
rect 66076 33940 66128 33992
rect 109592 33940 109644 33992
rect 69664 33872 69716 33924
rect 112168 33872 112220 33924
rect 72608 33804 72660 33856
rect 105912 33804 105964 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 81014 33702 81066 33754
rect 81078 33702 81130 33754
rect 81142 33702 81194 33754
rect 81206 33702 81258 33754
rect 81270 33702 81322 33754
rect 111734 33702 111786 33754
rect 111798 33702 111850 33754
rect 111862 33702 111914 33754
rect 111926 33702 111978 33754
rect 111990 33702 112042 33754
rect 142454 33702 142506 33754
rect 142518 33702 142570 33754
rect 142582 33702 142634 33754
rect 142646 33702 142698 33754
rect 142710 33702 142762 33754
rect 46204 33600 46256 33652
rect 79140 33600 79192 33652
rect 81900 33600 81952 33652
rect 89628 33600 89680 33652
rect 25964 33532 26016 33584
rect 86868 33532 86920 33584
rect 21364 33464 21416 33516
rect 83188 33464 83240 33516
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 65654 33158 65706 33210
rect 65718 33158 65770 33210
rect 65782 33158 65834 33210
rect 65846 33158 65898 33210
rect 65910 33158 65962 33210
rect 96374 33158 96426 33210
rect 96438 33158 96490 33210
rect 96502 33158 96554 33210
rect 96566 33158 96618 33210
rect 96630 33158 96682 33210
rect 127094 33158 127146 33210
rect 127158 33158 127210 33210
rect 127222 33158 127274 33210
rect 127286 33158 127338 33210
rect 127350 33158 127402 33210
rect 55864 33056 55916 33108
rect 56784 33056 56836 33108
rect 77760 33056 77812 33108
rect 147404 33056 147456 33108
rect 51540 32988 51592 33040
rect 114560 32988 114612 33040
rect 26516 32920 26568 32972
rect 88064 32920 88116 32972
rect 48136 32852 48188 32904
rect 108764 32852 108816 32904
rect 32496 32784 32548 32836
rect 91560 32784 91612 32836
rect 44824 32716 44876 32768
rect 98000 32716 98052 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 81014 32614 81066 32666
rect 81078 32614 81130 32666
rect 81142 32614 81194 32666
rect 81206 32614 81258 32666
rect 81270 32614 81322 32666
rect 111734 32614 111786 32666
rect 111798 32614 111850 32666
rect 111862 32614 111914 32666
rect 111926 32614 111978 32666
rect 111990 32614 112042 32666
rect 142454 32614 142506 32666
rect 142518 32614 142570 32666
rect 142582 32614 142634 32666
rect 142646 32614 142698 32666
rect 142710 32614 142762 32666
rect 49148 32376 49200 32428
rect 100760 32512 100812 32564
rect 52920 32444 52972 32496
rect 104440 32444 104492 32496
rect 57152 32308 57204 32360
rect 106280 32376 106332 32428
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 65654 32070 65706 32122
rect 65718 32070 65770 32122
rect 65782 32070 65834 32122
rect 65846 32070 65898 32122
rect 65910 32070 65962 32122
rect 96374 32070 96426 32122
rect 96438 32070 96490 32122
rect 96502 32070 96554 32122
rect 96566 32070 96618 32122
rect 96630 32070 96682 32122
rect 127094 32070 127146 32122
rect 127158 32070 127210 32122
rect 127222 32070 127274 32122
rect 127286 32070 127338 32122
rect 127350 32070 127402 32122
rect 62672 31696 62724 31748
rect 96160 31696 96212 31748
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 81014 31526 81066 31578
rect 81078 31526 81130 31578
rect 81142 31526 81194 31578
rect 81206 31526 81258 31578
rect 81270 31526 81322 31578
rect 111734 31526 111786 31578
rect 111798 31526 111850 31578
rect 111862 31526 111914 31578
rect 111926 31526 111978 31578
rect 111990 31526 112042 31578
rect 142454 31526 142506 31578
rect 142518 31526 142570 31578
rect 142582 31526 142634 31578
rect 142646 31526 142698 31578
rect 142710 31526 142762 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 65654 30982 65706 31034
rect 65718 30982 65770 31034
rect 65782 30982 65834 31034
rect 65846 30982 65898 31034
rect 65910 30982 65962 31034
rect 96374 30982 96426 31034
rect 96438 30982 96490 31034
rect 96502 30982 96554 31034
rect 96566 30982 96618 31034
rect 96630 30982 96682 31034
rect 127094 30982 127146 31034
rect 127158 30982 127210 31034
rect 127222 30982 127274 31034
rect 127286 30982 127338 31034
rect 127350 30982 127402 31034
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 81014 30438 81066 30490
rect 81078 30438 81130 30490
rect 81142 30438 81194 30490
rect 81206 30438 81258 30490
rect 81270 30438 81322 30490
rect 111734 30438 111786 30490
rect 111798 30438 111850 30490
rect 111862 30438 111914 30490
rect 111926 30438 111978 30490
rect 111990 30438 112042 30490
rect 142454 30438 142506 30490
rect 142518 30438 142570 30490
rect 142582 30438 142634 30490
rect 142646 30438 142698 30490
rect 142710 30438 142762 30490
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 65654 29894 65706 29946
rect 65718 29894 65770 29946
rect 65782 29894 65834 29946
rect 65846 29894 65898 29946
rect 65910 29894 65962 29946
rect 96374 29894 96426 29946
rect 96438 29894 96490 29946
rect 96502 29894 96554 29946
rect 96566 29894 96618 29946
rect 96630 29894 96682 29946
rect 127094 29894 127146 29946
rect 127158 29894 127210 29946
rect 127222 29894 127274 29946
rect 127286 29894 127338 29946
rect 127350 29894 127402 29946
rect 31760 29588 31812 29640
rect 61200 29588 61252 29640
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 81014 29350 81066 29402
rect 81078 29350 81130 29402
rect 81142 29350 81194 29402
rect 81206 29350 81258 29402
rect 81270 29350 81322 29402
rect 111734 29350 111786 29402
rect 111798 29350 111850 29402
rect 111862 29350 111914 29402
rect 111926 29350 111978 29402
rect 111990 29350 112042 29402
rect 142454 29350 142506 29402
rect 142518 29350 142570 29402
rect 142582 29350 142634 29402
rect 142646 29350 142698 29402
rect 142710 29350 142762 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 65654 28806 65706 28858
rect 65718 28806 65770 28858
rect 65782 28806 65834 28858
rect 65846 28806 65898 28858
rect 65910 28806 65962 28858
rect 96374 28806 96426 28858
rect 96438 28806 96490 28858
rect 96502 28806 96554 28858
rect 96566 28806 96618 28858
rect 96630 28806 96682 28858
rect 127094 28806 127146 28858
rect 127158 28806 127210 28858
rect 127222 28806 127274 28858
rect 127286 28806 127338 28858
rect 127350 28806 127402 28858
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 81014 28262 81066 28314
rect 81078 28262 81130 28314
rect 81142 28262 81194 28314
rect 81206 28262 81258 28314
rect 81270 28262 81322 28314
rect 111734 28262 111786 28314
rect 111798 28262 111850 28314
rect 111862 28262 111914 28314
rect 111926 28262 111978 28314
rect 111990 28262 112042 28314
rect 142454 28262 142506 28314
rect 142518 28262 142570 28314
rect 142582 28262 142634 28314
rect 142646 28262 142698 28314
rect 142710 28262 142762 28314
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 65654 27718 65706 27770
rect 65718 27718 65770 27770
rect 65782 27718 65834 27770
rect 65846 27718 65898 27770
rect 65910 27718 65962 27770
rect 96374 27718 96426 27770
rect 96438 27718 96490 27770
rect 96502 27718 96554 27770
rect 96566 27718 96618 27770
rect 96630 27718 96682 27770
rect 127094 27718 127146 27770
rect 127158 27718 127210 27770
rect 127222 27718 127274 27770
rect 127286 27718 127338 27770
rect 127350 27718 127402 27770
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 81014 27174 81066 27226
rect 81078 27174 81130 27226
rect 81142 27174 81194 27226
rect 81206 27174 81258 27226
rect 81270 27174 81322 27226
rect 111734 27174 111786 27226
rect 111798 27174 111850 27226
rect 111862 27174 111914 27226
rect 111926 27174 111978 27226
rect 111990 27174 112042 27226
rect 142454 27174 142506 27226
rect 142518 27174 142570 27226
rect 142582 27174 142634 27226
rect 142646 27174 142698 27226
rect 142710 27174 142762 27226
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 65654 26630 65706 26682
rect 65718 26630 65770 26682
rect 65782 26630 65834 26682
rect 65846 26630 65898 26682
rect 65910 26630 65962 26682
rect 96374 26630 96426 26682
rect 96438 26630 96490 26682
rect 96502 26630 96554 26682
rect 96566 26630 96618 26682
rect 96630 26630 96682 26682
rect 127094 26630 127146 26682
rect 127158 26630 127210 26682
rect 127222 26630 127274 26682
rect 127286 26630 127338 26682
rect 127350 26630 127402 26682
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 81014 26086 81066 26138
rect 81078 26086 81130 26138
rect 81142 26086 81194 26138
rect 81206 26086 81258 26138
rect 81270 26086 81322 26138
rect 111734 26086 111786 26138
rect 111798 26086 111850 26138
rect 111862 26086 111914 26138
rect 111926 26086 111978 26138
rect 111990 26086 112042 26138
rect 142454 26086 142506 26138
rect 142518 26086 142570 26138
rect 142582 26086 142634 26138
rect 142646 26086 142698 26138
rect 142710 26086 142762 26138
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 65654 25542 65706 25594
rect 65718 25542 65770 25594
rect 65782 25542 65834 25594
rect 65846 25542 65898 25594
rect 65910 25542 65962 25594
rect 96374 25542 96426 25594
rect 96438 25542 96490 25594
rect 96502 25542 96554 25594
rect 96566 25542 96618 25594
rect 96630 25542 96682 25594
rect 127094 25542 127146 25594
rect 127158 25542 127210 25594
rect 127222 25542 127274 25594
rect 127286 25542 127338 25594
rect 127350 25542 127402 25594
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 81014 24998 81066 25050
rect 81078 24998 81130 25050
rect 81142 24998 81194 25050
rect 81206 24998 81258 25050
rect 81270 24998 81322 25050
rect 111734 24998 111786 25050
rect 111798 24998 111850 25050
rect 111862 24998 111914 25050
rect 111926 24998 111978 25050
rect 111990 24998 112042 25050
rect 142454 24998 142506 25050
rect 142518 24998 142570 25050
rect 142582 24998 142634 25050
rect 142646 24998 142698 25050
rect 142710 24998 142762 25050
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 65654 24454 65706 24506
rect 65718 24454 65770 24506
rect 65782 24454 65834 24506
rect 65846 24454 65898 24506
rect 65910 24454 65962 24506
rect 96374 24454 96426 24506
rect 96438 24454 96490 24506
rect 96502 24454 96554 24506
rect 96566 24454 96618 24506
rect 96630 24454 96682 24506
rect 127094 24454 127146 24506
rect 127158 24454 127210 24506
rect 127222 24454 127274 24506
rect 127286 24454 127338 24506
rect 127350 24454 127402 24506
rect 73712 24148 73764 24200
rect 75092 24148 75144 24200
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 81014 23910 81066 23962
rect 81078 23910 81130 23962
rect 81142 23910 81194 23962
rect 81206 23910 81258 23962
rect 81270 23910 81322 23962
rect 111734 23910 111786 23962
rect 111798 23910 111850 23962
rect 111862 23910 111914 23962
rect 111926 23910 111978 23962
rect 111990 23910 112042 23962
rect 142454 23910 142506 23962
rect 142518 23910 142570 23962
rect 142582 23910 142634 23962
rect 142646 23910 142698 23962
rect 142710 23910 142762 23962
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 65654 23366 65706 23418
rect 65718 23366 65770 23418
rect 65782 23366 65834 23418
rect 65846 23366 65898 23418
rect 65910 23366 65962 23418
rect 96374 23366 96426 23418
rect 96438 23366 96490 23418
rect 96502 23366 96554 23418
rect 96566 23366 96618 23418
rect 96630 23366 96682 23418
rect 127094 23366 127146 23418
rect 127158 23366 127210 23418
rect 127222 23366 127274 23418
rect 127286 23366 127338 23418
rect 127350 23366 127402 23418
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 81014 22822 81066 22874
rect 81078 22822 81130 22874
rect 81142 22822 81194 22874
rect 81206 22822 81258 22874
rect 81270 22822 81322 22874
rect 111734 22822 111786 22874
rect 111798 22822 111850 22874
rect 111862 22822 111914 22874
rect 111926 22822 111978 22874
rect 111990 22822 112042 22874
rect 142454 22822 142506 22874
rect 142518 22822 142570 22874
rect 142582 22822 142634 22874
rect 142646 22822 142698 22874
rect 142710 22822 142762 22874
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 65654 22278 65706 22330
rect 65718 22278 65770 22330
rect 65782 22278 65834 22330
rect 65846 22278 65898 22330
rect 65910 22278 65962 22330
rect 96374 22278 96426 22330
rect 96438 22278 96490 22330
rect 96502 22278 96554 22330
rect 96566 22278 96618 22330
rect 96630 22278 96682 22330
rect 127094 22278 127146 22330
rect 127158 22278 127210 22330
rect 127222 22278 127274 22330
rect 127286 22278 127338 22330
rect 127350 22278 127402 22330
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 81014 21734 81066 21786
rect 81078 21734 81130 21786
rect 81142 21734 81194 21786
rect 81206 21734 81258 21786
rect 81270 21734 81322 21786
rect 111734 21734 111786 21786
rect 111798 21734 111850 21786
rect 111862 21734 111914 21786
rect 111926 21734 111978 21786
rect 111990 21734 112042 21786
rect 142454 21734 142506 21786
rect 142518 21734 142570 21786
rect 142582 21734 142634 21786
rect 142646 21734 142698 21786
rect 142710 21734 142762 21786
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 65654 21190 65706 21242
rect 65718 21190 65770 21242
rect 65782 21190 65834 21242
rect 65846 21190 65898 21242
rect 65910 21190 65962 21242
rect 96374 21190 96426 21242
rect 96438 21190 96490 21242
rect 96502 21190 96554 21242
rect 96566 21190 96618 21242
rect 96630 21190 96682 21242
rect 127094 21190 127146 21242
rect 127158 21190 127210 21242
rect 127222 21190 127274 21242
rect 127286 21190 127338 21242
rect 127350 21190 127402 21242
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 81014 20646 81066 20698
rect 81078 20646 81130 20698
rect 81142 20646 81194 20698
rect 81206 20646 81258 20698
rect 81270 20646 81322 20698
rect 111734 20646 111786 20698
rect 111798 20646 111850 20698
rect 111862 20646 111914 20698
rect 111926 20646 111978 20698
rect 111990 20646 112042 20698
rect 142454 20646 142506 20698
rect 142518 20646 142570 20698
rect 142582 20646 142634 20698
rect 142646 20646 142698 20698
rect 142710 20646 142762 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 65654 20102 65706 20154
rect 65718 20102 65770 20154
rect 65782 20102 65834 20154
rect 65846 20102 65898 20154
rect 65910 20102 65962 20154
rect 96374 20102 96426 20154
rect 96438 20102 96490 20154
rect 96502 20102 96554 20154
rect 96566 20102 96618 20154
rect 96630 20102 96682 20154
rect 127094 20102 127146 20154
rect 127158 20102 127210 20154
rect 127222 20102 127274 20154
rect 127286 20102 127338 20154
rect 127350 20102 127402 20154
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 81014 19558 81066 19610
rect 81078 19558 81130 19610
rect 81142 19558 81194 19610
rect 81206 19558 81258 19610
rect 81270 19558 81322 19610
rect 111734 19558 111786 19610
rect 111798 19558 111850 19610
rect 111862 19558 111914 19610
rect 111926 19558 111978 19610
rect 111990 19558 112042 19610
rect 142454 19558 142506 19610
rect 142518 19558 142570 19610
rect 142582 19558 142634 19610
rect 142646 19558 142698 19610
rect 142710 19558 142762 19610
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 65654 19014 65706 19066
rect 65718 19014 65770 19066
rect 65782 19014 65834 19066
rect 65846 19014 65898 19066
rect 65910 19014 65962 19066
rect 96374 19014 96426 19066
rect 96438 19014 96490 19066
rect 96502 19014 96554 19066
rect 96566 19014 96618 19066
rect 96630 19014 96682 19066
rect 127094 19014 127146 19066
rect 127158 19014 127210 19066
rect 127222 19014 127274 19066
rect 127286 19014 127338 19066
rect 127350 19014 127402 19066
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 81014 18470 81066 18522
rect 81078 18470 81130 18522
rect 81142 18470 81194 18522
rect 81206 18470 81258 18522
rect 81270 18470 81322 18522
rect 111734 18470 111786 18522
rect 111798 18470 111850 18522
rect 111862 18470 111914 18522
rect 111926 18470 111978 18522
rect 111990 18470 112042 18522
rect 142454 18470 142506 18522
rect 142518 18470 142570 18522
rect 142582 18470 142634 18522
rect 142646 18470 142698 18522
rect 142710 18470 142762 18522
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 65654 17926 65706 17978
rect 65718 17926 65770 17978
rect 65782 17926 65834 17978
rect 65846 17926 65898 17978
rect 65910 17926 65962 17978
rect 96374 17926 96426 17978
rect 96438 17926 96490 17978
rect 96502 17926 96554 17978
rect 96566 17926 96618 17978
rect 96630 17926 96682 17978
rect 127094 17926 127146 17978
rect 127158 17926 127210 17978
rect 127222 17926 127274 17978
rect 127286 17926 127338 17978
rect 127350 17926 127402 17978
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 81014 17382 81066 17434
rect 81078 17382 81130 17434
rect 81142 17382 81194 17434
rect 81206 17382 81258 17434
rect 81270 17382 81322 17434
rect 111734 17382 111786 17434
rect 111798 17382 111850 17434
rect 111862 17382 111914 17434
rect 111926 17382 111978 17434
rect 111990 17382 112042 17434
rect 142454 17382 142506 17434
rect 142518 17382 142570 17434
rect 142582 17382 142634 17434
rect 142646 17382 142698 17434
rect 142710 17382 142762 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 65654 16838 65706 16890
rect 65718 16838 65770 16890
rect 65782 16838 65834 16890
rect 65846 16838 65898 16890
rect 65910 16838 65962 16890
rect 96374 16838 96426 16890
rect 96438 16838 96490 16890
rect 96502 16838 96554 16890
rect 96566 16838 96618 16890
rect 96630 16838 96682 16890
rect 127094 16838 127146 16890
rect 127158 16838 127210 16890
rect 127222 16838 127274 16890
rect 127286 16838 127338 16890
rect 127350 16838 127402 16890
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 81014 16294 81066 16346
rect 81078 16294 81130 16346
rect 81142 16294 81194 16346
rect 81206 16294 81258 16346
rect 81270 16294 81322 16346
rect 111734 16294 111786 16346
rect 111798 16294 111850 16346
rect 111862 16294 111914 16346
rect 111926 16294 111978 16346
rect 111990 16294 112042 16346
rect 142454 16294 142506 16346
rect 142518 16294 142570 16346
rect 142582 16294 142634 16346
rect 142646 16294 142698 16346
rect 142710 16294 142762 16346
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 65654 15750 65706 15802
rect 65718 15750 65770 15802
rect 65782 15750 65834 15802
rect 65846 15750 65898 15802
rect 65910 15750 65962 15802
rect 96374 15750 96426 15802
rect 96438 15750 96490 15802
rect 96502 15750 96554 15802
rect 96566 15750 96618 15802
rect 96630 15750 96682 15802
rect 127094 15750 127146 15802
rect 127158 15750 127210 15802
rect 127222 15750 127274 15802
rect 127286 15750 127338 15802
rect 127350 15750 127402 15802
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 81014 15206 81066 15258
rect 81078 15206 81130 15258
rect 81142 15206 81194 15258
rect 81206 15206 81258 15258
rect 81270 15206 81322 15258
rect 111734 15206 111786 15258
rect 111798 15206 111850 15258
rect 111862 15206 111914 15258
rect 111926 15206 111978 15258
rect 111990 15206 112042 15258
rect 142454 15206 142506 15258
rect 142518 15206 142570 15258
rect 142582 15206 142634 15258
rect 142646 15206 142698 15258
rect 142710 15206 142762 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 65654 14662 65706 14714
rect 65718 14662 65770 14714
rect 65782 14662 65834 14714
rect 65846 14662 65898 14714
rect 65910 14662 65962 14714
rect 96374 14662 96426 14714
rect 96438 14662 96490 14714
rect 96502 14662 96554 14714
rect 96566 14662 96618 14714
rect 96630 14662 96682 14714
rect 127094 14662 127146 14714
rect 127158 14662 127210 14714
rect 127222 14662 127274 14714
rect 127286 14662 127338 14714
rect 127350 14662 127402 14714
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 81014 14118 81066 14170
rect 81078 14118 81130 14170
rect 81142 14118 81194 14170
rect 81206 14118 81258 14170
rect 81270 14118 81322 14170
rect 111734 14118 111786 14170
rect 111798 14118 111850 14170
rect 111862 14118 111914 14170
rect 111926 14118 111978 14170
rect 111990 14118 112042 14170
rect 142454 14118 142506 14170
rect 142518 14118 142570 14170
rect 142582 14118 142634 14170
rect 142646 14118 142698 14170
rect 142710 14118 142762 14170
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 65654 13574 65706 13626
rect 65718 13574 65770 13626
rect 65782 13574 65834 13626
rect 65846 13574 65898 13626
rect 65910 13574 65962 13626
rect 96374 13574 96426 13626
rect 96438 13574 96490 13626
rect 96502 13574 96554 13626
rect 96566 13574 96618 13626
rect 96630 13574 96682 13626
rect 127094 13574 127146 13626
rect 127158 13574 127210 13626
rect 127222 13574 127274 13626
rect 127286 13574 127338 13626
rect 127350 13574 127402 13626
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 81014 13030 81066 13082
rect 81078 13030 81130 13082
rect 81142 13030 81194 13082
rect 81206 13030 81258 13082
rect 81270 13030 81322 13082
rect 111734 13030 111786 13082
rect 111798 13030 111850 13082
rect 111862 13030 111914 13082
rect 111926 13030 111978 13082
rect 111990 13030 112042 13082
rect 142454 13030 142506 13082
rect 142518 13030 142570 13082
rect 142582 13030 142634 13082
rect 142646 13030 142698 13082
rect 142710 13030 142762 13082
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 65654 12486 65706 12538
rect 65718 12486 65770 12538
rect 65782 12486 65834 12538
rect 65846 12486 65898 12538
rect 65910 12486 65962 12538
rect 96374 12486 96426 12538
rect 96438 12486 96490 12538
rect 96502 12486 96554 12538
rect 96566 12486 96618 12538
rect 96630 12486 96682 12538
rect 127094 12486 127146 12538
rect 127158 12486 127210 12538
rect 127222 12486 127274 12538
rect 127286 12486 127338 12538
rect 127350 12486 127402 12538
rect 9588 12248 9640 12300
rect 15384 12248 15436 12300
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 81014 11942 81066 11994
rect 81078 11942 81130 11994
rect 81142 11942 81194 11994
rect 81206 11942 81258 11994
rect 81270 11942 81322 11994
rect 111734 11942 111786 11994
rect 111798 11942 111850 11994
rect 111862 11942 111914 11994
rect 111926 11942 111978 11994
rect 111990 11942 112042 11994
rect 142454 11942 142506 11994
rect 142518 11942 142570 11994
rect 142582 11942 142634 11994
rect 142646 11942 142698 11994
rect 142710 11942 142762 11994
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 65654 11398 65706 11450
rect 65718 11398 65770 11450
rect 65782 11398 65834 11450
rect 65846 11398 65898 11450
rect 65910 11398 65962 11450
rect 96374 11398 96426 11450
rect 96438 11398 96490 11450
rect 96502 11398 96554 11450
rect 96566 11398 96618 11450
rect 96630 11398 96682 11450
rect 127094 11398 127146 11450
rect 127158 11398 127210 11450
rect 127222 11398 127274 11450
rect 127286 11398 127338 11450
rect 127350 11398 127402 11450
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 81014 10854 81066 10906
rect 81078 10854 81130 10906
rect 81142 10854 81194 10906
rect 81206 10854 81258 10906
rect 81270 10854 81322 10906
rect 111734 10854 111786 10906
rect 111798 10854 111850 10906
rect 111862 10854 111914 10906
rect 111926 10854 111978 10906
rect 111990 10854 112042 10906
rect 142454 10854 142506 10906
rect 142518 10854 142570 10906
rect 142582 10854 142634 10906
rect 142646 10854 142698 10906
rect 142710 10854 142762 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 65654 10310 65706 10362
rect 65718 10310 65770 10362
rect 65782 10310 65834 10362
rect 65846 10310 65898 10362
rect 65910 10310 65962 10362
rect 96374 10310 96426 10362
rect 96438 10310 96490 10362
rect 96502 10310 96554 10362
rect 96566 10310 96618 10362
rect 96630 10310 96682 10362
rect 127094 10310 127146 10362
rect 127158 10310 127210 10362
rect 127222 10310 127274 10362
rect 127286 10310 127338 10362
rect 127350 10310 127402 10362
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 81014 9766 81066 9818
rect 81078 9766 81130 9818
rect 81142 9766 81194 9818
rect 81206 9766 81258 9818
rect 81270 9766 81322 9818
rect 111734 9766 111786 9818
rect 111798 9766 111850 9818
rect 111862 9766 111914 9818
rect 111926 9766 111978 9818
rect 111990 9766 112042 9818
rect 142454 9766 142506 9818
rect 142518 9766 142570 9818
rect 142582 9766 142634 9818
rect 142646 9766 142698 9818
rect 142710 9766 142762 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 65654 9222 65706 9274
rect 65718 9222 65770 9274
rect 65782 9222 65834 9274
rect 65846 9222 65898 9274
rect 65910 9222 65962 9274
rect 96374 9222 96426 9274
rect 96438 9222 96490 9274
rect 96502 9222 96554 9274
rect 96566 9222 96618 9274
rect 96630 9222 96682 9274
rect 127094 9222 127146 9274
rect 127158 9222 127210 9274
rect 127222 9222 127274 9274
rect 127286 9222 127338 9274
rect 127350 9222 127402 9274
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 81014 8678 81066 8730
rect 81078 8678 81130 8730
rect 81142 8678 81194 8730
rect 81206 8678 81258 8730
rect 81270 8678 81322 8730
rect 111734 8678 111786 8730
rect 111798 8678 111850 8730
rect 111862 8678 111914 8730
rect 111926 8678 111978 8730
rect 111990 8678 112042 8730
rect 142454 8678 142506 8730
rect 142518 8678 142570 8730
rect 142582 8678 142634 8730
rect 142646 8678 142698 8730
rect 142710 8678 142762 8730
rect 66812 8304 66864 8356
rect 67640 8304 67692 8356
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 65654 8134 65706 8186
rect 65718 8134 65770 8186
rect 65782 8134 65834 8186
rect 65846 8134 65898 8186
rect 65910 8134 65962 8186
rect 96374 8134 96426 8186
rect 96438 8134 96490 8186
rect 96502 8134 96554 8186
rect 96566 8134 96618 8186
rect 96630 8134 96682 8186
rect 127094 8134 127146 8186
rect 127158 8134 127210 8186
rect 127222 8134 127274 8186
rect 127286 8134 127338 8186
rect 127350 8134 127402 8186
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 81014 7590 81066 7642
rect 81078 7590 81130 7642
rect 81142 7590 81194 7642
rect 81206 7590 81258 7642
rect 81270 7590 81322 7642
rect 111734 7590 111786 7642
rect 111798 7590 111850 7642
rect 111862 7590 111914 7642
rect 111926 7590 111978 7642
rect 111990 7590 112042 7642
rect 142454 7590 142506 7642
rect 142518 7590 142570 7642
rect 142582 7590 142634 7642
rect 142646 7590 142698 7642
rect 142710 7590 142762 7642
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 65654 7046 65706 7098
rect 65718 7046 65770 7098
rect 65782 7046 65834 7098
rect 65846 7046 65898 7098
rect 65910 7046 65962 7098
rect 96374 7046 96426 7098
rect 96438 7046 96490 7098
rect 96502 7046 96554 7098
rect 96566 7046 96618 7098
rect 96630 7046 96682 7098
rect 127094 7046 127146 7098
rect 127158 7046 127210 7098
rect 127222 7046 127274 7098
rect 127286 7046 127338 7098
rect 127350 7046 127402 7098
rect 82452 6808 82504 6860
rect 83096 6808 83148 6860
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 81014 6502 81066 6554
rect 81078 6502 81130 6554
rect 81142 6502 81194 6554
rect 81206 6502 81258 6554
rect 81270 6502 81322 6554
rect 111734 6502 111786 6554
rect 111798 6502 111850 6554
rect 111862 6502 111914 6554
rect 111926 6502 111978 6554
rect 111990 6502 112042 6554
rect 142454 6502 142506 6554
rect 142518 6502 142570 6554
rect 142582 6502 142634 6554
rect 142646 6502 142698 6554
rect 142710 6502 142762 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 65654 5958 65706 6010
rect 65718 5958 65770 6010
rect 65782 5958 65834 6010
rect 65846 5958 65898 6010
rect 65910 5958 65962 6010
rect 96374 5958 96426 6010
rect 96438 5958 96490 6010
rect 96502 5958 96554 6010
rect 96566 5958 96618 6010
rect 96630 5958 96682 6010
rect 127094 5958 127146 6010
rect 127158 5958 127210 6010
rect 127222 5958 127274 6010
rect 127286 5958 127338 6010
rect 127350 5958 127402 6010
rect 64052 5899 64104 5908
rect 64052 5865 64061 5899
rect 64061 5865 64095 5899
rect 64095 5865 64104 5899
rect 64052 5856 64104 5865
rect 65524 5856 65576 5908
rect 80060 5899 80112 5908
rect 80060 5865 80069 5899
rect 80069 5865 80103 5899
rect 80103 5865 80112 5899
rect 80060 5856 80112 5865
rect 78220 5652 78272 5704
rect 79048 5652 79100 5704
rect 65156 5559 65208 5568
rect 65156 5525 65165 5559
rect 65165 5525 65199 5559
rect 65199 5525 65208 5559
rect 65156 5516 65208 5525
rect 69480 5559 69532 5568
rect 69480 5525 69489 5559
rect 69489 5525 69523 5559
rect 69523 5525 69532 5559
rect 69480 5516 69532 5525
rect 75736 5516 75788 5568
rect 76472 5516 76524 5568
rect 77208 5516 77260 5568
rect 78496 5516 78548 5568
rect 79140 5516 79192 5568
rect 80152 5516 80204 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 81014 5414 81066 5466
rect 81078 5414 81130 5466
rect 81142 5414 81194 5466
rect 81206 5414 81258 5466
rect 81270 5414 81322 5466
rect 111734 5414 111786 5466
rect 111798 5414 111850 5466
rect 111862 5414 111914 5466
rect 111926 5414 111978 5466
rect 111990 5414 112042 5466
rect 142454 5414 142506 5466
rect 142518 5414 142570 5466
rect 142582 5414 142634 5466
rect 142646 5414 142698 5466
rect 142710 5414 142762 5466
rect 28356 5355 28408 5364
rect 28356 5321 28365 5355
rect 28365 5321 28399 5355
rect 28399 5321 28408 5355
rect 28356 5312 28408 5321
rect 36084 5355 36136 5364
rect 36084 5321 36093 5355
rect 36093 5321 36127 5355
rect 36127 5321 36136 5355
rect 36084 5312 36136 5321
rect 38200 5312 38252 5364
rect 52092 5312 52144 5364
rect 52368 5312 52420 5364
rect 63500 5312 63552 5364
rect 66076 5312 66128 5364
rect 69112 5312 69164 5364
rect 69480 5312 69532 5364
rect 68192 5244 68244 5296
rect 34796 5040 34848 5092
rect 38568 5040 38620 5092
rect 35624 5015 35676 5024
rect 35624 4981 35633 5015
rect 35633 4981 35667 5015
rect 35667 4981 35676 5015
rect 35624 4972 35676 4981
rect 60832 5083 60884 5092
rect 60832 5049 60841 5083
rect 60841 5049 60875 5083
rect 60875 5049 60884 5083
rect 60832 5040 60884 5049
rect 79140 5040 79192 5092
rect 81716 5108 81768 5160
rect 81440 5040 81492 5092
rect 83372 5040 83424 5092
rect 42708 5015 42760 5024
rect 42708 4981 42717 5015
rect 42717 4981 42751 5015
rect 42751 4981 42760 5015
rect 42708 4972 42760 4981
rect 47124 5015 47176 5024
rect 47124 4981 47133 5015
rect 47133 4981 47167 5015
rect 47167 4981 47176 5015
rect 47124 4972 47176 4981
rect 48136 5015 48188 5024
rect 48136 4981 48145 5015
rect 48145 4981 48179 5015
rect 48179 4981 48188 5015
rect 48136 4972 48188 4981
rect 48320 4972 48372 5024
rect 49056 4972 49108 5024
rect 49608 4972 49660 5024
rect 53012 5015 53064 5024
rect 53012 4981 53021 5015
rect 53021 4981 53055 5015
rect 53055 4981 53064 5015
rect 53012 4972 53064 4981
rect 58072 5015 58124 5024
rect 58072 4981 58081 5015
rect 58081 4981 58115 5015
rect 58115 4981 58124 5015
rect 58072 4972 58124 4981
rect 58716 5015 58768 5024
rect 58716 4981 58725 5015
rect 58725 4981 58759 5015
rect 58759 4981 58768 5015
rect 58716 4972 58768 4981
rect 61844 5015 61896 5024
rect 61844 4981 61853 5015
rect 61853 4981 61887 5015
rect 61887 4981 61896 5015
rect 61844 4972 61896 4981
rect 64328 5015 64380 5024
rect 64328 4981 64337 5015
rect 64337 4981 64371 5015
rect 64371 4981 64380 5015
rect 64328 4972 64380 4981
rect 64880 5015 64932 5024
rect 64880 4981 64889 5015
rect 64889 4981 64923 5015
rect 64923 4981 64932 5015
rect 64880 4972 64932 4981
rect 65340 5015 65392 5024
rect 65340 4981 65349 5015
rect 65349 4981 65383 5015
rect 65383 4981 65392 5015
rect 65340 4972 65392 4981
rect 68928 4972 68980 5024
rect 69664 4972 69716 5024
rect 70308 4972 70360 5024
rect 79416 5015 79468 5024
rect 79416 4981 79425 5015
rect 79425 4981 79459 5015
rect 79459 4981 79468 5015
rect 79416 4972 79468 4981
rect 79508 4972 79560 5024
rect 80244 4972 80296 5024
rect 80796 4972 80848 5024
rect 81992 5015 82044 5024
rect 81992 4981 82001 5015
rect 82001 4981 82035 5015
rect 82035 4981 82044 5015
rect 81992 4972 82044 4981
rect 83004 5015 83056 5024
rect 83004 4981 83013 5015
rect 83013 4981 83047 5015
rect 83047 4981 83056 5015
rect 83004 4972 83056 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 65654 4870 65706 4922
rect 65718 4870 65770 4922
rect 65782 4870 65834 4922
rect 65846 4870 65898 4922
rect 65910 4870 65962 4922
rect 96374 4870 96426 4922
rect 96438 4870 96490 4922
rect 96502 4870 96554 4922
rect 96566 4870 96618 4922
rect 96630 4870 96682 4922
rect 127094 4870 127146 4922
rect 127158 4870 127210 4922
rect 127222 4870 127274 4922
rect 127286 4870 127338 4922
rect 127350 4870 127402 4922
rect 40592 4811 40644 4820
rect 40592 4777 40601 4811
rect 40601 4777 40635 4811
rect 40635 4777 40644 4811
rect 40592 4768 40644 4777
rect 42708 4768 42760 4820
rect 48596 4768 48648 4820
rect 48964 4811 49016 4820
rect 48964 4777 48973 4811
rect 48973 4777 49007 4811
rect 49007 4777 49016 4811
rect 48964 4768 49016 4777
rect 49516 4811 49568 4820
rect 49516 4777 49525 4811
rect 49525 4777 49559 4811
rect 49559 4777 49568 4811
rect 49516 4768 49568 4777
rect 53840 4811 53892 4820
rect 53840 4777 53849 4811
rect 53849 4777 53883 4811
rect 53883 4777 53892 4811
rect 53840 4768 53892 4777
rect 57980 4811 58032 4820
rect 57980 4777 57989 4811
rect 57989 4777 58023 4811
rect 58023 4777 58032 4811
rect 57980 4768 58032 4777
rect 58624 4768 58676 4820
rect 59084 4811 59136 4820
rect 59084 4777 59093 4811
rect 59093 4777 59127 4811
rect 59127 4777 59136 4811
rect 59084 4768 59136 4777
rect 61108 4811 61160 4820
rect 61108 4777 61117 4811
rect 61117 4777 61151 4811
rect 61151 4777 61160 4811
rect 61108 4768 61160 4777
rect 67640 4811 67692 4820
rect 67640 4777 67649 4811
rect 67649 4777 67683 4811
rect 67683 4777 67692 4811
rect 67640 4768 67692 4777
rect 68192 4811 68244 4820
rect 68192 4777 68201 4811
rect 68201 4777 68235 4811
rect 68235 4777 68244 4811
rect 68192 4768 68244 4777
rect 78220 4811 78272 4820
rect 78220 4777 78229 4811
rect 78229 4777 78263 4811
rect 78263 4777 78272 4811
rect 78220 4768 78272 4777
rect 83096 4811 83148 4820
rect 83096 4777 83105 4811
rect 83105 4777 83139 4811
rect 83139 4777 83148 4811
rect 83096 4768 83148 4777
rect 43444 4743 43496 4752
rect 43444 4709 43453 4743
rect 43453 4709 43487 4743
rect 43487 4709 43496 4743
rect 43444 4700 43496 4709
rect 36912 4632 36964 4684
rect 49608 4700 49660 4752
rect 66168 4700 66220 4752
rect 66536 4700 66588 4752
rect 81532 4700 81584 4752
rect 47584 4675 47636 4684
rect 47584 4641 47593 4675
rect 47593 4641 47627 4675
rect 47627 4641 47636 4675
rect 47584 4632 47636 4641
rect 48136 4632 48188 4684
rect 63316 4632 63368 4684
rect 78680 4632 78732 4684
rect 79784 4675 79836 4684
rect 79784 4641 79793 4675
rect 79793 4641 79827 4675
rect 79827 4641 79836 4675
rect 79784 4632 79836 4641
rect 26240 4564 26292 4616
rect 30288 4564 30340 4616
rect 38016 4607 38068 4616
rect 33692 4496 33744 4548
rect 38016 4573 38025 4607
rect 38025 4573 38059 4607
rect 38059 4573 38068 4607
rect 38016 4564 38068 4573
rect 39856 4564 39908 4616
rect 42432 4607 42484 4616
rect 42432 4573 42441 4607
rect 42441 4573 42475 4607
rect 42475 4573 42484 4607
rect 42432 4564 42484 4573
rect 47216 4564 47268 4616
rect 51448 4564 51500 4616
rect 58164 4564 58216 4616
rect 62212 4607 62264 4616
rect 62212 4573 62221 4607
rect 62221 4573 62255 4607
rect 62255 4573 62264 4607
rect 62212 4564 62264 4573
rect 65064 4607 65116 4616
rect 65064 4573 65073 4607
rect 65073 4573 65107 4607
rect 65107 4573 65116 4607
rect 65064 4564 65116 4573
rect 69848 4607 69900 4616
rect 69848 4573 69857 4607
rect 69857 4573 69891 4607
rect 69891 4573 69900 4607
rect 69848 4564 69900 4573
rect 36912 4496 36964 4548
rect 6368 4471 6420 4480
rect 6368 4437 6377 4471
rect 6377 4437 6411 4471
rect 6411 4437 6420 4471
rect 6368 4428 6420 4437
rect 23296 4428 23348 4480
rect 23848 4471 23900 4480
rect 23848 4437 23857 4471
rect 23857 4437 23891 4471
rect 23891 4437 23900 4471
rect 23848 4428 23900 4437
rect 27620 4471 27672 4480
rect 27620 4437 27629 4471
rect 27629 4437 27663 4471
rect 27663 4437 27672 4471
rect 27620 4428 27672 4437
rect 30196 4428 30248 4480
rect 32312 4428 32364 4480
rect 32772 4471 32824 4480
rect 32772 4437 32781 4471
rect 32781 4437 32815 4471
rect 32815 4437 32824 4471
rect 32772 4428 32824 4437
rect 35900 4471 35952 4480
rect 35900 4437 35909 4471
rect 35909 4437 35943 4471
rect 35943 4437 35952 4471
rect 37280 4471 37332 4480
rect 35900 4428 35952 4437
rect 37280 4437 37289 4471
rect 37289 4437 37323 4471
rect 37323 4437 37332 4471
rect 37280 4428 37332 4437
rect 38568 4428 38620 4480
rect 41328 4428 41380 4480
rect 42984 4428 43036 4480
rect 45928 4428 45980 4480
rect 47124 4496 47176 4548
rect 47584 4496 47636 4548
rect 48320 4496 48372 4548
rect 57796 4496 57848 4548
rect 71596 4564 71648 4616
rect 80060 4564 80112 4616
rect 80428 4607 80480 4616
rect 80428 4573 80437 4607
rect 80437 4573 80471 4607
rect 80471 4573 80480 4607
rect 80428 4564 80480 4573
rect 81992 4632 82044 4684
rect 82084 4607 82136 4616
rect 82084 4573 82093 4607
rect 82093 4573 82127 4607
rect 82127 4573 82136 4607
rect 82084 4564 82136 4573
rect 47032 4471 47084 4480
rect 47032 4437 47041 4471
rect 47041 4437 47075 4471
rect 47075 4437 47084 4471
rect 47032 4428 47084 4437
rect 50620 4428 50672 4480
rect 51632 4428 51684 4480
rect 52460 4428 52512 4480
rect 54300 4471 54352 4480
rect 54300 4437 54309 4471
rect 54309 4437 54343 4471
rect 54343 4437 54352 4471
rect 54300 4428 54352 4437
rect 56324 4428 56376 4480
rect 56416 4428 56468 4480
rect 58348 4428 58400 4480
rect 61476 4428 61528 4480
rect 62304 4471 62356 4480
rect 62304 4437 62313 4471
rect 62313 4437 62347 4471
rect 62347 4437 62356 4471
rect 62304 4428 62356 4437
rect 63408 4428 63460 4480
rect 70308 4496 70360 4548
rect 80336 4496 80388 4548
rect 64420 4471 64472 4480
rect 64420 4437 64429 4471
rect 64429 4437 64463 4471
rect 64463 4437 64472 4471
rect 64420 4428 64472 4437
rect 65248 4471 65300 4480
rect 65248 4437 65257 4471
rect 65257 4437 65291 4471
rect 65291 4437 65300 4471
rect 65248 4428 65300 4437
rect 68652 4471 68704 4480
rect 68652 4437 68661 4471
rect 68661 4437 68695 4471
rect 68695 4437 68704 4471
rect 68652 4428 68704 4437
rect 69204 4471 69256 4480
rect 69204 4437 69213 4471
rect 69213 4437 69247 4471
rect 69247 4437 69256 4471
rect 69204 4428 69256 4437
rect 70400 4428 70452 4480
rect 75092 4428 75144 4480
rect 77668 4471 77720 4480
rect 77668 4437 77677 4471
rect 77677 4437 77711 4471
rect 77711 4437 77720 4471
rect 77668 4428 77720 4437
rect 78680 4471 78732 4480
rect 78680 4437 78689 4471
rect 78689 4437 78723 4471
rect 78723 4437 78732 4471
rect 78680 4428 78732 4437
rect 78772 4428 78824 4480
rect 80152 4428 80204 4480
rect 81348 4471 81400 4480
rect 81348 4437 81357 4471
rect 81357 4437 81391 4471
rect 81391 4437 81400 4471
rect 81348 4428 81400 4437
rect 84200 4496 84252 4548
rect 82820 4428 82872 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 81014 4326 81066 4378
rect 81078 4326 81130 4378
rect 81142 4326 81194 4378
rect 81206 4326 81258 4378
rect 81270 4326 81322 4378
rect 111734 4326 111786 4378
rect 111798 4326 111850 4378
rect 111862 4326 111914 4378
rect 111926 4326 111978 4378
rect 111990 4326 112042 4378
rect 142454 4326 142506 4378
rect 142518 4326 142570 4378
rect 142582 4326 142634 4378
rect 142646 4326 142698 4378
rect 142710 4326 142762 4378
rect 32772 4224 32824 4276
rect 49056 4224 49108 4276
rect 54300 4224 54352 4276
rect 63408 4224 63460 4276
rect 64420 4224 64472 4276
rect 68284 4224 68336 4276
rect 68652 4224 68704 4276
rect 81440 4267 81492 4276
rect 81440 4233 81449 4267
rect 81449 4233 81483 4267
rect 81483 4233 81492 4267
rect 81440 4224 81492 4233
rect 82728 4224 82780 4276
rect 26332 4156 26384 4208
rect 6000 4088 6052 4140
rect 22744 4088 22796 4140
rect 27344 4131 27396 4140
rect 27344 4097 27353 4131
rect 27353 4097 27387 4131
rect 27387 4097 27396 4131
rect 27344 4088 27396 4097
rect 35624 4156 35676 4208
rect 37280 4156 37332 4208
rect 28448 4020 28500 4072
rect 6644 3952 6696 4004
rect 23756 3952 23808 4004
rect 26240 3952 26292 4004
rect 28816 4088 28868 4140
rect 33692 4088 33744 4140
rect 33784 4088 33836 4140
rect 34152 4088 34204 4140
rect 35992 4131 36044 4140
rect 35992 4097 36001 4131
rect 36001 4097 36035 4131
rect 36035 4097 36044 4131
rect 35992 4088 36044 4097
rect 37464 4088 37516 4140
rect 37648 4088 37700 4140
rect 38016 4088 38068 4140
rect 39856 4131 39908 4140
rect 39856 4097 39865 4131
rect 39865 4097 39899 4131
rect 39899 4097 39908 4131
rect 39856 4088 39908 4097
rect 40040 4088 40092 4140
rect 42156 4088 42208 4140
rect 43812 4088 43864 4140
rect 43904 4088 43956 4140
rect 49516 4156 49568 4208
rect 44364 4088 44416 4140
rect 47032 4131 47084 4140
rect 6276 3884 6328 3936
rect 6828 3884 6880 3936
rect 8024 3927 8076 3936
rect 8024 3893 8033 3927
rect 8033 3893 8067 3927
rect 8067 3893 8076 3927
rect 8024 3884 8076 3893
rect 22284 3927 22336 3936
rect 22284 3893 22293 3927
rect 22293 3893 22327 3927
rect 22327 3893 22336 3927
rect 22284 3884 22336 3893
rect 23204 3884 23256 3936
rect 24952 3884 25004 3936
rect 25964 3927 26016 3936
rect 25964 3893 25973 3927
rect 25973 3893 26007 3927
rect 26007 3893 26016 3927
rect 25964 3884 26016 3893
rect 27160 3927 27212 3936
rect 27160 3893 27169 3927
rect 27169 3893 27203 3927
rect 27203 3893 27212 3927
rect 27160 3884 27212 3893
rect 27896 3927 27948 3936
rect 27896 3893 27905 3927
rect 27905 3893 27939 3927
rect 27939 3893 27948 3927
rect 27896 3884 27948 3893
rect 27988 3884 28040 3936
rect 29828 4020 29880 4072
rect 46112 4020 46164 4072
rect 38568 3952 38620 4004
rect 41604 3952 41656 4004
rect 42432 3952 42484 4004
rect 47032 4097 47041 4131
rect 47041 4097 47075 4131
rect 47075 4097 47084 4131
rect 47032 4088 47084 4097
rect 48964 4088 49016 4140
rect 49424 4088 49476 4140
rect 49700 4088 49752 4140
rect 47584 4020 47636 4072
rect 51448 4156 51500 4208
rect 51356 4088 51408 4140
rect 52184 4088 52236 4140
rect 52460 4156 52512 4208
rect 53104 4088 53156 4140
rect 49332 3952 49384 4004
rect 51448 3952 51500 4004
rect 56324 4156 56376 4208
rect 55864 4131 55916 4140
rect 55864 4097 55873 4131
rect 55873 4097 55907 4131
rect 55907 4097 55916 4131
rect 55864 4088 55916 4097
rect 56600 4088 56652 4140
rect 57428 4088 57480 4140
rect 57152 4020 57204 4072
rect 56508 3952 56560 4004
rect 60464 4088 60516 4140
rect 60740 4088 60792 4140
rect 62212 4088 62264 4140
rect 63316 4131 63368 4140
rect 63316 4097 63325 4131
rect 63325 4097 63359 4131
rect 63359 4097 63368 4131
rect 63316 4088 63368 4097
rect 63868 4020 63920 4072
rect 59360 3952 59412 4004
rect 63960 3952 64012 4004
rect 66076 4156 66128 4208
rect 69296 4156 69348 4208
rect 79508 4156 79560 4208
rect 81348 4156 81400 4208
rect 66536 4131 66588 4140
rect 66536 4097 66545 4131
rect 66545 4097 66579 4131
rect 66579 4097 66588 4131
rect 66536 4088 66588 4097
rect 68836 4088 68888 4140
rect 71412 4088 71464 4140
rect 75736 4131 75788 4140
rect 75736 4097 75745 4131
rect 75745 4097 75779 4131
rect 75779 4097 75788 4131
rect 75736 4088 75788 4097
rect 78772 4088 78824 4140
rect 83096 4088 83148 4140
rect 83832 4131 83884 4140
rect 83832 4097 83841 4131
rect 83841 4097 83875 4131
rect 83875 4097 83884 4131
rect 83832 4088 83884 4097
rect 65156 4020 65208 4072
rect 69204 4020 69256 4072
rect 30288 3884 30340 3936
rect 31668 3927 31720 3936
rect 31668 3893 31677 3927
rect 31677 3893 31711 3927
rect 31711 3893 31720 3927
rect 31668 3884 31720 3893
rect 33324 3927 33376 3936
rect 33324 3893 33333 3927
rect 33333 3893 33367 3927
rect 33367 3893 33376 3927
rect 33324 3884 33376 3893
rect 33876 3927 33928 3936
rect 33876 3893 33885 3927
rect 33885 3893 33919 3927
rect 33919 3893 33928 3927
rect 33876 3884 33928 3893
rect 34244 3884 34296 3936
rect 37740 3884 37792 3936
rect 38752 3884 38804 3936
rect 39212 3927 39264 3936
rect 39212 3893 39221 3927
rect 39221 3893 39255 3927
rect 39255 3893 39264 3927
rect 39212 3884 39264 3893
rect 39948 3927 40000 3936
rect 39948 3893 39957 3927
rect 39957 3893 39991 3927
rect 39991 3893 40000 3927
rect 39948 3884 40000 3893
rect 41144 3884 41196 3936
rect 41880 3927 41932 3936
rect 41880 3893 41889 3927
rect 41889 3893 41923 3927
rect 41923 3893 41932 3927
rect 41880 3884 41932 3893
rect 42892 3884 42944 3936
rect 43904 3884 43956 3936
rect 45100 3927 45152 3936
rect 45100 3893 45109 3927
rect 45109 3893 45143 3927
rect 45143 3893 45152 3927
rect 45100 3884 45152 3893
rect 45468 3884 45520 3936
rect 46204 3927 46256 3936
rect 46204 3893 46213 3927
rect 46213 3893 46247 3927
rect 46247 3893 46256 3927
rect 46204 3884 46256 3893
rect 46296 3884 46348 3936
rect 46940 3884 46992 3936
rect 50620 3884 50672 3936
rect 50896 3927 50948 3936
rect 50896 3893 50905 3927
rect 50905 3893 50939 3927
rect 50939 3893 50948 3927
rect 50896 3884 50948 3893
rect 51540 3927 51592 3936
rect 51540 3893 51549 3927
rect 51549 3893 51583 3927
rect 51583 3893 51592 3927
rect 51540 3884 51592 3893
rect 52276 3927 52328 3936
rect 52276 3893 52285 3927
rect 52285 3893 52319 3927
rect 52319 3893 52328 3927
rect 52276 3884 52328 3893
rect 54024 3927 54076 3936
rect 54024 3893 54033 3927
rect 54033 3893 54067 3927
rect 54067 3893 54076 3927
rect 54024 3884 54076 3893
rect 55220 3927 55272 3936
rect 55220 3893 55229 3927
rect 55229 3893 55263 3927
rect 55263 3893 55272 3927
rect 55220 3884 55272 3893
rect 56600 3884 56652 3936
rect 59636 3884 59688 3936
rect 61384 3927 61436 3936
rect 61384 3893 61393 3927
rect 61393 3893 61427 3927
rect 61427 3893 61436 3927
rect 61384 3884 61436 3893
rect 63224 3884 63276 3936
rect 65340 3952 65392 4004
rect 67364 3952 67416 4004
rect 69756 4020 69808 4072
rect 72424 4020 72476 4072
rect 72516 4020 72568 4072
rect 79140 4063 79192 4072
rect 73528 3995 73580 4004
rect 65524 3927 65576 3936
rect 65524 3893 65533 3927
rect 65533 3893 65567 3927
rect 65567 3893 65576 3927
rect 65524 3884 65576 3893
rect 66536 3884 66588 3936
rect 68468 3884 68520 3936
rect 69204 3884 69256 3936
rect 73528 3961 73537 3995
rect 73537 3961 73571 3995
rect 73571 3961 73580 3995
rect 73528 3952 73580 3961
rect 77116 3995 77168 4004
rect 77116 3961 77125 3995
rect 77125 3961 77159 3995
rect 77159 3961 77168 3995
rect 77116 3952 77168 3961
rect 78680 3952 78732 4004
rect 71228 3884 71280 3936
rect 71596 3884 71648 3936
rect 75368 3884 75420 3936
rect 76472 3884 76524 3936
rect 78772 3884 78824 3936
rect 79140 4029 79149 4063
rect 79149 4029 79183 4063
rect 79183 4029 79192 4063
rect 79140 4020 79192 4029
rect 79784 4020 79836 4072
rect 81992 4063 82044 4072
rect 81992 4029 82001 4063
rect 82001 4029 82035 4063
rect 82035 4029 82044 4063
rect 81992 4020 82044 4029
rect 83004 4020 83056 4072
rect 83648 4020 83700 4072
rect 82728 3995 82780 4004
rect 82728 3961 82737 3995
rect 82737 3961 82771 3995
rect 82771 3961 82780 3995
rect 82728 3952 82780 3961
rect 81440 3884 81492 3936
rect 83464 3884 83516 3936
rect 117228 3884 117280 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 65654 3782 65706 3834
rect 65718 3782 65770 3834
rect 65782 3782 65834 3834
rect 65846 3782 65898 3834
rect 65910 3782 65962 3834
rect 96374 3782 96426 3834
rect 96438 3782 96490 3834
rect 96502 3782 96554 3834
rect 96566 3782 96618 3834
rect 96630 3782 96682 3834
rect 127094 3782 127146 3834
rect 127158 3782 127210 3834
rect 127222 3782 127274 3834
rect 127286 3782 127338 3834
rect 127350 3782 127402 3834
rect 22744 3723 22796 3732
rect 7012 3544 7064 3596
rect 5264 3476 5316 3528
rect 6276 3519 6328 3528
rect 6276 3485 6285 3519
rect 6285 3485 6319 3519
rect 6319 3485 6328 3519
rect 6276 3476 6328 3485
rect 6644 3476 6696 3528
rect 22744 3689 22753 3723
rect 22753 3689 22787 3723
rect 22787 3689 22796 3723
rect 22744 3680 22796 3689
rect 23940 3723 23992 3732
rect 23940 3689 23949 3723
rect 23949 3689 23983 3723
rect 23983 3689 23992 3723
rect 23940 3680 23992 3689
rect 24676 3723 24728 3732
rect 24676 3689 24685 3723
rect 24685 3689 24719 3723
rect 24719 3689 24728 3723
rect 24676 3680 24728 3689
rect 33140 3723 33192 3732
rect 27528 3612 27580 3664
rect 27988 3612 28040 3664
rect 28724 3612 28776 3664
rect 33140 3689 33149 3723
rect 33149 3689 33183 3723
rect 33183 3689 33192 3723
rect 33140 3680 33192 3689
rect 40224 3723 40276 3732
rect 40224 3689 40233 3723
rect 40233 3689 40267 3723
rect 40267 3689 40276 3723
rect 40224 3680 40276 3689
rect 40960 3723 41012 3732
rect 40960 3689 40969 3723
rect 40969 3689 41003 3723
rect 41003 3689 41012 3723
rect 40960 3680 41012 3689
rect 43812 3723 43864 3732
rect 43812 3689 43821 3723
rect 43821 3689 43855 3723
rect 43855 3689 43864 3723
rect 43812 3680 43864 3689
rect 46112 3680 46164 3732
rect 9404 3544 9456 3596
rect 22008 3544 22060 3596
rect 23296 3544 23348 3596
rect 24952 3544 25004 3596
rect 26240 3587 26292 3596
rect 26240 3553 26249 3587
rect 26249 3553 26283 3587
rect 26283 3553 26292 3587
rect 26240 3544 26292 3553
rect 27160 3544 27212 3596
rect 22100 3519 22152 3528
rect 5632 3408 5684 3460
rect 22100 3485 22109 3519
rect 22109 3485 22143 3519
rect 22143 3485 22152 3519
rect 22100 3476 22152 3485
rect 25872 3476 25924 3528
rect 27896 3544 27948 3596
rect 28080 3544 28132 3596
rect 30196 3544 30248 3596
rect 30380 3544 30432 3596
rect 35716 3587 35768 3596
rect 24216 3408 24268 3460
rect 5724 3340 5776 3392
rect 6736 3383 6788 3392
rect 6736 3349 6745 3383
rect 6745 3349 6779 3383
rect 6779 3349 6788 3383
rect 6736 3340 6788 3349
rect 7932 3383 7984 3392
rect 7932 3349 7941 3383
rect 7941 3349 7975 3383
rect 7975 3349 7984 3383
rect 7932 3340 7984 3349
rect 9220 3383 9272 3392
rect 9220 3349 9229 3383
rect 9229 3349 9263 3383
rect 9263 3349 9272 3383
rect 9220 3340 9272 3349
rect 20444 3383 20496 3392
rect 20444 3349 20453 3383
rect 20453 3349 20487 3383
rect 20487 3349 20496 3383
rect 20444 3340 20496 3349
rect 20996 3383 21048 3392
rect 20996 3349 21005 3383
rect 21005 3349 21039 3383
rect 21039 3349 21048 3383
rect 20996 3340 21048 3349
rect 21640 3383 21692 3392
rect 21640 3349 21649 3383
rect 21649 3349 21683 3383
rect 21683 3349 21692 3383
rect 21640 3340 21692 3349
rect 22744 3340 22796 3392
rect 23020 3340 23072 3392
rect 23940 3340 23992 3392
rect 24860 3340 24912 3392
rect 26424 3340 26476 3392
rect 27988 3383 28040 3392
rect 27988 3349 27997 3383
rect 27997 3349 28031 3383
rect 28031 3349 28040 3383
rect 32772 3476 32824 3528
rect 35716 3553 35725 3587
rect 35725 3553 35759 3587
rect 35759 3553 35768 3587
rect 35716 3544 35768 3553
rect 35992 3544 36044 3596
rect 38568 3612 38620 3664
rect 43352 3655 43404 3664
rect 43352 3621 43361 3655
rect 43361 3621 43395 3655
rect 43395 3621 43404 3655
rect 51356 3680 51408 3732
rect 53288 3680 53340 3732
rect 57428 3723 57480 3732
rect 53932 3655 53984 3664
rect 43352 3612 43404 3621
rect 41604 3587 41656 3596
rect 41604 3553 41613 3587
rect 41613 3553 41647 3587
rect 41647 3553 41656 3587
rect 41604 3544 41656 3553
rect 41880 3587 41932 3596
rect 41880 3553 41889 3587
rect 41889 3553 41923 3587
rect 41923 3553 41932 3587
rect 41880 3544 41932 3553
rect 43444 3544 43496 3596
rect 32864 3408 32916 3460
rect 37096 3476 37148 3528
rect 42984 3476 43036 3528
rect 27988 3340 28040 3349
rect 30748 3340 30800 3392
rect 32312 3340 32364 3392
rect 34704 3340 34756 3392
rect 35808 3408 35860 3460
rect 36084 3408 36136 3460
rect 38200 3451 38252 3460
rect 38200 3417 38209 3451
rect 38209 3417 38243 3451
rect 38243 3417 38252 3451
rect 38200 3408 38252 3417
rect 37096 3340 37148 3392
rect 38384 3340 38436 3392
rect 39764 3340 39816 3392
rect 41144 3408 41196 3460
rect 42524 3340 42576 3392
rect 45100 3476 45152 3528
rect 45928 3476 45980 3528
rect 46756 3476 46808 3528
rect 46848 3519 46900 3528
rect 46848 3485 46859 3519
rect 46859 3485 46893 3519
rect 46893 3485 46900 3519
rect 49056 3519 49108 3528
rect 46848 3476 46900 3485
rect 49056 3485 49065 3519
rect 49065 3485 49099 3519
rect 49099 3485 49108 3519
rect 49056 3476 49108 3485
rect 49332 3519 49384 3528
rect 49332 3485 49341 3519
rect 49341 3485 49375 3519
rect 49375 3485 49384 3519
rect 49332 3476 49384 3485
rect 44180 3451 44232 3460
rect 44180 3417 44189 3451
rect 44189 3417 44223 3451
rect 44223 3417 44232 3451
rect 44180 3408 44232 3417
rect 51908 3408 51960 3460
rect 45284 3383 45336 3392
rect 45284 3349 45293 3383
rect 45293 3349 45327 3383
rect 45327 3349 45336 3383
rect 45284 3340 45336 3349
rect 47676 3340 47728 3392
rect 47768 3340 47820 3392
rect 50620 3340 50672 3392
rect 50804 3340 50856 3392
rect 53932 3621 53941 3655
rect 53941 3621 53975 3655
rect 53975 3621 53984 3655
rect 53932 3612 53984 3621
rect 57428 3689 57437 3723
rect 57437 3689 57471 3723
rect 57471 3689 57480 3723
rect 57428 3680 57480 3689
rect 57704 3680 57756 3732
rect 52092 3544 52144 3596
rect 54208 3544 54260 3596
rect 52460 3476 52512 3528
rect 53012 3476 53064 3528
rect 53564 3408 53616 3460
rect 54300 3340 54352 3392
rect 54576 3340 54628 3392
rect 55864 3544 55916 3596
rect 55128 3476 55180 3528
rect 58624 3544 58676 3596
rect 61108 3587 61160 3596
rect 57152 3476 57204 3528
rect 61108 3553 61117 3587
rect 61117 3553 61151 3587
rect 61151 3553 61160 3587
rect 61108 3544 61160 3553
rect 62028 3519 62080 3528
rect 57704 3408 57756 3460
rect 57980 3408 58032 3460
rect 56048 3340 56100 3392
rect 56416 3340 56468 3392
rect 57428 3340 57480 3392
rect 57796 3383 57848 3392
rect 57796 3349 57805 3383
rect 57805 3349 57839 3383
rect 57839 3349 57848 3383
rect 57796 3340 57848 3349
rect 58716 3383 58768 3392
rect 58716 3349 58725 3383
rect 58725 3349 58759 3383
rect 58759 3349 58768 3383
rect 58716 3340 58768 3349
rect 59084 3340 59136 3392
rect 60004 3340 60056 3392
rect 61476 3408 61528 3460
rect 62028 3485 62037 3519
rect 62037 3485 62071 3519
rect 62071 3485 62080 3519
rect 62028 3476 62080 3485
rect 65064 3680 65116 3732
rect 66444 3680 66496 3732
rect 68836 3723 68888 3732
rect 62580 3544 62632 3596
rect 63500 3544 63552 3596
rect 63868 3587 63920 3596
rect 63868 3553 63877 3587
rect 63877 3553 63911 3587
rect 63911 3553 63920 3587
rect 63868 3544 63920 3553
rect 65432 3544 65484 3596
rect 66444 3587 66496 3596
rect 66444 3553 66453 3587
rect 66453 3553 66487 3587
rect 66487 3553 66496 3587
rect 66444 3544 66496 3553
rect 64880 3519 64932 3528
rect 64880 3485 64889 3519
rect 64889 3485 64923 3519
rect 64923 3485 64932 3519
rect 64880 3476 64932 3485
rect 66168 3476 66220 3528
rect 61200 3340 61252 3392
rect 62580 3340 62632 3392
rect 63500 3340 63552 3392
rect 65064 3408 65116 3460
rect 68836 3689 68845 3723
rect 68845 3689 68879 3723
rect 68879 3689 68888 3723
rect 68836 3680 68888 3689
rect 69848 3680 69900 3732
rect 70124 3680 70176 3732
rect 76472 3612 76524 3664
rect 80428 3680 80480 3732
rect 82084 3680 82136 3732
rect 82728 3680 82780 3732
rect 84844 3680 84896 3732
rect 145932 3680 145984 3732
rect 68008 3544 68060 3596
rect 68284 3587 68336 3596
rect 68284 3553 68293 3587
rect 68293 3553 68327 3587
rect 68327 3553 68336 3587
rect 68284 3544 68336 3553
rect 71412 3587 71464 3596
rect 71412 3553 71421 3587
rect 71421 3553 71455 3587
rect 71455 3553 71464 3587
rect 71412 3544 71464 3553
rect 71596 3587 71648 3596
rect 71596 3553 71605 3587
rect 71605 3553 71639 3587
rect 71639 3553 71648 3587
rect 71596 3544 71648 3553
rect 75368 3587 75420 3596
rect 75368 3553 75377 3587
rect 75377 3553 75411 3587
rect 75411 3553 75420 3587
rect 75368 3544 75420 3553
rect 77116 3544 77168 3596
rect 78772 3587 78824 3596
rect 78772 3553 78781 3587
rect 78781 3553 78815 3587
rect 78815 3553 78824 3587
rect 78772 3544 78824 3553
rect 80152 3544 80204 3596
rect 81348 3544 81400 3596
rect 81992 3544 82044 3596
rect 83280 3544 83332 3596
rect 104532 3612 104584 3664
rect 67640 3476 67692 3528
rect 68468 3519 68520 3528
rect 68468 3485 68477 3519
rect 68477 3485 68511 3519
rect 68511 3485 68520 3519
rect 68468 3476 68520 3485
rect 69112 3476 69164 3528
rect 69664 3519 69716 3528
rect 69664 3485 69673 3519
rect 69673 3485 69707 3519
rect 69707 3485 69716 3519
rect 69664 3476 69716 3485
rect 69940 3476 69992 3528
rect 70032 3476 70084 3528
rect 74080 3519 74132 3528
rect 74080 3485 74089 3519
rect 74089 3485 74123 3519
rect 74123 3485 74132 3519
rect 74080 3476 74132 3485
rect 74540 3476 74592 3528
rect 75736 3476 75788 3528
rect 75828 3476 75880 3528
rect 76564 3476 76616 3528
rect 69756 3408 69808 3460
rect 66812 3340 66864 3392
rect 67272 3383 67324 3392
rect 67272 3349 67281 3383
rect 67281 3349 67315 3383
rect 67315 3349 67324 3383
rect 67272 3340 67324 3349
rect 67364 3340 67416 3392
rect 70124 3408 70176 3460
rect 76196 3408 76248 3460
rect 69940 3340 69992 3392
rect 72700 3340 72752 3392
rect 72884 3340 72936 3392
rect 74448 3340 74500 3392
rect 75828 3340 75880 3392
rect 76380 3340 76432 3392
rect 78220 3476 78272 3528
rect 82820 3476 82872 3528
rect 83832 3476 83884 3528
rect 79416 3408 79468 3460
rect 81808 3408 81860 3460
rect 82360 3408 82412 3460
rect 108304 3408 108356 3460
rect 77668 3383 77720 3392
rect 77668 3349 77677 3383
rect 77677 3349 77711 3383
rect 77711 3349 77720 3383
rect 77668 3340 77720 3349
rect 78128 3340 78180 3392
rect 82728 3340 82780 3392
rect 83372 3340 83424 3392
rect 83648 3383 83700 3392
rect 83648 3349 83657 3383
rect 83657 3349 83691 3383
rect 83691 3349 83700 3383
rect 83648 3340 83700 3349
rect 85396 3383 85448 3392
rect 85396 3349 85405 3383
rect 85405 3349 85439 3383
rect 85439 3349 85448 3383
rect 85396 3340 85448 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 81014 3238 81066 3290
rect 81078 3238 81130 3290
rect 81142 3238 81194 3290
rect 81206 3238 81258 3290
rect 81270 3238 81322 3290
rect 111734 3238 111786 3290
rect 111798 3238 111850 3290
rect 111862 3238 111914 3290
rect 111926 3238 111978 3290
rect 111990 3238 112042 3290
rect 142454 3238 142506 3290
rect 142518 3238 142570 3290
rect 142582 3238 142634 3290
rect 142646 3238 142698 3290
rect 142710 3238 142762 3290
rect 5724 3179 5776 3188
rect 5724 3145 5733 3179
rect 5733 3145 5767 3179
rect 5767 3145 5776 3179
rect 5724 3136 5776 3145
rect 9404 3179 9456 3188
rect 9404 3145 9413 3179
rect 9413 3145 9447 3179
rect 9447 3145 9456 3179
rect 9404 3136 9456 3145
rect 21640 3136 21692 3188
rect 24216 3179 24268 3188
rect 4620 3068 4672 3120
rect 6000 3111 6052 3120
rect 6000 3077 6009 3111
rect 6009 3077 6043 3111
rect 6043 3077 6052 3111
rect 6000 3068 6052 3077
rect 6828 3068 6880 3120
rect 24216 3145 24225 3179
rect 24225 3145 24259 3179
rect 24259 3145 24268 3179
rect 24216 3136 24268 3145
rect 24676 3179 24728 3188
rect 24676 3145 24685 3179
rect 24685 3145 24719 3179
rect 24719 3145 24728 3179
rect 24676 3136 24728 3145
rect 6736 3043 6788 3052
rect 6736 3009 6745 3043
rect 6745 3009 6779 3043
rect 6779 3009 6788 3043
rect 6736 3000 6788 3009
rect 7012 3043 7064 3052
rect 7012 3009 7021 3043
rect 7021 3009 7055 3043
rect 7055 3009 7064 3043
rect 7012 3000 7064 3009
rect 8024 3000 8076 3052
rect 9404 3043 9456 3052
rect 9404 3009 9413 3043
rect 9413 3009 9447 3043
rect 9447 3009 9456 3043
rect 9404 3000 9456 3009
rect 20996 3000 21048 3052
rect 22100 3000 22152 3052
rect 23756 3043 23808 3052
rect 23756 3009 23765 3043
rect 23765 3009 23799 3043
rect 23799 3009 23808 3043
rect 23756 3000 23808 3009
rect 3884 2932 3936 2984
rect 21456 2932 21508 2984
rect 21916 2932 21968 2984
rect 24952 3136 25004 3188
rect 27344 3179 27396 3188
rect 27344 3145 27353 3179
rect 27353 3145 27387 3179
rect 27387 3145 27396 3179
rect 27344 3136 27396 3145
rect 27988 3136 28040 3188
rect 27528 3068 27580 3120
rect 28356 3068 28408 3120
rect 25872 3000 25924 3052
rect 26332 3000 26384 3052
rect 28816 3136 28868 3188
rect 30840 3179 30892 3188
rect 30840 3145 30849 3179
rect 30849 3145 30883 3179
rect 30883 3145 30892 3179
rect 30840 3136 30892 3145
rect 33784 3179 33836 3188
rect 28632 3068 28684 3120
rect 28908 3111 28960 3120
rect 28908 3077 28917 3111
rect 28917 3077 28951 3111
rect 28951 3077 28960 3111
rect 28908 3068 28960 3077
rect 29828 3111 29880 3120
rect 29828 3077 29837 3111
rect 29837 3077 29871 3111
rect 29871 3077 29880 3111
rect 29828 3068 29880 3077
rect 30104 3068 30156 3120
rect 30288 3068 30340 3120
rect 31484 3111 31536 3120
rect 31484 3077 31493 3111
rect 31493 3077 31527 3111
rect 31527 3077 31536 3111
rect 31484 3068 31536 3077
rect 31668 3111 31720 3120
rect 31668 3077 31677 3111
rect 31677 3077 31711 3111
rect 31711 3077 31720 3111
rect 31668 3068 31720 3077
rect 27620 2932 27672 2984
rect 33784 3145 33793 3179
rect 33793 3145 33827 3179
rect 33827 3145 33836 3179
rect 33784 3136 33836 3145
rect 34152 3179 34204 3188
rect 34152 3145 34161 3179
rect 34161 3145 34195 3179
rect 34195 3145 34204 3179
rect 34152 3136 34204 3145
rect 34428 3136 34480 3188
rect 37464 3179 37516 3188
rect 37464 3145 37473 3179
rect 37473 3145 37507 3179
rect 37507 3145 37516 3179
rect 37464 3136 37516 3145
rect 38108 3136 38160 3188
rect 46848 3136 46900 3188
rect 38200 3068 38252 3120
rect 39212 3111 39264 3120
rect 39212 3077 39221 3111
rect 39221 3077 39255 3111
rect 39255 3077 39264 3111
rect 39212 3068 39264 3077
rect 39948 3068 40000 3120
rect 41512 3068 41564 3120
rect 43352 3068 43404 3120
rect 46020 3068 46072 3120
rect 54024 3136 54076 3188
rect 57336 3179 57388 3188
rect 50896 3111 50948 3120
rect 50896 3077 50905 3111
rect 50905 3077 50939 3111
rect 50939 3077 50948 3111
rect 50896 3068 50948 3077
rect 51632 3068 51684 3120
rect 53288 3111 53340 3120
rect 53288 3077 53297 3111
rect 53297 3077 53331 3111
rect 53331 3077 53340 3111
rect 53288 3068 53340 3077
rect 53840 3068 53892 3120
rect 32772 3000 32824 3052
rect 33692 2932 33744 2984
rect 34796 2932 34848 2984
rect 35992 2932 36044 2984
rect 36912 2932 36964 2984
rect 38568 3000 38620 3052
rect 42524 3000 42576 3052
rect 42616 3000 42668 3052
rect 45468 3000 45520 3052
rect 39212 2932 39264 2984
rect 41420 2975 41472 2984
rect 41420 2941 41429 2975
rect 41429 2941 41463 2975
rect 41463 2941 41472 2975
rect 49332 3000 49384 3052
rect 50620 3043 50672 3052
rect 50620 3009 50629 3043
rect 50629 3009 50663 3043
rect 50663 3009 50672 3043
rect 50620 3000 50672 3009
rect 57336 3145 57345 3179
rect 57345 3145 57379 3179
rect 57379 3145 57388 3179
rect 57336 3136 57388 3145
rect 58716 3136 58768 3188
rect 54576 3111 54628 3120
rect 54576 3077 54585 3111
rect 54585 3077 54619 3111
rect 54619 3077 54628 3111
rect 54576 3068 54628 3077
rect 55220 3068 55272 3120
rect 57704 3068 57756 3120
rect 58072 3068 58124 3120
rect 58992 3068 59044 3120
rect 41420 2932 41472 2941
rect 5356 2796 5408 2848
rect 14924 2796 14976 2848
rect 20628 2796 20680 2848
rect 21824 2796 21876 2848
rect 26332 2796 26384 2848
rect 27896 2796 27948 2848
rect 41696 2864 41748 2916
rect 40684 2839 40736 2848
rect 40684 2805 40693 2839
rect 40693 2805 40727 2839
rect 40727 2805 40736 2839
rect 52460 2932 52512 2984
rect 54208 2932 54260 2984
rect 52184 2864 52236 2916
rect 40684 2796 40736 2805
rect 42156 2796 42208 2848
rect 42524 2796 42576 2848
rect 46664 2796 46716 2848
rect 50068 2839 50120 2848
rect 50068 2805 50077 2839
rect 50077 2805 50111 2839
rect 50111 2805 50120 2839
rect 50068 2796 50120 2805
rect 56508 3000 56560 3052
rect 59636 3000 59688 3052
rect 65156 3136 65208 3188
rect 60004 3111 60056 3120
rect 60004 3077 60013 3111
rect 60013 3077 60047 3111
rect 60047 3077 60056 3111
rect 60004 3068 60056 3077
rect 61384 3068 61436 3120
rect 62120 3068 62172 3120
rect 64052 3068 64104 3120
rect 64328 3068 64380 3120
rect 64604 3111 64656 3120
rect 64604 3077 64613 3111
rect 64613 3077 64647 3111
rect 64647 3077 64656 3111
rect 64604 3068 64656 3077
rect 64788 3111 64840 3120
rect 64788 3077 64797 3111
rect 64797 3077 64831 3111
rect 64831 3077 64840 3111
rect 64788 3068 64840 3077
rect 61844 3000 61896 3052
rect 63592 3043 63644 3052
rect 63592 3009 63601 3043
rect 63601 3009 63635 3043
rect 63635 3009 63644 3043
rect 66168 3136 66220 3188
rect 65524 3111 65576 3120
rect 65524 3077 65533 3111
rect 65533 3077 65567 3111
rect 65567 3077 65576 3111
rect 65524 3068 65576 3077
rect 67272 3068 67324 3120
rect 69296 3136 69348 3188
rect 69664 3136 69716 3188
rect 72516 3136 72568 3188
rect 73712 3179 73764 3188
rect 73712 3145 73721 3179
rect 73721 3145 73755 3179
rect 73755 3145 73764 3179
rect 73712 3136 73764 3145
rect 77208 3179 77260 3188
rect 77208 3145 77217 3179
rect 77217 3145 77251 3179
rect 77251 3145 77260 3179
rect 77208 3136 77260 3145
rect 79784 3136 79836 3188
rect 81716 3179 81768 3188
rect 81716 3145 81725 3179
rect 81725 3145 81759 3179
rect 81759 3145 81768 3179
rect 81716 3136 81768 3145
rect 82360 3136 82412 3188
rect 83188 3136 83240 3188
rect 83372 3136 83424 3188
rect 84108 3136 84160 3188
rect 125508 3136 125560 3188
rect 145932 3179 145984 3188
rect 145932 3145 145941 3179
rect 145941 3145 145975 3179
rect 145975 3145 145984 3179
rect 145932 3136 145984 3145
rect 69848 3068 69900 3120
rect 70400 3111 70452 3120
rect 70400 3077 70409 3111
rect 70409 3077 70443 3111
rect 70443 3077 70452 3111
rect 70400 3068 70452 3077
rect 70492 3068 70544 3120
rect 63592 3000 63644 3009
rect 58624 2975 58676 2984
rect 58624 2941 58633 2975
rect 58633 2941 58667 2975
rect 58667 2941 58676 2975
rect 58624 2932 58676 2941
rect 61476 2975 61528 2984
rect 61476 2941 61485 2975
rect 61485 2941 61519 2975
rect 61519 2941 61528 2975
rect 61476 2932 61528 2941
rect 63868 2975 63920 2984
rect 63868 2941 63877 2975
rect 63877 2941 63911 2975
rect 63911 2941 63920 2975
rect 63868 2932 63920 2941
rect 58164 2864 58216 2916
rect 62028 2864 62080 2916
rect 55680 2796 55732 2848
rect 56048 2839 56100 2848
rect 56048 2805 56057 2839
rect 56057 2805 56091 2839
rect 56091 2805 56100 2839
rect 56048 2796 56100 2805
rect 56692 2839 56744 2848
rect 56692 2805 56701 2839
rect 56701 2805 56735 2839
rect 56735 2805 56744 2839
rect 56692 2796 56744 2805
rect 66812 3000 66864 3052
rect 68008 3000 68060 3052
rect 68836 3043 68888 3052
rect 68836 3009 68845 3043
rect 68845 3009 68879 3043
rect 68879 3009 68888 3043
rect 68836 3000 68888 3009
rect 69756 3000 69808 3052
rect 72424 3043 72476 3052
rect 65064 2932 65116 2984
rect 69940 2932 69992 2984
rect 72424 3009 72433 3043
rect 72433 3009 72467 3043
rect 72467 3009 72476 3043
rect 72424 3000 72476 3009
rect 72884 3000 72936 3052
rect 74448 3043 74500 3052
rect 74448 3009 74457 3043
rect 74457 3009 74491 3043
rect 74491 3009 74500 3043
rect 74448 3000 74500 3009
rect 75092 3043 75144 3052
rect 75092 3009 75101 3043
rect 75101 3009 75135 3043
rect 75135 3009 75144 3043
rect 75092 3000 75144 3009
rect 75736 3043 75788 3052
rect 75736 3009 75745 3043
rect 75745 3009 75779 3043
rect 75779 3009 75788 3043
rect 75736 3000 75788 3009
rect 77024 3000 77076 3052
rect 82820 3068 82872 3120
rect 137284 3068 137336 3120
rect 74080 2932 74132 2984
rect 76196 2932 76248 2984
rect 83280 3000 83332 3052
rect 84200 3000 84252 3052
rect 84936 3000 84988 3052
rect 85396 3000 85448 3052
rect 104532 3043 104584 3052
rect 104532 3009 104541 3043
rect 104541 3009 104575 3043
rect 104575 3009 104584 3043
rect 104532 3000 104584 3009
rect 78680 2932 78732 2984
rect 79140 2932 79192 2984
rect 80244 2932 80296 2984
rect 81992 2932 82044 2984
rect 83648 2932 83700 2984
rect 70032 2864 70084 2916
rect 70124 2864 70176 2916
rect 71504 2864 71556 2916
rect 76840 2864 76892 2916
rect 67272 2796 67324 2848
rect 67364 2796 67416 2848
rect 71136 2796 71188 2848
rect 73804 2796 73856 2848
rect 75644 2796 75696 2848
rect 76472 2839 76524 2848
rect 76472 2805 76481 2839
rect 76481 2805 76515 2839
rect 76515 2805 76524 2839
rect 76472 2796 76524 2805
rect 76564 2796 76616 2848
rect 84844 2864 84896 2916
rect 83188 2796 83240 2848
rect 85672 2839 85724 2848
rect 85672 2805 85681 2839
rect 85681 2805 85715 2839
rect 85715 2805 85724 2839
rect 85672 2796 85724 2805
rect 97724 2839 97776 2848
rect 97724 2805 97733 2839
rect 97733 2805 97767 2839
rect 97767 2805 97776 2839
rect 97724 2796 97776 2805
rect 101864 2839 101916 2848
rect 101864 2805 101873 2839
rect 101873 2805 101907 2839
rect 101907 2805 101916 2839
rect 101864 2796 101916 2805
rect 110420 2796 110472 2848
rect 118424 2839 118476 2848
rect 118424 2805 118433 2839
rect 118433 2805 118467 2839
rect 118467 2805 118476 2839
rect 118424 2796 118476 2805
rect 122564 2839 122616 2848
rect 122564 2805 122573 2839
rect 122573 2805 122607 2839
rect 122607 2805 122616 2839
rect 122564 2796 122616 2805
rect 125416 2796 125468 2848
rect 130844 2839 130896 2848
rect 130844 2805 130853 2839
rect 130853 2805 130887 2839
rect 130887 2805 130896 2839
rect 130844 2796 130896 2805
rect 143264 2839 143316 2848
rect 143264 2805 143273 2839
rect 143273 2805 143307 2839
rect 143307 2805 143316 2839
rect 143264 2796 143316 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 65654 2694 65706 2746
rect 65718 2694 65770 2746
rect 65782 2694 65834 2746
rect 65846 2694 65898 2746
rect 65910 2694 65962 2746
rect 96374 2694 96426 2746
rect 96438 2694 96490 2746
rect 96502 2694 96554 2746
rect 96566 2694 96618 2746
rect 96630 2694 96682 2746
rect 127094 2694 127146 2746
rect 127158 2694 127210 2746
rect 127222 2694 127274 2746
rect 127286 2694 127338 2746
rect 127350 2694 127402 2746
rect 4620 2592 4672 2644
rect 9404 2592 9456 2644
rect 14464 2635 14516 2644
rect 14464 2601 14473 2635
rect 14473 2601 14507 2635
rect 14507 2601 14516 2635
rect 14464 2592 14516 2601
rect 15384 2635 15436 2644
rect 15384 2601 15393 2635
rect 15393 2601 15427 2635
rect 15427 2601 15436 2635
rect 15384 2592 15436 2601
rect 21272 2635 21324 2644
rect 21272 2601 21281 2635
rect 21281 2601 21315 2635
rect 21315 2601 21324 2635
rect 21272 2592 21324 2601
rect 24768 2635 24820 2644
rect 24768 2601 24777 2635
rect 24777 2601 24811 2635
rect 24811 2601 24820 2635
rect 24768 2592 24820 2601
rect 25688 2635 25740 2644
rect 25688 2601 25697 2635
rect 25697 2601 25731 2635
rect 25731 2601 25740 2635
rect 25688 2592 25740 2601
rect 26516 2635 26568 2644
rect 26516 2601 26525 2635
rect 26525 2601 26559 2635
rect 26559 2601 26568 2635
rect 26516 2592 26568 2601
rect 28908 2635 28960 2644
rect 28908 2601 28917 2635
rect 28917 2601 28951 2635
rect 28951 2601 28960 2635
rect 28908 2592 28960 2601
rect 34152 2592 34204 2644
rect 37096 2592 37148 2644
rect 39212 2635 39264 2644
rect 39212 2601 39221 2635
rect 39221 2601 39255 2635
rect 39255 2601 39264 2635
rect 39212 2592 39264 2601
rect 40040 2635 40092 2644
rect 40040 2601 40049 2635
rect 40049 2601 40083 2635
rect 40083 2601 40092 2635
rect 40040 2592 40092 2601
rect 41512 2592 41564 2644
rect 44180 2592 44232 2644
rect 47216 2635 47268 2644
rect 47216 2601 47225 2635
rect 47225 2601 47259 2635
rect 47259 2601 47268 2635
rect 47216 2592 47268 2601
rect 49516 2635 49568 2644
rect 49516 2601 49525 2635
rect 49525 2601 49559 2635
rect 49559 2601 49568 2635
rect 49516 2592 49568 2601
rect 50620 2592 50672 2644
rect 60832 2592 60884 2644
rect 19984 2524 20036 2576
rect 20720 2567 20772 2576
rect 20720 2533 20729 2567
rect 20729 2533 20763 2567
rect 20763 2533 20772 2567
rect 20720 2524 20772 2533
rect 6368 2456 6420 2508
rect 9220 2456 9272 2508
rect 23848 2456 23900 2508
rect 26240 2456 26292 2508
rect 32312 2499 32364 2508
rect 32312 2465 32321 2499
rect 32321 2465 32355 2499
rect 32355 2465 32364 2499
rect 32312 2456 32364 2465
rect 34796 2456 34848 2508
rect 38476 2456 38528 2508
rect 41420 2456 41472 2508
rect 7932 2388 7984 2440
rect 9404 2388 9456 2440
rect 5632 2320 5684 2372
rect 6828 2363 6880 2372
rect 2504 2252 2556 2304
rect 5356 2252 5408 2304
rect 6828 2329 6837 2363
rect 6837 2329 6871 2363
rect 6871 2329 6880 2363
rect 6828 2320 6880 2329
rect 8576 2363 8628 2372
rect 8576 2329 8585 2363
rect 8585 2329 8619 2363
rect 8619 2329 8628 2363
rect 8576 2320 8628 2329
rect 12164 2252 12216 2304
rect 13544 2252 13596 2304
rect 14924 2388 14976 2440
rect 20628 2388 20680 2440
rect 21456 2431 21508 2440
rect 21456 2397 21465 2431
rect 21465 2397 21499 2431
rect 21499 2397 21508 2431
rect 21456 2388 21508 2397
rect 21824 2388 21876 2440
rect 26332 2388 26384 2440
rect 30288 2431 30340 2440
rect 19432 2320 19484 2372
rect 17684 2252 17736 2304
rect 19064 2252 19116 2304
rect 19616 2320 19668 2372
rect 20444 2320 20496 2372
rect 22284 2363 22336 2372
rect 22284 2329 22293 2363
rect 22293 2329 22327 2363
rect 22327 2329 22336 2363
rect 22284 2320 22336 2329
rect 22744 2320 22796 2372
rect 24860 2363 24912 2372
rect 24860 2329 24869 2363
rect 24869 2329 24903 2363
rect 24903 2329 24912 2363
rect 24860 2320 24912 2329
rect 25964 2320 26016 2372
rect 26424 2363 26476 2372
rect 26424 2329 26433 2363
rect 26433 2329 26467 2363
rect 26467 2329 26476 2363
rect 26424 2320 26476 2329
rect 30288 2397 30297 2431
rect 30297 2397 30331 2431
rect 30331 2397 30340 2431
rect 30288 2388 30340 2397
rect 31760 2431 31812 2440
rect 31760 2397 31769 2431
rect 31769 2397 31803 2431
rect 31803 2397 31812 2431
rect 31760 2388 31812 2397
rect 40684 2388 40736 2440
rect 42616 2499 42668 2508
rect 42616 2465 42625 2499
rect 42625 2465 42659 2499
rect 42659 2465 42668 2499
rect 42616 2456 42668 2465
rect 46296 2456 46348 2508
rect 47768 2499 47820 2508
rect 47768 2465 47777 2499
rect 47777 2465 47811 2499
rect 47811 2465 47820 2499
rect 47768 2456 47820 2465
rect 53288 2524 53340 2576
rect 54944 2524 54996 2576
rect 51540 2456 51592 2508
rect 51908 2456 51960 2508
rect 54208 2499 54260 2508
rect 54208 2465 54217 2499
rect 54217 2465 54251 2499
rect 54251 2465 54260 2499
rect 54208 2456 54260 2465
rect 55128 2456 55180 2508
rect 55680 2499 55732 2508
rect 55680 2465 55689 2499
rect 55689 2465 55723 2499
rect 55723 2465 55732 2499
rect 55680 2456 55732 2465
rect 58716 2456 58768 2508
rect 63592 2592 63644 2644
rect 65064 2592 65116 2644
rect 69020 2635 69072 2644
rect 69020 2601 69029 2635
rect 69029 2601 69063 2635
rect 69063 2601 69072 2635
rect 69020 2592 69072 2601
rect 69112 2592 69164 2644
rect 70124 2592 70176 2644
rect 70952 2592 71004 2644
rect 68836 2524 68888 2576
rect 69112 2456 69164 2508
rect 54300 2388 54352 2440
rect 62304 2388 62356 2440
rect 70492 2524 70544 2576
rect 70952 2499 71004 2508
rect 70952 2465 70961 2499
rect 70961 2465 70995 2499
rect 70995 2465 71004 2499
rect 73528 2499 73580 2508
rect 70952 2456 71004 2465
rect 73528 2465 73537 2499
rect 73537 2465 73571 2499
rect 73571 2465 73580 2499
rect 73528 2456 73580 2465
rect 76472 2456 76524 2508
rect 78680 2499 78732 2508
rect 78680 2465 78689 2499
rect 78689 2465 78723 2499
rect 78723 2465 78732 2499
rect 78680 2456 78732 2465
rect 80244 2456 80296 2508
rect 81348 2592 81400 2644
rect 85488 2635 85540 2644
rect 82912 2524 82964 2576
rect 84108 2524 84160 2576
rect 84200 2456 84252 2508
rect 27896 2320 27948 2372
rect 30748 2320 30800 2372
rect 23112 2252 23164 2304
rect 27344 2252 27396 2304
rect 33324 2320 33376 2372
rect 34704 2320 34756 2372
rect 35900 2320 35952 2372
rect 37740 2363 37792 2372
rect 37740 2329 37749 2363
rect 37749 2329 37783 2363
rect 37783 2329 37792 2363
rect 37740 2320 37792 2329
rect 38752 2320 38804 2372
rect 40592 2320 40644 2372
rect 42892 2363 42944 2372
rect 42892 2329 42901 2363
rect 42901 2329 42935 2363
rect 42935 2329 42944 2363
rect 42892 2320 42944 2329
rect 45284 2320 45336 2372
rect 46204 2320 46256 2372
rect 47676 2320 47728 2372
rect 50068 2320 50120 2372
rect 52276 2320 52328 2372
rect 33876 2252 33928 2304
rect 42524 2252 42576 2304
rect 56692 2320 56744 2372
rect 58348 2363 58400 2372
rect 58348 2329 58357 2363
rect 58357 2329 58391 2363
rect 58391 2329 58400 2363
rect 58348 2320 58400 2329
rect 59360 2320 59412 2372
rect 61200 2363 61252 2372
rect 61200 2329 61209 2363
rect 61209 2329 61243 2363
rect 61243 2329 61252 2363
rect 61200 2320 61252 2329
rect 63500 2363 63552 2372
rect 63500 2329 63509 2363
rect 63509 2329 63543 2363
rect 63543 2329 63552 2363
rect 63500 2320 63552 2329
rect 63960 2320 64012 2372
rect 65248 2320 65300 2372
rect 66536 2320 66588 2372
rect 56600 2252 56652 2304
rect 57428 2295 57480 2304
rect 57428 2261 57437 2295
rect 57437 2261 57471 2295
rect 57471 2261 57480 2295
rect 57428 2252 57480 2261
rect 59820 2295 59872 2304
rect 59820 2261 59829 2295
rect 59829 2261 59863 2295
rect 59863 2261 59872 2295
rect 59820 2252 59872 2261
rect 61476 2252 61528 2304
rect 68928 2363 68980 2372
rect 68928 2329 68937 2363
rect 68937 2329 68971 2363
rect 68971 2329 68980 2363
rect 68928 2320 68980 2329
rect 75828 2388 75880 2440
rect 80796 2388 80848 2440
rect 82820 2388 82872 2440
rect 67548 2295 67600 2304
rect 67548 2261 67557 2295
rect 67557 2261 67591 2295
rect 67591 2261 67600 2295
rect 67548 2252 67600 2261
rect 70952 2252 71004 2304
rect 71136 2320 71188 2372
rect 71688 2320 71740 2372
rect 73804 2363 73856 2372
rect 72700 2295 72752 2304
rect 72700 2261 72709 2295
rect 72709 2261 72743 2295
rect 72743 2261 72752 2295
rect 72700 2252 72752 2261
rect 73804 2329 73813 2363
rect 73813 2329 73847 2363
rect 73847 2329 73856 2363
rect 73804 2320 73856 2329
rect 74540 2320 74592 2372
rect 76380 2363 76432 2372
rect 76380 2329 76389 2363
rect 76389 2329 76423 2363
rect 76423 2329 76432 2363
rect 76380 2320 76432 2329
rect 76840 2320 76892 2372
rect 78128 2363 78180 2372
rect 78128 2329 78137 2363
rect 78137 2329 78171 2363
rect 78171 2329 78180 2363
rect 78128 2320 78180 2329
rect 81348 2252 81400 2304
rect 81624 2320 81676 2372
rect 83096 2320 83148 2372
rect 85488 2601 85497 2635
rect 85497 2601 85531 2635
rect 85531 2601 85540 2635
rect 85488 2592 85540 2601
rect 89720 2635 89772 2644
rect 89720 2601 89729 2635
rect 89729 2601 89763 2635
rect 89763 2601 89772 2635
rect 89720 2592 89772 2601
rect 94320 2635 94372 2644
rect 94320 2601 94329 2635
rect 94329 2601 94363 2635
rect 94363 2601 94372 2635
rect 94320 2592 94372 2601
rect 97816 2592 97868 2644
rect 102140 2635 102192 2644
rect 102140 2601 102149 2635
rect 102149 2601 102183 2635
rect 102183 2601 102192 2635
rect 102140 2592 102192 2601
rect 106280 2635 106332 2644
rect 106280 2601 106289 2635
rect 106289 2601 106323 2635
rect 106323 2601 106332 2635
rect 106280 2592 106332 2601
rect 110512 2635 110564 2644
rect 110512 2601 110521 2635
rect 110521 2601 110555 2635
rect 110555 2601 110564 2635
rect 110512 2592 110564 2601
rect 114836 2592 114888 2644
rect 118700 2635 118752 2644
rect 118700 2601 118709 2635
rect 118709 2601 118743 2635
rect 118743 2601 118752 2635
rect 118700 2592 118752 2601
rect 122840 2635 122892 2644
rect 122840 2601 122849 2635
rect 122849 2601 122883 2635
rect 122883 2601 122892 2635
rect 126980 2635 127032 2644
rect 122840 2592 122892 2601
rect 126980 2601 126989 2635
rect 126989 2601 127023 2635
rect 127023 2601 127032 2635
rect 126980 2592 127032 2601
rect 131120 2635 131172 2644
rect 131120 2601 131129 2635
rect 131129 2601 131163 2635
rect 131163 2601 131172 2635
rect 131120 2592 131172 2601
rect 137284 2635 137336 2644
rect 137284 2601 137293 2635
rect 137293 2601 137327 2635
rect 137327 2601 137336 2635
rect 137284 2592 137336 2601
rect 141332 2592 141384 2644
rect 143540 2635 143592 2644
rect 143540 2601 143549 2635
rect 143549 2601 143583 2635
rect 143583 2601 143592 2635
rect 143540 2592 143592 2601
rect 147312 2635 147364 2644
rect 147312 2601 147321 2635
rect 147321 2601 147355 2635
rect 147355 2601 147364 2635
rect 147312 2592 147364 2601
rect 108764 2524 108816 2576
rect 117228 2524 117280 2576
rect 108304 2456 108356 2508
rect 84936 2431 84988 2440
rect 84936 2397 84945 2431
rect 84945 2397 84979 2431
rect 84979 2397 84988 2431
rect 84936 2388 84988 2397
rect 85304 2320 85356 2372
rect 89444 2320 89496 2372
rect 82820 2252 82872 2304
rect 83004 2295 83056 2304
rect 83004 2261 83013 2295
rect 83013 2261 83047 2295
rect 83047 2261 83056 2295
rect 83004 2252 83056 2261
rect 83924 2252 83976 2304
rect 84200 2252 84252 2304
rect 85672 2252 85724 2304
rect 87604 2295 87656 2304
rect 87604 2261 87613 2295
rect 87613 2261 87647 2295
rect 87647 2261 87656 2295
rect 87604 2252 87656 2261
rect 88064 2252 88116 2304
rect 91744 2295 91796 2304
rect 91744 2261 91753 2295
rect 91753 2261 91787 2295
rect 91787 2261 91796 2295
rect 91744 2252 91796 2261
rect 92204 2252 92256 2304
rect 93584 2295 93636 2304
rect 93584 2261 93593 2295
rect 93593 2261 93627 2295
rect 93627 2261 93636 2295
rect 97724 2320 97776 2372
rect 104532 2388 104584 2440
rect 101864 2320 101916 2372
rect 106004 2320 106056 2372
rect 110420 2363 110472 2372
rect 110420 2329 110429 2363
rect 110429 2329 110463 2363
rect 110463 2329 110472 2363
rect 110420 2320 110472 2329
rect 96068 2295 96120 2304
rect 93584 2252 93636 2261
rect 96068 2261 96077 2295
rect 96077 2261 96111 2295
rect 96111 2261 96120 2295
rect 96068 2252 96120 2261
rect 96344 2252 96396 2304
rect 100024 2295 100076 2304
rect 100024 2261 100033 2295
rect 100033 2261 100067 2295
rect 100067 2261 100076 2295
rect 100024 2252 100076 2261
rect 100484 2252 100536 2304
rect 104624 2252 104676 2304
rect 109040 2295 109092 2304
rect 109040 2261 109049 2295
rect 109049 2261 109083 2295
rect 109083 2261 109092 2295
rect 109040 2252 109092 2261
rect 112444 2295 112496 2304
rect 112444 2261 112453 2295
rect 112453 2261 112487 2295
rect 112487 2261 112496 2295
rect 112444 2252 112496 2261
rect 112904 2252 112956 2304
rect 114284 2252 114336 2304
rect 125416 2431 125468 2440
rect 125416 2397 125425 2431
rect 125425 2397 125459 2431
rect 125459 2397 125468 2431
rect 125416 2388 125468 2397
rect 125508 2388 125560 2440
rect 139492 2524 139544 2576
rect 118424 2320 118476 2372
rect 122564 2320 122616 2372
rect 126704 2320 126756 2372
rect 130844 2320 130896 2372
rect 137284 2388 137336 2440
rect 139124 2388 139176 2440
rect 145932 2388 145984 2440
rect 143264 2320 143316 2372
rect 147404 2320 147456 2372
rect 116676 2295 116728 2304
rect 116676 2261 116685 2295
rect 116685 2261 116719 2295
rect 116719 2261 116728 2295
rect 116676 2252 116728 2261
rect 117044 2252 117096 2304
rect 121184 2252 121236 2304
rect 125324 2252 125376 2304
rect 129648 2252 129700 2304
rect 133604 2252 133656 2304
rect 134984 2252 135036 2304
rect 137744 2252 137796 2304
rect 141424 2295 141476 2304
rect 141424 2261 141433 2295
rect 141433 2261 141467 2295
rect 141467 2261 141476 2295
rect 141424 2252 141476 2261
rect 141884 2252 141936 2304
rect 146024 2252 146076 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 81014 2150 81066 2202
rect 81078 2150 81130 2202
rect 81142 2150 81194 2202
rect 81206 2150 81258 2202
rect 81270 2150 81322 2202
rect 111734 2150 111786 2202
rect 111798 2150 111850 2202
rect 111862 2150 111914 2202
rect 111926 2150 111978 2202
rect 111990 2150 112042 2202
rect 142454 2150 142506 2202
rect 142518 2150 142570 2202
rect 142582 2150 142634 2202
rect 142646 2150 142698 2202
rect 142710 2150 142762 2202
rect 8576 2048 8628 2100
rect 23296 2048 23348 2100
rect 57428 2048 57480 2100
rect 96068 2048 96120 2100
rect 56048 1980 56100 2032
rect 91744 1980 91796 2032
rect 64880 1912 64932 1964
rect 67548 1912 67600 1964
rect 100024 1912 100076 1964
rect 70952 1844 71004 1896
rect 71688 1844 71740 1896
rect 81164 1844 81216 1896
rect 83280 1844 83332 1896
rect 72700 1776 72752 1828
rect 116676 1776 116728 1828
rect 71228 1708 71280 1760
rect 109040 1708 109092 1760
rect 78128 1640 78180 1692
rect 141424 1640 141476 1692
rect 59820 1572 59872 1624
rect 87604 1572 87656 1624
rect 83004 1504 83056 1556
rect 125416 1504 125468 1556
rect 81440 1436 81492 1488
rect 112444 1436 112496 1488
<< metal2 >>
rect 2686 39200 2742 40000
rect 3606 39200 3662 40000
rect 4526 39200 4582 40000
rect 5446 39200 5502 40000
rect 6366 39200 6422 40000
rect 7286 39200 7342 40000
rect 8206 39200 8262 40000
rect 9126 39200 9182 40000
rect 10046 39200 10102 40000
rect 10966 39200 11022 40000
rect 11886 39200 11942 40000
rect 12806 39200 12862 40000
rect 13726 39200 13782 40000
rect 14646 39200 14702 40000
rect 15566 39200 15622 40000
rect 16486 39200 16542 40000
rect 17406 39200 17462 40000
rect 18326 39200 18382 40000
rect 19246 39200 19302 40000
rect 20166 39200 20222 40000
rect 21086 39200 21142 40000
rect 22006 39200 22062 40000
rect 22926 39200 22982 40000
rect 23846 39200 23902 40000
rect 24766 39200 24822 40000
rect 25686 39200 25742 40000
rect 26606 39200 26662 40000
rect 27526 39200 27582 40000
rect 28446 39200 28502 40000
rect 29366 39200 29422 40000
rect 30286 39200 30342 40000
rect 31206 39200 31262 40000
rect 32126 39200 32182 40000
rect 33046 39200 33102 40000
rect 33966 39200 34022 40000
rect 34532 39222 34836 39250
rect 2700 38298 2728 39200
rect 2700 38270 2820 38298
rect 2792 37466 2820 38270
rect 2780 37460 2832 37466
rect 2780 37402 2832 37408
rect 3620 36922 3648 39200
rect 4540 37754 4568 39200
rect 4540 37726 4660 37754
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4528 37392 4580 37398
rect 4528 37334 4580 37340
rect 4540 36922 4568 37334
rect 4632 37126 4660 37726
rect 4896 37256 4948 37262
rect 4896 37198 4948 37204
rect 4620 37120 4672 37126
rect 4620 37062 4672 37068
rect 3608 36916 3660 36922
rect 3608 36858 3660 36864
rect 4528 36916 4580 36922
rect 4528 36858 4580 36864
rect 4908 36854 4936 37198
rect 5460 37108 5488 39200
rect 5540 37120 5592 37126
rect 5460 37080 5540 37108
rect 5540 37062 5592 37068
rect 4896 36848 4948 36854
rect 4896 36790 4948 36796
rect 6380 36786 6408 39200
rect 6920 37256 6972 37262
rect 6920 37198 6972 37204
rect 6368 36780 6420 36786
rect 6368 36722 6420 36728
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 6932 36106 6960 37198
rect 7300 37126 7328 39200
rect 8220 37346 8248 39200
rect 8220 37318 8340 37346
rect 8208 37256 8260 37262
rect 8208 37198 8260 37204
rect 7288 37120 7340 37126
rect 7288 37062 7340 37068
rect 8220 36922 8248 37198
rect 8312 37126 8340 37318
rect 8576 37256 8628 37262
rect 8576 37198 8628 37204
rect 8300 37120 8352 37126
rect 8300 37062 8352 37068
rect 8208 36916 8260 36922
rect 8208 36858 8260 36864
rect 8392 36780 8444 36786
rect 8392 36722 8444 36728
rect 8404 36582 8432 36722
rect 8392 36576 8444 36582
rect 8392 36518 8444 36524
rect 6920 36100 6972 36106
rect 6920 36042 6972 36048
rect 8588 36038 8616 37198
rect 9140 37126 9168 39200
rect 10060 37262 10088 39200
rect 9772 37256 9824 37262
rect 9772 37198 9824 37204
rect 10048 37256 10100 37262
rect 10048 37198 10100 37204
rect 9128 37120 9180 37126
rect 9128 37062 9180 37068
rect 9784 36922 9812 37198
rect 9772 36916 9824 36922
rect 9772 36858 9824 36864
rect 9588 36576 9640 36582
rect 9588 36518 9640 36524
rect 8576 36032 8628 36038
rect 8576 35974 8628 35980
rect 9600 35698 9628 36518
rect 10060 36378 10088 37198
rect 10980 37126 11008 39200
rect 11900 37126 11928 39200
rect 12256 37256 12308 37262
rect 12256 37198 12308 37204
rect 10324 37120 10376 37126
rect 10324 37062 10376 37068
rect 10968 37120 11020 37126
rect 10968 37062 11020 37068
rect 11888 37120 11940 37126
rect 11888 37062 11940 37068
rect 10048 36372 10100 36378
rect 10048 36314 10100 36320
rect 10336 36174 10364 37062
rect 12268 36922 12296 37198
rect 12820 37126 12848 39200
rect 13176 37256 13228 37262
rect 13176 37198 13228 37204
rect 12808 37120 12860 37126
rect 12808 37062 12860 37068
rect 12256 36916 12308 36922
rect 12256 36858 12308 36864
rect 13188 36854 13216 37198
rect 13740 36904 13768 39200
rect 14660 37126 14688 39200
rect 15580 37126 15608 39200
rect 15936 37256 15988 37262
rect 15936 37198 15988 37204
rect 14648 37120 14700 37126
rect 14648 37062 14700 37068
rect 15476 37120 15528 37126
rect 15476 37062 15528 37068
rect 15568 37120 15620 37126
rect 15568 37062 15620 37068
rect 13740 36876 13860 36904
rect 13176 36848 13228 36854
rect 13176 36790 13228 36796
rect 13832 36786 13860 36876
rect 10508 36780 10560 36786
rect 10508 36722 10560 36728
rect 13820 36780 13872 36786
rect 13820 36722 13872 36728
rect 10520 36582 10548 36722
rect 12898 36680 12954 36689
rect 12898 36615 12900 36624
rect 12952 36615 12954 36624
rect 12900 36586 12952 36592
rect 10508 36576 10560 36582
rect 10508 36518 10560 36524
rect 10520 36242 10548 36518
rect 10508 36236 10560 36242
rect 10508 36178 10560 36184
rect 14832 36236 14884 36242
rect 14832 36178 14884 36184
rect 10324 36168 10376 36174
rect 10324 36110 10376 36116
rect 14464 36100 14516 36106
rect 14464 36042 14516 36048
rect 9588 35692 9640 35698
rect 9588 35634 9640 35640
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 9600 12306 9628 35634
rect 9588 12300 9640 12306
rect 9588 12242 9640 12248
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 6368 4480 6420 4486
rect 6368 4422 6420 4428
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 4620 3120 4672 3126
rect 4620 3062 4672 3068
rect 3884 2984 3936 2990
rect 3884 2926 3936 2932
rect 2504 2304 2556 2310
rect 2504 2246 2556 2252
rect 2516 800 2544 2246
rect 3896 800 3924 2926
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2650 4660 3062
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 5276 800 5304 3470
rect 5632 3460 5684 3466
rect 5632 3402 5684 3408
rect 5356 2848 5408 2854
rect 5356 2790 5408 2796
rect 5368 2310 5396 2790
rect 5644 2378 5672 3402
rect 5724 3392 5776 3398
rect 5724 3334 5776 3340
rect 5736 3194 5764 3334
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 6012 3126 6040 4082
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 6288 3534 6316 3878
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 6000 3120 6052 3126
rect 6000 3062 6052 3068
rect 6380 2514 6408 4422
rect 6644 4004 6696 4010
rect 6644 3946 6696 3952
rect 6656 3534 6684 3946
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 6368 2508 6420 2514
rect 6368 2450 6420 2456
rect 5632 2372 5684 2378
rect 5632 2314 5684 2320
rect 5356 2304 5408 2310
rect 5356 2246 5408 2252
rect 6656 800 6684 3470
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 6748 3058 6776 3334
rect 6840 3126 6868 3878
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 6828 3120 6880 3126
rect 6828 3062 6880 3068
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6840 2378 6868 3062
rect 7024 3058 7052 3538
rect 7932 3392 7984 3398
rect 7932 3334 7984 3340
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 7944 2446 7972 3334
rect 8036 3058 8064 3878
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9220 3392 9272 3398
rect 9220 3334 9272 3340
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 6828 2372 6880 2378
rect 6828 2314 6880 2320
rect 8036 800 8064 2994
rect 9232 2514 9260 3334
rect 9416 3194 9444 3538
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9416 2650 9444 2994
rect 14476 2650 14504 36042
rect 14844 36038 14872 36178
rect 15488 36174 15516 37062
rect 15948 36582 15976 37198
rect 16500 37108 16528 39200
rect 17420 37262 17448 39200
rect 17316 37256 17368 37262
rect 17316 37198 17368 37204
rect 17408 37256 17460 37262
rect 17408 37198 17460 37204
rect 16580 37120 16632 37126
rect 16500 37080 16580 37108
rect 16580 37062 16632 37068
rect 17328 36922 17356 37198
rect 16580 36916 16632 36922
rect 16580 36858 16632 36864
rect 17316 36916 17368 36922
rect 17316 36858 17368 36864
rect 16592 36825 16620 36858
rect 16578 36816 16634 36825
rect 16578 36751 16634 36760
rect 15936 36576 15988 36582
rect 15936 36518 15988 36524
rect 17420 36378 17448 37198
rect 18340 37126 18368 39200
rect 19064 37256 19116 37262
rect 19064 37198 19116 37204
rect 17776 37120 17828 37126
rect 17776 37062 17828 37068
rect 18328 37120 18380 37126
rect 18328 37062 18380 37068
rect 17684 36576 17736 36582
rect 17684 36518 17736 36524
rect 17408 36372 17460 36378
rect 17408 36314 17460 36320
rect 15016 36168 15068 36174
rect 14936 36116 15016 36122
rect 15476 36168 15528 36174
rect 14936 36110 15068 36116
rect 15106 36136 15162 36145
rect 14936 36094 15056 36110
rect 15476 36110 15528 36116
rect 17696 36122 17724 36518
rect 17788 36378 17816 37062
rect 19076 36922 19104 37198
rect 19260 37108 19288 39200
rect 19432 37664 19484 37670
rect 19432 37606 19484 37612
rect 19340 37120 19392 37126
rect 19260 37080 19340 37108
rect 19340 37062 19392 37068
rect 19064 36916 19116 36922
rect 19064 36858 19116 36864
rect 19156 36916 19208 36922
rect 19156 36858 19208 36864
rect 19168 36786 19196 36858
rect 17960 36780 18012 36786
rect 17960 36722 18012 36728
rect 18052 36780 18104 36786
rect 18052 36722 18104 36728
rect 19156 36780 19208 36786
rect 19156 36722 19208 36728
rect 17972 36582 18000 36722
rect 18064 36650 18092 36722
rect 18052 36644 18104 36650
rect 18052 36586 18104 36592
rect 17960 36576 18012 36582
rect 17960 36518 18012 36524
rect 17776 36372 17828 36378
rect 17776 36314 17828 36320
rect 17972 36242 18000 36518
rect 17960 36236 18012 36242
rect 17960 36178 18012 36184
rect 14740 36032 14792 36038
rect 14740 35974 14792 35980
rect 14832 36032 14884 36038
rect 14832 35974 14884 35980
rect 14752 35850 14780 35974
rect 14936 35850 14964 36094
rect 17696 36094 18000 36122
rect 19444 36106 19472 37606
rect 19708 37256 19760 37262
rect 19706 37224 19708 37233
rect 19760 37224 19762 37233
rect 19706 37159 19762 37168
rect 19982 37224 20038 37233
rect 19982 37159 20038 37168
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19524 36712 19576 36718
rect 19524 36654 19576 36660
rect 19536 36174 19564 36654
rect 19524 36168 19576 36174
rect 19524 36110 19576 36116
rect 15106 36071 15108 36080
rect 15160 36071 15162 36080
rect 15108 36042 15160 36048
rect 14752 35822 14964 35850
rect 17972 35086 18000 36094
rect 19432 36100 19484 36106
rect 19432 36042 19484 36048
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19996 35834 20024 37159
rect 20180 37126 20208 39200
rect 20442 37496 20498 37505
rect 20442 37431 20498 37440
rect 20168 37120 20220 37126
rect 20168 37062 20220 37068
rect 20456 36922 20484 37431
rect 20548 37318 20760 37346
rect 20444 36916 20496 36922
rect 20444 36858 20496 36864
rect 20168 36712 20220 36718
rect 20168 36654 20220 36660
rect 20180 36174 20208 36654
rect 20260 36576 20312 36582
rect 20258 36544 20260 36553
rect 20312 36544 20314 36553
rect 20258 36479 20314 36488
rect 20168 36168 20220 36174
rect 20168 36110 20220 36116
rect 20548 36038 20576 37318
rect 20732 37262 20760 37318
rect 20628 37256 20680 37262
rect 20628 37198 20680 37204
rect 20720 37256 20772 37262
rect 20720 37198 20772 37204
rect 20640 36922 20668 37198
rect 20628 36916 20680 36922
rect 20628 36858 20680 36864
rect 20720 36780 20772 36786
rect 20720 36722 20772 36728
rect 20732 36106 20760 36722
rect 20812 36576 20864 36582
rect 20810 36544 20812 36553
rect 20864 36544 20866 36553
rect 20810 36479 20866 36488
rect 21100 36174 21128 39200
rect 21548 37188 21600 37194
rect 21548 37130 21600 37136
rect 21364 37120 21416 37126
rect 21364 37062 21416 37068
rect 21272 36780 21324 36786
rect 21272 36722 21324 36728
rect 21284 36281 21312 36722
rect 21270 36272 21326 36281
rect 21270 36207 21326 36216
rect 21088 36168 21140 36174
rect 21088 36110 21140 36116
rect 20720 36100 20772 36106
rect 20720 36042 20772 36048
rect 20536 36032 20588 36038
rect 20536 35974 20588 35980
rect 19984 35828 20036 35834
rect 19984 35770 20036 35776
rect 20548 35290 20576 35974
rect 19984 35284 20036 35290
rect 19984 35226 20036 35232
rect 20536 35284 20588 35290
rect 20536 35226 20588 35232
rect 17960 35080 18012 35086
rect 17960 35022 18012 35028
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 15384 12300 15436 12306
rect 15384 12242 15436 12248
rect 14924 2848 14976 2854
rect 14924 2790 14976 2796
rect 9404 2644 9456 2650
rect 9404 2586 9456 2592
rect 14464 2644 14516 2650
rect 14464 2586 14516 2592
rect 9220 2508 9272 2514
rect 9220 2450 9272 2456
rect 14936 2446 14964 2790
rect 15396 2650 15424 12242
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 19996 2582 20024 35226
rect 20444 3392 20496 3398
rect 20444 3334 20496 3340
rect 19984 2576 20036 2582
rect 19984 2518 20036 2524
rect 9404 2440 9456 2446
rect 9404 2382 9456 2388
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 8576 2372 8628 2378
rect 8576 2314 8628 2320
rect 8588 2106 8616 2314
rect 8576 2100 8628 2106
rect 8576 2042 8628 2048
rect 9416 800 9444 2382
rect 12164 2304 12216 2310
rect 12164 2246 12216 2252
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 12176 800 12204 2246
rect 13556 800 13584 2246
rect 14936 800 14964 2382
rect 20456 2378 20484 3334
rect 20628 2848 20680 2854
rect 20628 2790 20680 2796
rect 20640 2446 20668 2790
rect 20732 2582 20760 36042
rect 21100 35834 21128 36110
rect 21284 36038 21312 36207
rect 21272 36032 21324 36038
rect 21272 35974 21324 35980
rect 21088 35828 21140 35834
rect 21088 35770 21140 35776
rect 20996 3392 21048 3398
rect 20996 3334 21048 3340
rect 21008 3058 21036 3334
rect 20996 3052 21048 3058
rect 20996 2994 21048 3000
rect 21284 2650 21312 35974
rect 21376 33522 21404 37062
rect 21560 36854 21588 37130
rect 22020 37108 22048 39200
rect 22192 39160 22244 39166
rect 22192 39102 22244 39108
rect 22100 37120 22152 37126
rect 22020 37080 22100 37108
rect 22100 37062 22152 37068
rect 21548 36848 21600 36854
rect 21548 36790 21600 36796
rect 21824 36780 21876 36786
rect 21824 36722 21876 36728
rect 21732 36712 21784 36718
rect 21732 36654 21784 36660
rect 21744 36310 21772 36654
rect 21732 36304 21784 36310
rect 21732 36246 21784 36252
rect 21836 36174 21864 36722
rect 22204 36582 22232 39102
rect 22284 37256 22336 37262
rect 22282 37224 22284 37233
rect 22468 37256 22520 37262
rect 22336 37224 22338 37233
rect 22468 37198 22520 37204
rect 22282 37159 22338 37168
rect 22192 36576 22244 36582
rect 22192 36518 22244 36524
rect 22480 36378 22508 37198
rect 22940 37126 22968 39200
rect 23296 37256 23348 37262
rect 23296 37198 23348 37204
rect 23388 37256 23440 37262
rect 23388 37198 23440 37204
rect 22928 37120 22980 37126
rect 23308 37097 23336 37198
rect 22928 37062 22980 37068
rect 23294 37088 23350 37097
rect 23294 37023 23350 37032
rect 22744 36780 22796 36786
rect 22744 36722 22796 36728
rect 22756 36689 22784 36722
rect 23400 36689 23428 37198
rect 23860 36786 23888 39200
rect 24676 37256 24728 37262
rect 24676 37198 24728 37204
rect 23940 37188 23992 37194
rect 23940 37130 23992 37136
rect 23952 36854 23980 37130
rect 24032 37120 24084 37126
rect 24032 37062 24084 37068
rect 23940 36848 23992 36854
rect 23940 36790 23992 36796
rect 23480 36780 23532 36786
rect 23480 36722 23532 36728
rect 23848 36780 23900 36786
rect 23848 36722 23900 36728
rect 22742 36680 22798 36689
rect 22742 36615 22798 36624
rect 23386 36680 23442 36689
rect 23386 36615 23442 36624
rect 23492 36378 23520 36722
rect 23940 36576 23992 36582
rect 23940 36518 23992 36524
rect 22468 36372 22520 36378
rect 22468 36314 22520 36320
rect 23480 36372 23532 36378
rect 23480 36314 23532 36320
rect 23952 36242 23980 36518
rect 23940 36236 23992 36242
rect 23940 36178 23992 36184
rect 21824 36168 21876 36174
rect 21824 36110 21876 36116
rect 21364 33516 21416 33522
rect 21364 33458 21416 33464
rect 24044 26234 24072 37062
rect 24490 36952 24546 36961
rect 24490 36887 24546 36896
rect 24504 36854 24532 36887
rect 24688 36854 24716 37198
rect 24492 36848 24544 36854
rect 24492 36790 24544 36796
rect 24676 36848 24728 36854
rect 24676 36790 24728 36796
rect 24124 36780 24176 36786
rect 24124 36722 24176 36728
rect 24136 36378 24164 36722
rect 24124 36372 24176 36378
rect 24124 36314 24176 36320
rect 24504 35290 24532 36790
rect 24688 36666 24716 36790
rect 24596 36638 24716 36666
rect 24596 35494 24624 36638
rect 24676 36576 24728 36582
rect 24676 36518 24728 36524
rect 24584 35488 24636 35494
rect 24584 35430 24636 35436
rect 24492 35284 24544 35290
rect 24492 35226 24544 35232
rect 24596 34542 24624 35430
rect 24584 34536 24636 34542
rect 24584 34478 24636 34484
rect 23952 26206 24072 26234
rect 23296 4480 23348 4486
rect 23296 4422 23348 4428
rect 23848 4480 23900 4486
rect 23848 4422 23900 4428
rect 22744 4140 22796 4146
rect 22744 4082 22796 4088
rect 22284 3936 22336 3942
rect 22284 3878 22336 3884
rect 22006 3632 22062 3641
rect 22006 3567 22008 3576
rect 22060 3567 22062 3576
rect 22008 3538 22060 3544
rect 22100 3528 22152 3534
rect 22100 3470 22152 3476
rect 21640 3392 21692 3398
rect 21640 3334 21692 3340
rect 21652 3194 21680 3334
rect 21640 3188 21692 3194
rect 21640 3130 21692 3136
rect 22112 3058 22140 3470
rect 22100 3052 22152 3058
rect 22100 2994 22152 3000
rect 21456 2984 21508 2990
rect 21456 2926 21508 2932
rect 21916 2984 21968 2990
rect 21916 2926 21968 2932
rect 21272 2644 21324 2650
rect 21272 2586 21324 2592
rect 20720 2576 20772 2582
rect 20720 2518 20772 2524
rect 21468 2446 21496 2926
rect 21824 2848 21876 2854
rect 21928 2836 21956 2926
rect 21876 2808 21956 2836
rect 21824 2790 21876 2796
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 21456 2440 21508 2446
rect 21456 2382 21508 2388
rect 21824 2440 21876 2446
rect 21824 2382 21876 2388
rect 19432 2372 19484 2378
rect 19616 2372 19668 2378
rect 19484 2332 19616 2360
rect 19432 2314 19484 2320
rect 19616 2314 19668 2320
rect 20444 2372 20496 2378
rect 20444 2314 20496 2320
rect 17684 2304 17736 2310
rect 17684 2246 17736 2252
rect 19064 2304 19116 2310
rect 19064 2246 19116 2252
rect 17696 800 17724 2246
rect 19076 800 19104 2246
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 20456 800 20484 2314
rect 21836 800 21864 2382
rect 22296 2378 22324 3878
rect 22756 3738 22784 4082
rect 23204 3936 23256 3942
rect 23204 3878 23256 3884
rect 22744 3732 22796 3738
rect 22744 3674 22796 3680
rect 22744 3392 22796 3398
rect 22744 3334 22796 3340
rect 23020 3392 23072 3398
rect 23020 3334 23072 3340
rect 22756 2378 22784 3334
rect 23032 2774 23060 3334
rect 23032 2746 23152 2774
rect 22284 2372 22336 2378
rect 22284 2314 22336 2320
rect 22744 2372 22796 2378
rect 22744 2314 22796 2320
rect 23124 2310 23152 2746
rect 23112 2304 23164 2310
rect 23112 2246 23164 2252
rect 23216 800 23244 3878
rect 23308 3602 23336 4422
rect 23756 4004 23808 4010
rect 23756 3946 23808 3952
rect 23296 3596 23348 3602
rect 23296 3538 23348 3544
rect 23308 2106 23336 3538
rect 23768 3058 23796 3946
rect 23756 3052 23808 3058
rect 23756 2994 23808 3000
rect 23860 2514 23888 4422
rect 23952 3738 23980 26206
rect 24688 3738 24716 36518
rect 24780 36394 24808 39200
rect 25136 37664 25188 37670
rect 25136 37606 25188 37612
rect 25148 37330 25176 37606
rect 25136 37324 25188 37330
rect 25136 37266 25188 37272
rect 24858 37224 24914 37233
rect 24858 37159 24914 37168
rect 25044 37188 25096 37194
rect 24872 36582 24900 37159
rect 25044 37130 25096 37136
rect 25504 37188 25556 37194
rect 25504 37130 25556 37136
rect 25056 36718 25084 37130
rect 25136 37120 25188 37126
rect 25136 37062 25188 37068
rect 25320 37120 25372 37126
rect 25320 37062 25372 37068
rect 25044 36712 25096 36718
rect 25044 36654 25096 36660
rect 24860 36576 24912 36582
rect 24860 36518 24912 36524
rect 24780 36378 24900 36394
rect 24780 36372 24912 36378
rect 24780 36366 24860 36372
rect 24860 36314 24912 36320
rect 25148 36310 25176 37062
rect 25332 36786 25360 37062
rect 25320 36780 25372 36786
rect 25320 36722 25372 36728
rect 25136 36304 25188 36310
rect 25188 36252 25268 36258
rect 25136 36246 25268 36252
rect 25148 36230 25268 36246
rect 25136 36168 25188 36174
rect 25136 36110 25188 36116
rect 25148 35834 25176 36110
rect 25136 35828 25188 35834
rect 25136 35770 25188 35776
rect 25148 35630 25176 35770
rect 25136 35624 25188 35630
rect 25136 35566 25188 35572
rect 24860 35488 24912 35494
rect 24860 35430 24912 35436
rect 24872 35290 24900 35430
rect 24860 35284 24912 35290
rect 24860 35226 24912 35232
rect 25240 35222 25268 36230
rect 25228 35216 25280 35222
rect 25228 35158 25280 35164
rect 25332 34950 25360 36722
rect 25412 36304 25464 36310
rect 25412 36246 25464 36252
rect 25424 36106 25452 36246
rect 25412 36100 25464 36106
rect 25412 36042 25464 36048
rect 25516 35290 25544 37130
rect 25700 36378 25728 39200
rect 25872 37256 25924 37262
rect 25872 37198 25924 37204
rect 25884 36854 25912 37198
rect 25964 37188 26016 37194
rect 25964 37130 26016 37136
rect 25872 36848 25924 36854
rect 25872 36790 25924 36796
rect 25976 36718 26004 37130
rect 26516 37120 26568 37126
rect 26516 37062 26568 37068
rect 25964 36712 26016 36718
rect 25964 36654 26016 36660
rect 25964 36576 26016 36582
rect 25964 36518 26016 36524
rect 25688 36372 25740 36378
rect 25688 36314 25740 36320
rect 25504 35284 25556 35290
rect 25504 35226 25556 35232
rect 25320 34944 25372 34950
rect 25320 34886 25372 34892
rect 25688 34944 25740 34950
rect 25688 34886 25740 34892
rect 24768 34536 24820 34542
rect 24768 34478 24820 34484
rect 23940 3732 23992 3738
rect 23940 3674 23992 3680
rect 24676 3732 24728 3738
rect 24676 3674 24728 3680
rect 23952 3398 23980 3674
rect 24216 3460 24268 3466
rect 24216 3402 24268 3408
rect 23940 3392 23992 3398
rect 23940 3334 23992 3340
rect 24228 3194 24256 3402
rect 24688 3194 24716 3674
rect 24216 3188 24268 3194
rect 24216 3130 24268 3136
rect 24676 3188 24728 3194
rect 24676 3130 24728 3136
rect 24780 2650 24808 34478
rect 24952 3936 25004 3942
rect 24952 3878 25004 3884
rect 24964 3602 24992 3878
rect 24952 3596 25004 3602
rect 24952 3538 25004 3544
rect 24860 3392 24912 3398
rect 24860 3334 24912 3340
rect 24768 2644 24820 2650
rect 24768 2586 24820 2592
rect 23848 2508 23900 2514
rect 23848 2450 23900 2456
rect 24872 2378 24900 3334
rect 24964 3194 24992 3538
rect 24952 3188 25004 3194
rect 24952 3130 25004 3136
rect 25700 2650 25728 34886
rect 25976 33590 26004 36518
rect 26332 36304 26384 36310
rect 26332 36246 26384 36252
rect 26344 36106 26372 36246
rect 26332 36100 26384 36106
rect 26332 36042 26384 36048
rect 25964 33584 26016 33590
rect 25964 33526 26016 33532
rect 26528 32978 26556 37062
rect 26620 36174 26648 39200
rect 27344 37256 27396 37262
rect 27344 37198 27396 37204
rect 27252 37188 27304 37194
rect 27172 37148 27252 37176
rect 27172 36650 27200 37148
rect 27252 37130 27304 37136
rect 27356 36854 27384 37198
rect 27252 36848 27304 36854
rect 27252 36790 27304 36796
rect 27344 36848 27396 36854
rect 27344 36790 27396 36796
rect 27264 36650 27292 36790
rect 27160 36644 27212 36650
rect 27160 36586 27212 36592
rect 27252 36644 27304 36650
rect 27252 36586 27304 36592
rect 27356 36582 27384 36790
rect 26700 36576 26752 36582
rect 26700 36518 26752 36524
rect 27344 36576 27396 36582
rect 27344 36518 27396 36524
rect 26608 36168 26660 36174
rect 26608 36110 26660 36116
rect 26620 35834 26648 36110
rect 26608 35828 26660 35834
rect 26608 35770 26660 35776
rect 26516 32972 26568 32978
rect 26516 32914 26568 32920
rect 26712 26234 26740 36518
rect 27540 36394 27568 39200
rect 28170 37496 28226 37505
rect 28170 37431 28226 37440
rect 27988 37324 28040 37330
rect 27988 37266 28040 37272
rect 28000 36650 28028 37266
rect 28184 37126 28212 37431
rect 28172 37120 28224 37126
rect 28172 37062 28224 37068
rect 28460 36922 28488 39200
rect 29092 37664 29144 37670
rect 29092 37606 29144 37612
rect 29104 37398 29132 37606
rect 29092 37392 29144 37398
rect 28998 37360 29054 37369
rect 29092 37334 29144 37340
rect 28998 37295 29054 37304
rect 28724 37256 28776 37262
rect 28724 37198 28776 37204
rect 28908 37256 28960 37262
rect 29012 37210 29040 37295
rect 28960 37204 29040 37210
rect 28908 37198 29040 37204
rect 28632 37120 28684 37126
rect 28632 37062 28684 37068
rect 28356 36916 28408 36922
rect 28356 36858 28408 36864
rect 28448 36916 28500 36922
rect 28448 36858 28500 36864
rect 27988 36644 28040 36650
rect 27988 36586 28040 36592
rect 27540 36378 27660 36394
rect 27540 36372 27672 36378
rect 27540 36366 27620 36372
rect 27620 36314 27672 36320
rect 27896 36168 27948 36174
rect 27896 36110 27948 36116
rect 26792 36032 26844 36038
rect 26792 35974 26844 35980
rect 26804 35766 26832 35974
rect 26792 35760 26844 35766
rect 26792 35702 26844 35708
rect 27908 35562 27936 36110
rect 27896 35556 27948 35562
rect 27896 35498 27948 35504
rect 26620 26206 26740 26234
rect 26620 12434 26648 26206
rect 26528 12406 26648 12434
rect 26240 4616 26292 4622
rect 26240 4558 26292 4564
rect 26252 4010 26280 4558
rect 26332 4208 26384 4214
rect 26332 4150 26384 4156
rect 26240 4004 26292 4010
rect 26240 3946 26292 3952
rect 25964 3936 26016 3942
rect 25964 3878 26016 3884
rect 25872 3528 25924 3534
rect 25872 3470 25924 3476
rect 25884 3058 25912 3470
rect 25872 3052 25924 3058
rect 25872 2994 25924 3000
rect 25688 2644 25740 2650
rect 25688 2586 25740 2592
rect 25976 2378 26004 3878
rect 26252 3602 26280 3946
rect 26240 3596 26292 3602
rect 26240 3538 26292 3544
rect 26252 2514 26280 3538
rect 26344 3058 26372 4150
rect 26424 3392 26476 3398
rect 26424 3334 26476 3340
rect 26332 3052 26384 3058
rect 26332 2994 26384 3000
rect 26332 2848 26384 2854
rect 26332 2790 26384 2796
rect 26240 2508 26292 2514
rect 26240 2450 26292 2456
rect 26344 2446 26372 2790
rect 26332 2440 26384 2446
rect 26332 2382 26384 2388
rect 26436 2378 26464 3334
rect 26528 2650 26556 12406
rect 28368 5370 28396 36858
rect 28644 36786 28672 37062
rect 28632 36780 28684 36786
rect 28632 36722 28684 36728
rect 28540 36712 28592 36718
rect 28540 36654 28592 36660
rect 28552 35834 28580 36654
rect 28632 36644 28684 36650
rect 28632 36586 28684 36592
rect 28644 36038 28672 36586
rect 28632 36032 28684 36038
rect 28632 35974 28684 35980
rect 28644 35834 28672 35974
rect 28540 35828 28592 35834
rect 28540 35770 28592 35776
rect 28632 35828 28684 35834
rect 28632 35770 28684 35776
rect 28736 35290 28764 37198
rect 28920 37182 29040 37198
rect 29380 37194 29408 39200
rect 29644 37392 29696 37398
rect 29644 37334 29696 37340
rect 29368 37188 29420 37194
rect 29368 37130 29420 37136
rect 28816 36780 28868 36786
rect 28816 36722 28868 36728
rect 29092 36780 29144 36786
rect 29092 36722 29144 36728
rect 28724 35284 28776 35290
rect 28724 35226 28776 35232
rect 28356 5364 28408 5370
rect 28356 5306 28408 5312
rect 27620 4480 27672 4486
rect 27620 4422 27672 4428
rect 27344 4140 27396 4146
rect 27344 4082 27396 4088
rect 27160 3936 27212 3942
rect 27160 3878 27212 3884
rect 27172 3602 27200 3878
rect 27160 3596 27212 3602
rect 27160 3538 27212 3544
rect 27356 3194 27384 4082
rect 27528 3664 27580 3670
rect 27528 3606 27580 3612
rect 27344 3188 27396 3194
rect 27344 3130 27396 3136
rect 27540 3126 27568 3606
rect 27528 3120 27580 3126
rect 27528 3062 27580 3068
rect 27632 2990 27660 4422
rect 27896 3936 27948 3942
rect 27896 3878 27948 3884
rect 27988 3936 28040 3942
rect 27988 3878 28040 3884
rect 27908 3602 27936 3878
rect 28000 3670 28028 3878
rect 27988 3664 28040 3670
rect 27988 3606 28040 3612
rect 28078 3632 28134 3641
rect 27896 3596 27948 3602
rect 28078 3567 28080 3576
rect 27896 3538 27948 3544
rect 28132 3567 28134 3576
rect 28080 3538 28132 3544
rect 27988 3392 28040 3398
rect 27988 3334 28040 3340
rect 28000 3194 28028 3334
rect 27988 3188 28040 3194
rect 27988 3130 28040 3136
rect 28368 3126 28396 5306
rect 28828 4146 28856 36722
rect 28908 36644 28960 36650
rect 28908 36586 28960 36592
rect 28920 35766 28948 36586
rect 28908 35760 28960 35766
rect 28908 35702 28960 35708
rect 29104 34746 29132 36722
rect 29380 36378 29408 37130
rect 29656 36650 29684 37334
rect 30012 37324 30064 37330
rect 30012 37266 30064 37272
rect 29828 37188 29880 37194
rect 29828 37130 29880 37136
rect 29840 36922 29868 37130
rect 29828 36916 29880 36922
rect 29828 36858 29880 36864
rect 29644 36644 29696 36650
rect 29644 36586 29696 36592
rect 29368 36372 29420 36378
rect 29368 36314 29420 36320
rect 29276 36032 29328 36038
rect 29276 35974 29328 35980
rect 29288 35834 29316 35974
rect 29276 35828 29328 35834
rect 29276 35770 29328 35776
rect 30024 35737 30052 37266
rect 30300 36904 30328 39200
rect 31024 37664 31076 37670
rect 31024 37606 31076 37612
rect 31036 37466 31064 37606
rect 31024 37460 31076 37466
rect 31024 37402 31076 37408
rect 30748 37188 30800 37194
rect 30800 37148 30880 37176
rect 30748 37130 30800 37136
rect 30380 36916 30432 36922
rect 30300 36876 30380 36904
rect 30380 36858 30432 36864
rect 30564 36916 30616 36922
rect 30564 36858 30616 36864
rect 30576 36825 30604 36858
rect 30562 36816 30618 36825
rect 30562 36751 30618 36760
rect 30656 36780 30708 36786
rect 30656 36722 30708 36728
rect 30668 36378 30696 36722
rect 30656 36372 30708 36378
rect 30656 36314 30708 36320
rect 30010 35728 30066 35737
rect 30010 35663 30066 35672
rect 30668 35018 30696 36314
rect 30852 36174 30880 37148
rect 31220 37126 31248 39200
rect 31300 37256 31352 37262
rect 31300 37198 31352 37204
rect 31116 37120 31168 37126
rect 31116 37062 31168 37068
rect 31208 37120 31260 37126
rect 31208 37062 31260 37068
rect 31128 36786 31156 37062
rect 31116 36780 31168 36786
rect 31116 36722 31168 36728
rect 30840 36168 30892 36174
rect 30840 36110 30892 36116
rect 30852 35494 30880 36110
rect 31312 35562 31340 37198
rect 31760 37188 31812 37194
rect 31760 37130 31812 37136
rect 31484 37120 31536 37126
rect 31484 37062 31536 37068
rect 31496 36786 31524 37062
rect 31484 36780 31536 36786
rect 31484 36722 31536 36728
rect 31300 35556 31352 35562
rect 31300 35498 31352 35504
rect 30840 35488 30892 35494
rect 30840 35430 30892 35436
rect 30656 35012 30708 35018
rect 30656 34954 30708 34960
rect 29092 34740 29144 34746
rect 29092 34682 29144 34688
rect 30288 4616 30340 4622
rect 30340 4564 30420 4570
rect 30288 4558 30420 4564
rect 30300 4542 30420 4558
rect 30196 4480 30248 4486
rect 30196 4422 30248 4428
rect 28816 4140 28868 4146
rect 28816 4082 28868 4088
rect 28448 4072 28500 4078
rect 28448 4014 28500 4020
rect 28460 3210 28488 4014
rect 28724 3664 28776 3670
rect 28724 3606 28776 3612
rect 28460 3182 28672 3210
rect 28644 3126 28672 3182
rect 28356 3120 28408 3126
rect 28356 3062 28408 3068
rect 28632 3120 28684 3126
rect 28632 3062 28684 3068
rect 27620 2984 27672 2990
rect 27620 2926 27672 2932
rect 27896 2848 27948 2854
rect 27896 2790 27948 2796
rect 26516 2644 26568 2650
rect 26516 2586 26568 2592
rect 27908 2378 27936 2790
rect 24860 2372 24912 2378
rect 24860 2314 24912 2320
rect 25964 2372 26016 2378
rect 25964 2314 26016 2320
rect 26424 2372 26476 2378
rect 26424 2314 26476 2320
rect 27896 2372 27948 2378
rect 27896 2314 27948 2320
rect 23296 2100 23348 2106
rect 23296 2042 23348 2048
rect 24872 1986 24900 2314
rect 24596 1958 24900 1986
rect 24596 800 24624 1958
rect 25976 800 26004 2314
rect 27344 2304 27396 2310
rect 27344 2246 27396 2252
rect 27356 800 27384 2246
rect 28736 800 28764 3606
rect 28828 3194 28856 4082
rect 29828 4072 29880 4078
rect 29828 4014 29880 4020
rect 28816 3188 28868 3194
rect 28816 3130 28868 3136
rect 29840 3126 29868 4014
rect 30208 3602 30236 4422
rect 30288 3936 30340 3942
rect 30288 3878 30340 3884
rect 30196 3596 30248 3602
rect 30196 3538 30248 3544
rect 28908 3120 28960 3126
rect 28908 3062 28960 3068
rect 29828 3120 29880 3126
rect 29828 3062 29880 3068
rect 30104 3120 30156 3126
rect 30104 3062 30156 3068
rect 28920 2650 28948 3062
rect 28908 2644 28960 2650
rect 28908 2586 28960 2592
rect 30116 800 30144 3062
rect 30208 2774 30236 3538
rect 30300 3126 30328 3878
rect 30392 3602 30420 4542
rect 30380 3596 30432 3602
rect 30380 3538 30432 3544
rect 30748 3392 30800 3398
rect 30748 3334 30800 3340
rect 30288 3120 30340 3126
rect 30288 3062 30340 3068
rect 30208 2746 30328 2774
rect 30300 2446 30328 2746
rect 30288 2440 30340 2446
rect 30288 2382 30340 2388
rect 30760 2378 30788 3334
rect 30852 3194 30880 35430
rect 30840 3188 30892 3194
rect 30840 3130 30892 3136
rect 31496 3126 31524 36722
rect 31772 33969 31800 37130
rect 32140 36174 32168 39200
rect 32956 37188 33008 37194
rect 32956 37130 33008 37136
rect 32496 37120 32548 37126
rect 32496 37062 32548 37068
rect 32312 36372 32364 36378
rect 32312 36314 32364 36320
rect 32128 36168 32180 36174
rect 32128 36110 32180 36116
rect 32324 36038 32352 36314
rect 32312 36032 32364 36038
rect 32312 35974 32364 35980
rect 31944 35828 31996 35834
rect 31944 35770 31996 35776
rect 31956 35562 31984 35770
rect 31944 35556 31996 35562
rect 31944 35498 31996 35504
rect 31758 33960 31814 33969
rect 31758 33895 31814 33904
rect 32508 32842 32536 37062
rect 32968 36768 32996 37130
rect 33060 36904 33088 39200
rect 33600 37868 33652 37874
rect 33600 37810 33652 37816
rect 33416 37664 33468 37670
rect 33416 37606 33468 37612
rect 33140 36916 33192 36922
rect 33060 36876 33140 36904
rect 33140 36858 33192 36864
rect 33428 36786 33456 37606
rect 33612 37330 33640 37810
rect 33600 37324 33652 37330
rect 33600 37266 33652 37272
rect 33600 37188 33652 37194
rect 33600 37130 33652 37136
rect 33048 36780 33100 36786
rect 32968 36740 33048 36768
rect 33048 36722 33100 36728
rect 33140 36780 33192 36786
rect 33140 36722 33192 36728
rect 33416 36780 33468 36786
rect 33416 36722 33468 36728
rect 32956 35692 33008 35698
rect 32956 35634 33008 35640
rect 32968 35494 32996 35634
rect 32956 35488 33008 35494
rect 33060 35476 33088 36722
rect 33152 36038 33180 36722
rect 33612 36650 33640 37130
rect 33980 36786 34008 39200
rect 34336 37256 34388 37262
rect 34336 37198 34388 37204
rect 33968 36780 34020 36786
rect 33968 36722 34020 36728
rect 34244 36780 34296 36786
rect 34244 36722 34296 36728
rect 33600 36644 33652 36650
rect 33600 36586 33652 36592
rect 33232 36576 33284 36582
rect 33232 36518 33284 36524
rect 33784 36576 33836 36582
rect 33784 36518 33836 36524
rect 33244 36038 33272 36518
rect 33692 36372 33744 36378
rect 33796 36360 33824 36518
rect 33980 36378 34008 36722
rect 33744 36332 33824 36360
rect 33968 36372 34020 36378
rect 33692 36314 33744 36320
rect 33968 36314 34020 36320
rect 34256 36310 34284 36722
rect 34244 36304 34296 36310
rect 34244 36246 34296 36252
rect 33140 36032 33192 36038
rect 33140 35974 33192 35980
rect 33232 36032 33284 36038
rect 33232 35974 33284 35980
rect 34256 35766 34284 36246
rect 34348 35766 34376 37198
rect 34428 37120 34480 37126
rect 34532 37108 34560 39222
rect 34808 39114 34836 39222
rect 34886 39200 34942 40000
rect 35806 39200 35862 40000
rect 36726 39200 36782 40000
rect 37646 39200 37702 40000
rect 38566 39200 38622 40000
rect 39396 39296 39448 39302
rect 39396 39238 39448 39244
rect 34900 39114 34928 39200
rect 34808 39086 34928 39114
rect 35532 38820 35584 38826
rect 35532 38762 35584 38768
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34704 37256 34756 37262
rect 34704 37198 34756 37204
rect 34480 37080 34560 37108
rect 34428 37062 34480 37068
rect 34612 36576 34664 36582
rect 34612 36518 34664 36524
rect 34426 36272 34482 36281
rect 34624 36242 34652 36518
rect 34426 36207 34428 36216
rect 34480 36207 34482 36216
rect 34612 36236 34664 36242
rect 34428 36178 34480 36184
rect 34612 36178 34664 36184
rect 34716 36174 34744 37198
rect 35544 37194 35572 38762
rect 35532 37188 35584 37194
rect 35716 37188 35768 37194
rect 35532 37130 35584 37136
rect 35636 37148 35716 37176
rect 34796 37120 34848 37126
rect 34796 37062 34848 37068
rect 34704 36168 34756 36174
rect 34704 36110 34756 36116
rect 34244 35760 34296 35766
rect 34244 35702 34296 35708
rect 34336 35760 34388 35766
rect 34336 35702 34388 35708
rect 34704 35556 34756 35562
rect 34704 35498 34756 35504
rect 33140 35488 33192 35494
rect 33060 35448 33140 35476
rect 32956 35430 33008 35436
rect 33140 35430 33192 35436
rect 32496 32836 32548 32842
rect 32496 32778 32548 32784
rect 31760 29640 31812 29646
rect 31760 29582 31812 29588
rect 31668 3936 31720 3942
rect 31668 3878 31720 3884
rect 31680 3126 31708 3878
rect 31484 3120 31536 3126
rect 31484 3062 31536 3068
rect 31668 3120 31720 3126
rect 31668 3062 31720 3068
rect 31680 2774 31708 3062
rect 31496 2746 31708 2774
rect 30748 2372 30800 2378
rect 30748 2314 30800 2320
rect 31496 800 31524 2746
rect 31772 2446 31800 29582
rect 32312 4480 32364 4486
rect 32312 4422 32364 4428
rect 32772 4480 32824 4486
rect 32772 4422 32824 4428
rect 32324 3398 32352 4422
rect 32784 4282 32812 4422
rect 32772 4276 32824 4282
rect 32772 4218 32824 4224
rect 32784 3534 32812 4218
rect 33152 3738 33180 35430
rect 34716 35193 34744 35498
rect 34702 35184 34758 35193
rect 34702 35119 34758 35128
rect 34808 6914 34836 37062
rect 35348 36576 35400 36582
rect 35348 36518 35400 36524
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 35360 35154 35388 36518
rect 35544 35222 35572 37130
rect 35636 36650 35664 37148
rect 35716 37130 35768 37136
rect 35714 37088 35770 37097
rect 35714 37023 35770 37032
rect 35728 36650 35756 37023
rect 35624 36644 35676 36650
rect 35624 36586 35676 36592
rect 35716 36644 35768 36650
rect 35716 36586 35768 36592
rect 35820 36122 35848 39200
rect 36084 37120 36136 37126
rect 36084 37062 36136 37068
rect 36544 37120 36596 37126
rect 36636 37120 36688 37126
rect 36544 37062 36596 37068
rect 36634 37088 36636 37097
rect 36688 37088 36690 37097
rect 35992 36780 36044 36786
rect 35992 36722 36044 36728
rect 35900 36168 35952 36174
rect 35820 36116 35900 36122
rect 35820 36110 35952 36116
rect 35820 36094 35940 36110
rect 35820 35562 35848 36094
rect 36004 36038 36032 36722
rect 35992 36032 36044 36038
rect 35992 35974 36044 35980
rect 35808 35556 35860 35562
rect 35808 35498 35860 35504
rect 35532 35216 35584 35222
rect 35532 35158 35584 35164
rect 35348 35148 35400 35154
rect 35348 35090 35400 35096
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34440 6886 34836 6914
rect 33692 4548 33744 4554
rect 33692 4490 33744 4496
rect 33704 4146 33732 4490
rect 33692 4140 33744 4146
rect 33692 4082 33744 4088
rect 33784 4140 33836 4146
rect 33784 4082 33836 4088
rect 34152 4140 34204 4146
rect 34152 4082 34204 4088
rect 33324 3936 33376 3942
rect 33324 3878 33376 3884
rect 33140 3732 33192 3738
rect 33140 3674 33192 3680
rect 32772 3528 32824 3534
rect 32772 3470 32824 3476
rect 32312 3392 32364 3398
rect 32312 3334 32364 3340
rect 32324 2514 32352 3334
rect 32784 3058 32812 3470
rect 32864 3460 32916 3466
rect 32864 3402 32916 3408
rect 32772 3052 32824 3058
rect 32772 2994 32824 3000
rect 32312 2508 32364 2514
rect 32312 2450 32364 2456
rect 31760 2440 31812 2446
rect 31760 2382 31812 2388
rect 32876 800 32904 3402
rect 33336 2378 33364 3878
rect 33704 2990 33732 4082
rect 33796 3194 33824 4082
rect 33876 3936 33928 3942
rect 33876 3878 33928 3884
rect 33784 3188 33836 3194
rect 33784 3130 33836 3136
rect 33692 2984 33744 2990
rect 33692 2926 33744 2932
rect 33324 2372 33376 2378
rect 33324 2314 33376 2320
rect 33888 2310 33916 3878
rect 34164 3194 34192 4082
rect 34244 3936 34296 3942
rect 34244 3878 34296 3884
rect 34152 3188 34204 3194
rect 34152 3130 34204 3136
rect 34164 2650 34192 3130
rect 34152 2644 34204 2650
rect 34152 2586 34204 2592
rect 33876 2304 33928 2310
rect 33876 2246 33928 2252
rect 34256 800 34284 3878
rect 34440 3194 34468 6886
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34796 5092 34848 5098
rect 34796 5034 34848 5040
rect 34704 3392 34756 3398
rect 34704 3334 34756 3340
rect 34428 3188 34480 3194
rect 34428 3130 34480 3136
rect 34716 2378 34744 3334
rect 34808 2990 34836 5034
rect 35624 5024 35676 5030
rect 35624 4966 35676 4972
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 35636 4214 35664 4966
rect 35900 4480 35952 4486
rect 35900 4422 35952 4428
rect 35624 4208 35676 4214
rect 35624 4150 35676 4156
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34796 2984 34848 2990
rect 34796 2926 34848 2932
rect 34808 2514 34836 2926
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34796 2508 34848 2514
rect 34796 2450 34848 2456
rect 34704 2372 34756 2378
rect 34704 2314 34756 2320
rect 35636 800 35664 4150
rect 35716 3596 35768 3602
rect 35716 3538 35768 3544
rect 35728 3448 35756 3538
rect 35808 3460 35860 3466
rect 35728 3420 35808 3448
rect 35808 3402 35860 3408
rect 35912 2378 35940 4422
rect 36004 4146 36032 35974
rect 36096 5370 36124 37062
rect 36452 36916 36504 36922
rect 36452 36858 36504 36864
rect 36464 36825 36492 36858
rect 36450 36816 36506 36825
rect 36450 36751 36506 36760
rect 36556 36378 36584 37062
rect 36634 37023 36690 37032
rect 36544 36372 36596 36378
rect 36544 36314 36596 36320
rect 36360 36304 36412 36310
rect 36412 36264 36492 36292
rect 36360 36246 36412 36252
rect 36464 36258 36492 36264
rect 36464 36242 36584 36258
rect 36464 36236 36596 36242
rect 36464 36230 36544 36236
rect 36544 36178 36596 36184
rect 36544 36032 36596 36038
rect 36544 35974 36596 35980
rect 36556 35086 36584 35974
rect 36648 35222 36676 37023
rect 36740 36922 36768 39200
rect 36818 37360 36874 37369
rect 36818 37295 36874 37304
rect 37556 37324 37608 37330
rect 36832 36922 36860 37295
rect 37556 37266 37608 37272
rect 36728 36916 36780 36922
rect 36728 36858 36780 36864
rect 36820 36916 36872 36922
rect 36820 36858 36872 36864
rect 37280 36848 37332 36854
rect 37094 36816 37150 36825
rect 36912 36780 36964 36786
rect 37280 36790 37332 36796
rect 37094 36751 37096 36760
rect 36912 36722 36964 36728
rect 37148 36751 37150 36760
rect 37096 36722 37148 36728
rect 36636 35216 36688 35222
rect 36636 35158 36688 35164
rect 36924 35086 36952 36722
rect 37188 36576 37240 36582
rect 37188 36518 37240 36524
rect 36544 35080 36596 35086
rect 36544 35022 36596 35028
rect 36912 35080 36964 35086
rect 36912 35022 36964 35028
rect 37200 34513 37228 36518
rect 37292 36310 37320 36790
rect 37568 36582 37596 37266
rect 37556 36576 37608 36582
rect 37556 36518 37608 36524
rect 37280 36304 37332 36310
rect 37280 36246 37332 36252
rect 37280 36168 37332 36174
rect 37280 36110 37332 36116
rect 37292 35494 37320 36110
rect 37568 35850 37596 36518
rect 37660 36174 37688 39200
rect 38200 37120 38252 37126
rect 38200 37062 38252 37068
rect 38476 37120 38528 37126
rect 38580 37108 38608 39200
rect 39408 37262 39436 39238
rect 39486 39200 39542 40000
rect 40406 39200 40462 40000
rect 41326 39200 41382 40000
rect 42246 39200 42302 40000
rect 42616 39364 42668 39370
rect 42616 39306 42668 39312
rect 39396 37256 39448 37262
rect 39396 37198 39448 37204
rect 38660 37120 38712 37126
rect 38580 37080 38660 37108
rect 38476 37062 38528 37068
rect 38660 37062 38712 37068
rect 38108 36848 38160 36854
rect 38108 36790 38160 36796
rect 37648 36168 37700 36174
rect 37648 36110 37700 36116
rect 37476 35834 37596 35850
rect 37660 35834 37688 36110
rect 37464 35828 37596 35834
rect 37516 35822 37596 35828
rect 37648 35828 37700 35834
rect 37464 35770 37516 35776
rect 37648 35770 37700 35776
rect 38120 35494 38148 36790
rect 37280 35488 37332 35494
rect 37280 35430 37332 35436
rect 38108 35488 38160 35494
rect 38108 35430 38160 35436
rect 37186 34504 37242 34513
rect 37186 34439 37242 34448
rect 37292 26234 37320 35430
rect 37292 26206 37688 26234
rect 36084 5364 36136 5370
rect 36084 5306 36136 5312
rect 35992 4140 36044 4146
rect 35992 4082 36044 4088
rect 35992 3596 36044 3602
rect 35992 3538 36044 3544
rect 36004 2990 36032 3538
rect 36096 3466 36124 5306
rect 36912 4684 36964 4690
rect 36912 4626 36964 4632
rect 36924 4554 36952 4626
rect 36912 4548 36964 4554
rect 36912 4490 36964 4496
rect 36084 3460 36136 3466
rect 36084 3402 36136 3408
rect 36924 2990 36952 4490
rect 37280 4480 37332 4486
rect 37280 4422 37332 4428
rect 37292 4214 37320 4422
rect 37280 4208 37332 4214
rect 37280 4150 37332 4156
rect 37292 4026 37320 4150
rect 37660 4146 37688 26206
rect 38212 5370 38240 37062
rect 38488 36530 38516 37062
rect 38844 36780 38896 36786
rect 38844 36722 38896 36728
rect 38566 36544 38622 36553
rect 38488 36502 38566 36530
rect 38566 36479 38622 36488
rect 38580 35850 38608 36479
rect 38580 35834 38700 35850
rect 38580 35828 38712 35834
rect 38580 35822 38660 35828
rect 38660 35770 38712 35776
rect 38856 34134 38884 36722
rect 39304 36576 39356 36582
rect 39304 36518 39356 36524
rect 39316 36378 39344 36518
rect 39304 36372 39356 36378
rect 39304 36314 39356 36320
rect 39408 35834 39436 37198
rect 39500 36378 39528 39200
rect 40040 37732 40092 37738
rect 40040 37674 40092 37680
rect 40052 37262 40080 37674
rect 40040 37256 40092 37262
rect 40040 37198 40092 37204
rect 40132 37256 40184 37262
rect 40132 37198 40184 37204
rect 40314 37224 40370 37233
rect 39946 36408 40002 36417
rect 39488 36372 39540 36378
rect 39946 36343 40002 36352
rect 39488 36314 39540 36320
rect 39500 36174 39528 36314
rect 39960 36242 39988 36343
rect 39948 36236 40000 36242
rect 39948 36178 40000 36184
rect 39488 36168 39540 36174
rect 39488 36110 39540 36116
rect 40052 36038 40080 37198
rect 40144 36854 40172 37198
rect 40314 37159 40370 37168
rect 40132 36848 40184 36854
rect 40132 36790 40184 36796
rect 40224 36780 40276 36786
rect 40224 36722 40276 36728
rect 40040 36032 40092 36038
rect 40040 35974 40092 35980
rect 39396 35828 39448 35834
rect 39396 35770 39448 35776
rect 40236 35494 40264 36722
rect 40328 36650 40356 37159
rect 40420 37126 40448 39200
rect 40868 37324 40920 37330
rect 40868 37266 40920 37272
rect 40408 37120 40460 37126
rect 40408 37062 40460 37068
rect 40592 37120 40644 37126
rect 40592 37062 40644 37068
rect 40316 36644 40368 36650
rect 40316 36586 40368 36592
rect 40224 35488 40276 35494
rect 40224 35430 40276 35436
rect 38844 34128 38896 34134
rect 38844 34070 38896 34076
rect 38200 5364 38252 5370
rect 38200 5306 38252 5312
rect 38016 4616 38068 4622
rect 38016 4558 38068 4564
rect 38028 4146 38056 4558
rect 37464 4140 37516 4146
rect 37464 4082 37516 4088
rect 37648 4140 37700 4146
rect 37648 4082 37700 4088
rect 38016 4140 38068 4146
rect 38016 4082 38068 4088
rect 37016 3998 37320 4026
rect 35992 2984 36044 2990
rect 35992 2926 36044 2932
rect 36912 2984 36964 2990
rect 36912 2926 36964 2932
rect 35900 2372 35952 2378
rect 35900 2314 35952 2320
rect 37016 800 37044 3998
rect 37096 3528 37148 3534
rect 37096 3470 37148 3476
rect 37108 3398 37136 3470
rect 37096 3392 37148 3398
rect 37096 3334 37148 3340
rect 37108 2650 37136 3334
rect 37476 3194 37504 4082
rect 37740 3936 37792 3942
rect 37740 3878 37792 3884
rect 37464 3188 37516 3194
rect 37464 3130 37516 3136
rect 37096 2644 37148 2650
rect 37096 2586 37148 2592
rect 37752 2378 37780 3878
rect 38212 3618 38240 5306
rect 38568 5092 38620 5098
rect 38568 5034 38620 5040
rect 38580 4486 38608 5034
rect 39856 4616 39908 4622
rect 39856 4558 39908 4564
rect 38568 4480 38620 4486
rect 38568 4422 38620 4428
rect 38580 4010 38608 4422
rect 39868 4146 39896 4558
rect 39856 4140 39908 4146
rect 39856 4082 39908 4088
rect 40040 4140 40092 4146
rect 40040 4082 40092 4088
rect 38568 4004 38620 4010
rect 38568 3946 38620 3952
rect 38580 3670 38608 3946
rect 38752 3936 38804 3942
rect 38752 3878 38804 3884
rect 39212 3936 39264 3942
rect 39212 3878 39264 3884
rect 39948 3936 40000 3942
rect 39948 3878 40000 3884
rect 38120 3590 38240 3618
rect 38568 3664 38620 3670
rect 38568 3606 38620 3612
rect 38120 3194 38148 3590
rect 38200 3460 38252 3466
rect 38200 3402 38252 3408
rect 38108 3188 38160 3194
rect 38108 3130 38160 3136
rect 38212 3126 38240 3402
rect 38384 3392 38436 3398
rect 38384 3334 38436 3340
rect 38200 3120 38252 3126
rect 38200 3062 38252 3068
rect 37740 2372 37792 2378
rect 37740 2314 37792 2320
rect 38396 800 38424 3334
rect 38580 3058 38608 3606
rect 38568 3052 38620 3058
rect 38568 2994 38620 3000
rect 38476 2508 38528 2514
rect 38580 2496 38608 2994
rect 38528 2468 38608 2496
rect 38476 2450 38528 2456
rect 38764 2378 38792 3878
rect 39224 3126 39252 3878
rect 39764 3392 39816 3398
rect 39764 3334 39816 3340
rect 39212 3120 39264 3126
rect 39212 3062 39264 3068
rect 39212 2984 39264 2990
rect 39212 2926 39264 2932
rect 39224 2650 39252 2926
rect 39212 2644 39264 2650
rect 39212 2586 39264 2592
rect 38752 2372 38804 2378
rect 38752 2314 38804 2320
rect 39776 800 39804 3334
rect 39960 3126 39988 3878
rect 39948 3120 40000 3126
rect 39948 3062 40000 3068
rect 40052 2650 40080 4082
rect 40236 3738 40264 35430
rect 40604 4826 40632 37062
rect 40880 34950 40908 37266
rect 41340 37210 41368 39200
rect 41156 37182 41368 37210
rect 40960 36780 41012 36786
rect 40960 36722 41012 36728
rect 40972 35494 41000 36722
rect 41050 36680 41106 36689
rect 41050 36615 41052 36624
rect 41104 36615 41106 36624
rect 41052 36586 41104 36592
rect 41156 36174 41184 37182
rect 41236 37120 41288 37126
rect 41236 37062 41288 37068
rect 41512 37120 41564 37126
rect 41512 37062 41564 37068
rect 41144 36168 41196 36174
rect 41050 36136 41106 36145
rect 41248 36145 41276 37062
rect 41328 36644 41380 36650
rect 41328 36586 41380 36592
rect 41144 36110 41196 36116
rect 41234 36136 41290 36145
rect 41050 36071 41052 36080
rect 41104 36071 41106 36080
rect 41234 36071 41290 36080
rect 41052 36042 41104 36048
rect 41236 35828 41288 35834
rect 41236 35770 41288 35776
rect 41248 35698 41276 35770
rect 41236 35692 41288 35698
rect 41236 35634 41288 35640
rect 41144 35624 41196 35630
rect 41142 35592 41144 35601
rect 41196 35592 41198 35601
rect 41142 35527 41198 35536
rect 40960 35488 41012 35494
rect 40960 35430 41012 35436
rect 40868 34944 40920 34950
rect 40868 34886 40920 34892
rect 40592 4820 40644 4826
rect 40592 4762 40644 4768
rect 40224 3732 40276 3738
rect 40224 3674 40276 3680
rect 40040 2644 40092 2650
rect 40040 2586 40092 2592
rect 40604 2378 40632 4762
rect 40972 3738 41000 35430
rect 41340 33561 41368 36586
rect 41524 36242 41552 37062
rect 41604 36916 41656 36922
rect 41604 36858 41656 36864
rect 41512 36236 41564 36242
rect 41512 36178 41564 36184
rect 41420 35624 41472 35630
rect 41418 35592 41420 35601
rect 41472 35592 41474 35601
rect 41418 35527 41474 35536
rect 41326 33552 41382 33561
rect 41326 33487 41382 33496
rect 41616 12434 41644 36858
rect 41972 36576 42024 36582
rect 41972 36518 42024 36524
rect 42064 36576 42116 36582
rect 42064 36518 42116 36524
rect 41694 36136 41750 36145
rect 41694 36071 41750 36080
rect 41708 35222 41736 36071
rect 41696 35216 41748 35222
rect 41696 35158 41748 35164
rect 41984 34105 42012 36518
rect 42076 36038 42104 36518
rect 42260 36378 42288 39200
rect 42248 36372 42300 36378
rect 42248 36314 42300 36320
rect 42628 36174 42656 39306
rect 43166 39200 43222 40000
rect 44086 39200 44142 40000
rect 45006 39200 45062 40000
rect 45926 39200 45982 40000
rect 46296 39228 46348 39234
rect 42708 37256 42760 37262
rect 42708 37198 42760 37204
rect 42800 37256 42852 37262
rect 42800 37198 42852 37204
rect 42720 36922 42748 37198
rect 42708 36916 42760 36922
rect 42708 36858 42760 36864
rect 42812 36786 42840 37198
rect 43074 36816 43130 36825
rect 42800 36780 42852 36786
rect 43074 36751 43130 36760
rect 42800 36722 42852 36728
rect 42616 36168 42668 36174
rect 42616 36110 42668 36116
rect 42064 36032 42116 36038
rect 42064 35974 42116 35980
rect 42628 35834 42656 36110
rect 42524 35828 42576 35834
rect 42524 35770 42576 35776
rect 42616 35828 42668 35834
rect 42616 35770 42668 35776
rect 42536 35562 42564 35770
rect 42524 35556 42576 35562
rect 42524 35498 42576 35504
rect 42812 35494 42840 36722
rect 43088 36718 43116 36751
rect 43076 36712 43128 36718
rect 43076 36654 43128 36660
rect 42892 36372 42944 36378
rect 42892 36314 42944 36320
rect 42904 36281 42932 36314
rect 42890 36272 42946 36281
rect 42890 36207 42946 36216
rect 42800 35488 42852 35494
rect 42800 35430 42852 35436
rect 42812 34950 42840 35430
rect 43088 35222 43116 36654
rect 43180 35834 43208 39200
rect 43996 39024 44048 39030
rect 43996 38966 44048 38972
rect 43812 37188 43864 37194
rect 43812 37130 43864 37136
rect 43444 37120 43496 37126
rect 43444 37062 43496 37068
rect 43720 37120 43772 37126
rect 43720 37062 43772 37068
rect 43168 35828 43220 35834
rect 43168 35770 43220 35776
rect 43076 35216 43128 35222
rect 43076 35158 43128 35164
rect 43352 35080 43404 35086
rect 43350 35048 43352 35057
rect 43404 35048 43406 35057
rect 43350 34983 43406 34992
rect 42800 34944 42852 34950
rect 42800 34886 42852 34892
rect 41970 34096 42026 34105
rect 41970 34031 42026 34040
rect 41524 12406 41644 12434
rect 41328 4480 41380 4486
rect 41380 4428 41460 4434
rect 41328 4422 41460 4428
rect 41340 4406 41460 4422
rect 41144 3936 41196 3942
rect 41144 3878 41196 3884
rect 40960 3732 41012 3738
rect 40960 3674 41012 3680
rect 41156 3466 41184 3878
rect 41144 3460 41196 3466
rect 41144 3402 41196 3408
rect 40684 2848 40736 2854
rect 40684 2790 40736 2796
rect 40696 2446 40724 2790
rect 40684 2440 40736 2446
rect 40684 2382 40736 2388
rect 40592 2372 40644 2378
rect 40592 2314 40644 2320
rect 41156 800 41184 3402
rect 41432 2990 41460 4406
rect 41524 3126 41552 12406
rect 42708 5024 42760 5030
rect 42708 4966 42760 4972
rect 42720 4826 42748 4966
rect 42708 4820 42760 4826
rect 42708 4762 42760 4768
rect 42432 4616 42484 4622
rect 42432 4558 42484 4564
rect 42156 4140 42208 4146
rect 42156 4082 42208 4088
rect 41604 4004 41656 4010
rect 41604 3946 41656 3952
rect 41616 3602 41644 3946
rect 41880 3936 41932 3942
rect 41880 3878 41932 3884
rect 41892 3602 41920 3878
rect 41604 3596 41656 3602
rect 41604 3538 41656 3544
rect 41880 3596 41932 3602
rect 41880 3538 41932 3544
rect 41512 3120 41564 3126
rect 41512 3062 41564 3068
rect 41420 2984 41472 2990
rect 41420 2926 41472 2932
rect 41432 2514 41460 2926
rect 41524 2650 41552 3062
rect 41694 2952 41750 2961
rect 41694 2887 41696 2896
rect 41748 2887 41750 2896
rect 41696 2858 41748 2864
rect 42168 2854 42196 4082
rect 42444 4010 42472 4558
rect 42432 4004 42484 4010
rect 42432 3946 42484 3952
rect 42524 3392 42576 3398
rect 42524 3334 42576 3340
rect 42536 3058 42564 3334
rect 42524 3052 42576 3058
rect 42524 2994 42576 3000
rect 42616 3052 42668 3058
rect 42616 2994 42668 3000
rect 42536 2854 42564 2994
rect 42628 2961 42656 2994
rect 42614 2952 42670 2961
rect 42614 2887 42670 2896
rect 42156 2848 42208 2854
rect 42156 2790 42208 2796
rect 42524 2848 42576 2854
rect 42524 2790 42576 2796
rect 42720 2774 42748 4762
rect 43456 4758 43484 37062
rect 43732 36417 43760 37062
rect 43718 36408 43774 36417
rect 43718 36343 43774 36352
rect 43824 36281 43852 37130
rect 44008 36786 44036 38966
rect 44100 36922 44128 39200
rect 44088 36916 44140 36922
rect 44088 36858 44140 36864
rect 44180 36916 44232 36922
rect 44180 36858 44232 36864
rect 43996 36780 44048 36786
rect 43996 36722 44048 36728
rect 43810 36272 43866 36281
rect 43810 36207 43866 36216
rect 43824 34678 43852 36207
rect 44008 35222 44036 36722
rect 44192 36689 44220 36858
rect 45020 36786 45048 39200
rect 45376 37800 45428 37806
rect 45376 37742 45428 37748
rect 45388 37466 45416 37742
rect 45376 37460 45428 37466
rect 45376 37402 45428 37408
rect 45376 37256 45428 37262
rect 45296 37204 45376 37210
rect 45296 37198 45428 37204
rect 45296 37182 45416 37198
rect 45652 37188 45704 37194
rect 44640 36780 44692 36786
rect 44640 36722 44692 36728
rect 45008 36780 45060 36786
rect 45008 36722 45060 36728
rect 44178 36680 44234 36689
rect 44178 36615 44234 36624
rect 44178 36408 44234 36417
rect 44178 36343 44234 36352
rect 44088 36168 44140 36174
rect 44088 36110 44140 36116
rect 44100 35834 44128 36110
rect 44192 36038 44220 36343
rect 44652 36106 44680 36722
rect 44824 36644 44876 36650
rect 44824 36586 44876 36592
rect 44364 36100 44416 36106
rect 44364 36042 44416 36048
rect 44640 36100 44692 36106
rect 44640 36042 44692 36048
rect 44180 36032 44232 36038
rect 44180 35974 44232 35980
rect 44088 35828 44140 35834
rect 44088 35770 44140 35776
rect 44376 35494 44404 36042
rect 44364 35488 44416 35494
rect 44364 35430 44416 35436
rect 43996 35216 44048 35222
rect 43996 35158 44048 35164
rect 43812 34672 43864 34678
rect 43812 34614 43864 34620
rect 43444 4752 43496 4758
rect 43444 4694 43496 4700
rect 42984 4480 43036 4486
rect 42984 4422 43036 4428
rect 42892 3936 42944 3942
rect 42892 3878 42944 3884
rect 42628 2746 42748 2774
rect 41512 2644 41564 2650
rect 41512 2586 41564 2592
rect 42628 2514 42656 2746
rect 41420 2508 41472 2514
rect 41420 2450 41472 2456
rect 42616 2508 42668 2514
rect 42616 2450 42668 2456
rect 42904 2378 42932 3878
rect 42996 3534 43024 4422
rect 43352 3664 43404 3670
rect 43352 3606 43404 3612
rect 42984 3528 43036 3534
rect 42984 3470 43036 3476
rect 43364 3126 43392 3606
rect 43456 3602 43484 4694
rect 44376 4146 44404 35430
rect 44456 35148 44508 35154
rect 44456 35090 44508 35096
rect 44468 35018 44496 35090
rect 44548 35080 44600 35086
rect 44546 35048 44548 35057
rect 44600 35048 44602 35057
rect 44456 35012 44508 35018
rect 44546 34983 44602 34992
rect 44456 34954 44508 34960
rect 44836 32774 44864 36586
rect 45020 35834 45048 36722
rect 45296 36038 45324 37182
rect 45652 37130 45704 37136
rect 45836 37188 45888 37194
rect 45836 37130 45888 37136
rect 45284 36032 45336 36038
rect 45282 36000 45284 36009
rect 45336 36000 45338 36009
rect 45282 35935 45338 35944
rect 45008 35828 45060 35834
rect 45008 35770 45060 35776
rect 45664 34950 45692 37130
rect 45848 36650 45876 37130
rect 45940 36650 45968 39200
rect 46846 39200 46902 40000
rect 47766 39200 47822 40000
rect 48686 39200 48742 40000
rect 49606 39200 49662 40000
rect 50526 39200 50582 40000
rect 51446 39200 51502 40000
rect 52366 39200 52422 40000
rect 53286 39200 53342 40000
rect 54206 39200 54262 40000
rect 55126 39200 55182 40000
rect 56046 39200 56102 40000
rect 56612 39222 56916 39250
rect 46296 39170 46348 39176
rect 46204 37324 46256 37330
rect 46204 37266 46256 37272
rect 45836 36644 45888 36650
rect 45836 36586 45888 36592
rect 45928 36644 45980 36650
rect 45928 36586 45980 36592
rect 45652 34944 45704 34950
rect 45652 34886 45704 34892
rect 46020 34944 46072 34950
rect 46020 34886 46072 34892
rect 44824 32768 44876 32774
rect 44824 32710 44876 32716
rect 45928 4480 45980 4486
rect 45928 4422 45980 4428
rect 43812 4140 43864 4146
rect 43812 4082 43864 4088
rect 43904 4140 43956 4146
rect 43904 4082 43956 4088
rect 44364 4140 44416 4146
rect 44364 4082 44416 4088
rect 43824 3738 43852 4082
rect 43916 3942 43944 4082
rect 43904 3936 43956 3942
rect 43904 3878 43956 3884
rect 45100 3936 45152 3942
rect 45100 3878 45152 3884
rect 45468 3936 45520 3942
rect 45468 3878 45520 3884
rect 43812 3732 43864 3738
rect 43812 3674 43864 3680
rect 43444 3596 43496 3602
rect 43444 3538 43496 3544
rect 43352 3120 43404 3126
rect 43352 3062 43404 3068
rect 42892 2372 42944 2378
rect 42892 2314 42944 2320
rect 42524 2304 42576 2310
rect 42524 2246 42576 2252
rect 42536 800 42564 2246
rect 43916 800 43944 3878
rect 45112 3534 45140 3878
rect 45100 3528 45152 3534
rect 45100 3470 45152 3476
rect 44180 3460 44232 3466
rect 44180 3402 44232 3408
rect 44192 2650 44220 3402
rect 45284 3392 45336 3398
rect 45284 3334 45336 3340
rect 44180 2644 44232 2650
rect 44180 2586 44232 2592
rect 45296 2378 45324 3334
rect 45480 3058 45508 3878
rect 45940 3534 45968 4422
rect 45928 3528 45980 3534
rect 45928 3470 45980 3476
rect 46032 3126 46060 34886
rect 46216 33658 46244 37266
rect 46308 36786 46336 39170
rect 46296 36780 46348 36786
rect 46296 36722 46348 36728
rect 46308 35834 46336 36722
rect 46756 36576 46808 36582
rect 46756 36518 46808 36524
rect 46296 35828 46348 35834
rect 46296 35770 46348 35776
rect 46768 35766 46796 36518
rect 46860 36174 46888 39200
rect 46940 38956 46992 38962
rect 46940 38898 46992 38904
rect 46952 37262 46980 38898
rect 46940 37256 46992 37262
rect 46940 37198 46992 37204
rect 46848 36168 46900 36174
rect 46848 36110 46900 36116
rect 46952 35834 46980 37198
rect 47780 37126 47808 39200
rect 48044 38276 48096 38282
rect 48044 38218 48096 38224
rect 47860 37460 47912 37466
rect 47860 37402 47912 37408
rect 47872 37330 47900 37402
rect 47860 37324 47912 37330
rect 47860 37266 47912 37272
rect 47768 37120 47820 37126
rect 47768 37062 47820 37068
rect 47216 36780 47268 36786
rect 47216 36722 47268 36728
rect 47308 36780 47360 36786
rect 47308 36722 47360 36728
rect 47032 36576 47084 36582
rect 47032 36518 47084 36524
rect 47124 36576 47176 36582
rect 47124 36518 47176 36524
rect 46940 35828 46992 35834
rect 46940 35770 46992 35776
rect 46756 35760 46808 35766
rect 46756 35702 46808 35708
rect 47044 34746 47072 36518
rect 47136 35494 47164 36518
rect 47228 36242 47256 36722
rect 47320 36310 47348 36722
rect 47872 36718 47900 37266
rect 48056 36718 48084 38218
rect 48136 37324 48188 37330
rect 48136 37266 48188 37272
rect 47860 36712 47912 36718
rect 47860 36654 47912 36660
rect 48044 36712 48096 36718
rect 48044 36654 48096 36660
rect 47872 36582 47900 36654
rect 48056 36582 48084 36654
rect 47860 36576 47912 36582
rect 47860 36518 47912 36524
rect 48044 36576 48096 36582
rect 48044 36518 48096 36524
rect 47308 36304 47360 36310
rect 47308 36246 47360 36252
rect 47216 36236 47268 36242
rect 47216 36178 47268 36184
rect 48148 35494 48176 37266
rect 48504 37256 48556 37262
rect 48504 37198 48556 37204
rect 48228 36576 48280 36582
rect 48228 36518 48280 36524
rect 47124 35488 47176 35494
rect 47124 35430 47176 35436
rect 48136 35488 48188 35494
rect 48136 35430 48188 35436
rect 47136 35018 47164 35430
rect 47124 35012 47176 35018
rect 47124 34954 47176 34960
rect 47032 34740 47084 34746
rect 47032 34682 47084 34688
rect 46204 33652 46256 33658
rect 46204 33594 46256 33600
rect 48148 32910 48176 35430
rect 48240 35018 48268 36518
rect 48516 36174 48544 37198
rect 48596 36780 48648 36786
rect 48596 36722 48648 36728
rect 48608 36310 48636 36722
rect 48596 36304 48648 36310
rect 48596 36246 48648 36252
rect 48504 36168 48556 36174
rect 48504 36110 48556 36116
rect 48412 36100 48464 36106
rect 48412 36042 48464 36048
rect 48424 35630 48452 36042
rect 48412 35624 48464 35630
rect 48412 35566 48464 35572
rect 48608 35494 48636 36246
rect 48700 36174 48728 39200
rect 49620 37126 49648 39200
rect 49792 38888 49844 38894
rect 49792 38830 49844 38836
rect 49804 37262 49832 38830
rect 49792 37256 49844 37262
rect 49792 37198 49844 37204
rect 50540 37210 50568 39200
rect 51172 38004 51224 38010
rect 51172 37946 51224 37952
rect 51184 37262 51212 37946
rect 51172 37256 51224 37262
rect 48964 37120 49016 37126
rect 48964 37062 49016 37068
rect 49608 37120 49660 37126
rect 49608 37062 49660 37068
rect 48688 36168 48740 36174
rect 48688 36110 48740 36116
rect 48700 35834 48728 36110
rect 48688 35828 48740 35834
rect 48688 35770 48740 35776
rect 48596 35488 48648 35494
rect 48596 35430 48648 35436
rect 48228 35012 48280 35018
rect 48228 34954 48280 34960
rect 48136 32904 48188 32910
rect 48136 32846 48188 32852
rect 47124 5024 47176 5030
rect 47124 4966 47176 4972
rect 48136 5024 48188 5030
rect 48136 4966 48188 4972
rect 48320 5024 48372 5030
rect 48320 4966 48372 4972
rect 47136 4554 47164 4966
rect 48148 4690 48176 4966
rect 47584 4684 47636 4690
rect 47584 4626 47636 4632
rect 48136 4684 48188 4690
rect 48136 4626 48188 4632
rect 47216 4616 47268 4622
rect 47216 4558 47268 4564
rect 47124 4548 47176 4554
rect 47124 4490 47176 4496
rect 47032 4480 47084 4486
rect 47032 4422 47084 4428
rect 47044 4146 47072 4422
rect 47032 4140 47084 4146
rect 47032 4082 47084 4088
rect 46112 4072 46164 4078
rect 46112 4014 46164 4020
rect 46124 3738 46152 4014
rect 46204 3936 46256 3942
rect 46204 3878 46256 3884
rect 46296 3936 46348 3942
rect 46940 3936 46992 3942
rect 46296 3878 46348 3884
rect 46768 3896 46940 3924
rect 46112 3732 46164 3738
rect 46112 3674 46164 3680
rect 46020 3120 46072 3126
rect 46020 3062 46072 3068
rect 45468 3052 45520 3058
rect 45468 2994 45520 3000
rect 45480 2774 45508 2994
rect 45388 2746 45508 2774
rect 45284 2372 45336 2378
rect 45284 2314 45336 2320
rect 45388 2258 45416 2746
rect 46216 2378 46244 3878
rect 46308 2514 46336 3878
rect 46768 3534 46796 3896
rect 46940 3878 46992 3884
rect 46756 3528 46808 3534
rect 46756 3470 46808 3476
rect 46848 3528 46900 3534
rect 46848 3470 46900 3476
rect 46860 3194 46888 3470
rect 46848 3188 46900 3194
rect 46848 3130 46900 3136
rect 46664 2848 46716 2854
rect 46664 2790 46716 2796
rect 46296 2508 46348 2514
rect 46296 2450 46348 2456
rect 46204 2372 46256 2378
rect 46204 2314 46256 2320
rect 45296 2230 45416 2258
rect 45296 800 45324 2230
rect 46676 800 46704 2790
rect 47228 2650 47256 4558
rect 47596 4554 47624 4626
rect 48332 4554 48360 4966
rect 48608 4826 48636 35430
rect 48976 4826 49004 37062
rect 49516 36644 49568 36650
rect 49516 36586 49568 36592
rect 49148 36576 49200 36582
rect 49148 36518 49200 36524
rect 49160 32434 49188 36518
rect 49148 32428 49200 32434
rect 49148 32370 49200 32376
rect 49056 5024 49108 5030
rect 49056 4966 49108 4972
rect 48596 4820 48648 4826
rect 48596 4762 48648 4768
rect 48964 4820 49016 4826
rect 48964 4762 49016 4768
rect 47584 4548 47636 4554
rect 47584 4490 47636 4496
rect 48320 4548 48372 4554
rect 48320 4490 48372 4496
rect 47596 4078 47624 4490
rect 47584 4072 47636 4078
rect 47584 4014 47636 4020
rect 47676 3392 47728 3398
rect 47676 3334 47728 3340
rect 47768 3392 47820 3398
rect 47768 3334 47820 3340
rect 47216 2644 47268 2650
rect 47216 2586 47268 2592
rect 47688 2378 47716 3334
rect 47780 2514 47808 3334
rect 48332 2774 48360 4490
rect 48976 4146 49004 4762
rect 49068 4282 49096 4966
rect 49528 4826 49556 36586
rect 49700 36100 49752 36106
rect 49700 36042 49752 36048
rect 49712 35494 49740 36042
rect 49700 35488 49752 35494
rect 49700 35430 49752 35436
rect 49608 5024 49660 5030
rect 49608 4966 49660 4972
rect 49516 4820 49568 4826
rect 49516 4762 49568 4768
rect 49620 4758 49648 4966
rect 49608 4752 49660 4758
rect 49608 4694 49660 4700
rect 49056 4276 49108 4282
rect 49056 4218 49108 4224
rect 48964 4140 49016 4146
rect 48964 4082 49016 4088
rect 49068 3534 49096 4218
rect 49516 4208 49568 4214
rect 49516 4150 49568 4156
rect 49424 4140 49476 4146
rect 49424 4082 49476 4088
rect 49332 4004 49384 4010
rect 49332 3946 49384 3952
rect 49344 3534 49372 3946
rect 49056 3528 49108 3534
rect 49056 3470 49108 3476
rect 49332 3528 49384 3534
rect 49332 3470 49384 3476
rect 49344 3058 49372 3470
rect 49332 3052 49384 3058
rect 49332 2994 49384 3000
rect 48056 2746 48360 2774
rect 47768 2508 47820 2514
rect 47768 2450 47820 2456
rect 47676 2372 47728 2378
rect 47676 2314 47728 2320
rect 48056 800 48084 2746
rect 49436 800 49464 4082
rect 49528 2650 49556 4150
rect 49712 4146 49740 35430
rect 49804 35018 49832 37198
rect 50540 37182 50660 37210
rect 51172 37198 51224 37204
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 50252 36780 50304 36786
rect 50252 36722 50304 36728
rect 50264 36106 50292 36722
rect 50632 36174 50660 37182
rect 50896 36780 50948 36786
rect 50896 36722 50948 36728
rect 50620 36168 50672 36174
rect 50620 36110 50672 36116
rect 50252 36100 50304 36106
rect 50252 36042 50304 36048
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 50632 35834 50660 36110
rect 50712 36032 50764 36038
rect 50710 36000 50712 36009
rect 50764 36000 50766 36009
rect 50710 35935 50766 35944
rect 50620 35828 50672 35834
rect 50620 35770 50672 35776
rect 50908 35601 50936 36722
rect 50894 35592 50950 35601
rect 50894 35527 50950 35536
rect 51184 35018 51212 37198
rect 51460 37126 51488 39200
rect 51724 37460 51776 37466
rect 51724 37402 51776 37408
rect 51736 37330 51764 37402
rect 51724 37324 51776 37330
rect 51724 37266 51776 37272
rect 51448 37120 51500 37126
rect 51448 37062 51500 37068
rect 51540 37120 51592 37126
rect 51540 37062 51592 37068
rect 51262 36680 51318 36689
rect 51262 36615 51318 36624
rect 51276 36310 51304 36615
rect 51448 36576 51500 36582
rect 51448 36518 51500 36524
rect 51264 36304 51316 36310
rect 51264 36246 51316 36252
rect 51460 35193 51488 36518
rect 51552 36038 51580 37062
rect 51632 36780 51684 36786
rect 51632 36722 51684 36728
rect 51540 36032 51592 36038
rect 51540 35974 51592 35980
rect 51446 35184 51502 35193
rect 51446 35119 51502 35128
rect 49792 35012 49844 35018
rect 49792 34954 49844 34960
rect 51172 35012 51224 35018
rect 51172 34954 51224 34960
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 51552 33046 51580 35974
rect 51644 35494 51672 36722
rect 51736 35834 51764 37266
rect 52380 37210 52408 39200
rect 53196 38412 53248 38418
rect 53196 38354 53248 38360
rect 52288 37182 52408 37210
rect 53010 37224 53066 37233
rect 52092 36780 52144 36786
rect 52092 36722 52144 36728
rect 51816 36712 51868 36718
rect 51816 36654 51868 36660
rect 51828 36582 51856 36654
rect 51816 36576 51868 36582
rect 51816 36518 51868 36524
rect 51724 35828 51776 35834
rect 51724 35770 51776 35776
rect 52104 35562 52132 36722
rect 52288 36174 52316 37182
rect 53010 37159 53066 37168
rect 52368 37120 52420 37126
rect 52368 37062 52420 37068
rect 52276 36168 52328 36174
rect 52276 36110 52328 36116
rect 52288 35834 52316 36110
rect 52276 35828 52328 35834
rect 52276 35770 52328 35776
rect 52092 35556 52144 35562
rect 52092 35498 52144 35504
rect 51632 35488 51684 35494
rect 51632 35430 51684 35436
rect 51540 33040 51592 33046
rect 51540 32982 51592 32988
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 52380 5370 52408 37062
rect 53024 36922 53052 37159
rect 53208 37126 53236 38354
rect 53196 37120 53248 37126
rect 53196 37062 53248 37068
rect 53012 36916 53064 36922
rect 53012 36858 53064 36864
rect 53104 36916 53156 36922
rect 53104 36858 53156 36864
rect 53012 36780 53064 36786
rect 53012 36722 53064 36728
rect 53024 36650 53052 36722
rect 53012 36644 53064 36650
rect 53012 36586 53064 36592
rect 53024 36417 53052 36586
rect 53010 36408 53066 36417
rect 53010 36343 53066 36352
rect 53012 36304 53064 36310
rect 53012 36246 53064 36252
rect 52736 36100 52788 36106
rect 52736 36042 52788 36048
rect 52920 36100 52972 36106
rect 52920 36042 52972 36048
rect 52748 35494 52776 36042
rect 52736 35488 52788 35494
rect 52736 35430 52788 35436
rect 52932 32502 52960 36042
rect 53024 36038 53052 36246
rect 53116 36174 53144 36858
rect 53104 36168 53156 36174
rect 53104 36110 53156 36116
rect 53012 36032 53064 36038
rect 53012 35974 53064 35980
rect 53104 35488 53156 35494
rect 53104 35430 53156 35436
rect 52920 32496 52972 32502
rect 52920 32438 52972 32444
rect 52092 5364 52144 5370
rect 52092 5306 52144 5312
rect 52368 5364 52420 5370
rect 52368 5306 52420 5312
rect 51448 4616 51500 4622
rect 51448 4558 51500 4564
rect 50620 4480 50672 4486
rect 50620 4422 50672 4428
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 49700 4140 49752 4146
rect 49700 4082 49752 4088
rect 50632 3942 50660 4422
rect 51460 4214 51488 4558
rect 51632 4480 51684 4486
rect 51632 4422 51684 4428
rect 51448 4208 51500 4214
rect 51448 4150 51500 4156
rect 51356 4140 51408 4146
rect 51356 4082 51408 4088
rect 50620 3936 50672 3942
rect 50620 3878 50672 3884
rect 50896 3936 50948 3942
rect 50896 3878 50948 3884
rect 50632 3398 50660 3878
rect 50620 3392 50672 3398
rect 50620 3334 50672 3340
rect 50804 3392 50856 3398
rect 50804 3334 50856 3340
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 50632 3058 50660 3334
rect 50620 3052 50672 3058
rect 50620 2994 50672 3000
rect 50068 2848 50120 2854
rect 50068 2790 50120 2796
rect 49516 2644 49568 2650
rect 49516 2586 49568 2592
rect 50080 2378 50108 2790
rect 50632 2650 50660 2994
rect 50620 2644 50672 2650
rect 50620 2586 50672 2592
rect 50068 2372 50120 2378
rect 50068 2314 50120 2320
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50816 800 50844 3334
rect 50908 3126 50936 3878
rect 51368 3738 51396 4082
rect 51460 4010 51488 4150
rect 51448 4004 51500 4010
rect 51448 3946 51500 3952
rect 51540 3936 51592 3942
rect 51540 3878 51592 3884
rect 51356 3732 51408 3738
rect 51356 3674 51408 3680
rect 50896 3120 50948 3126
rect 50896 3062 50948 3068
rect 51552 2514 51580 3878
rect 51644 3126 51672 4422
rect 52104 3602 52132 5306
rect 53012 5024 53064 5030
rect 53012 4966 53064 4972
rect 52460 4480 52512 4486
rect 52460 4422 52512 4428
rect 52472 4214 52500 4422
rect 52460 4208 52512 4214
rect 52460 4150 52512 4156
rect 52184 4140 52236 4146
rect 52184 4082 52236 4088
rect 52092 3596 52144 3602
rect 52092 3538 52144 3544
rect 51908 3460 51960 3466
rect 51908 3402 51960 3408
rect 51632 3120 51684 3126
rect 51632 3062 51684 3068
rect 51920 2514 51948 3402
rect 52196 2922 52224 4082
rect 52472 4026 52500 4150
rect 52380 3998 52500 4026
rect 52276 3936 52328 3942
rect 52276 3878 52328 3884
rect 52184 2916 52236 2922
rect 52184 2858 52236 2864
rect 51540 2508 51592 2514
rect 51540 2450 51592 2456
rect 51908 2508 51960 2514
rect 51908 2450 51960 2456
rect 52288 2378 52316 3878
rect 52276 2372 52328 2378
rect 52276 2314 52328 2320
rect 52380 2258 52408 3998
rect 53024 3534 53052 4966
rect 53116 4146 53144 35430
rect 53208 35018 53236 37062
rect 53300 36360 53328 39200
rect 53564 37664 53616 37670
rect 53564 37606 53616 37612
rect 53576 37194 53604 37606
rect 53564 37188 53616 37194
rect 53564 37130 53616 37136
rect 53656 37120 53708 37126
rect 53656 37062 53708 37068
rect 53380 36372 53432 36378
rect 53300 36332 53380 36360
rect 53380 36314 53432 36320
rect 53196 35012 53248 35018
rect 53196 34954 53248 34960
rect 53668 6914 53696 37062
rect 53932 36780 53984 36786
rect 53932 36722 53984 36728
rect 53748 36576 53800 36582
rect 53748 36518 53800 36524
rect 53760 35873 53788 36518
rect 53746 35864 53802 35873
rect 53746 35799 53802 35808
rect 53944 35494 53972 36722
rect 54220 36718 54248 39200
rect 54944 38752 54996 38758
rect 54944 38694 54996 38700
rect 54300 37936 54352 37942
rect 54300 37878 54352 37884
rect 54208 36712 54260 36718
rect 54208 36654 54260 36660
rect 54312 36378 54340 37878
rect 54956 37262 54984 38694
rect 54944 37256 54996 37262
rect 54944 37198 54996 37204
rect 54760 36712 54812 36718
rect 54760 36654 54812 36660
rect 54392 36576 54444 36582
rect 54392 36518 54444 36524
rect 54300 36372 54352 36378
rect 54300 36314 54352 36320
rect 54312 36174 54340 36314
rect 54300 36168 54352 36174
rect 54300 36110 54352 36116
rect 53932 35488 53984 35494
rect 53932 35430 53984 35436
rect 53668 6886 53880 6914
rect 53852 4826 53880 6886
rect 53840 4820 53892 4826
rect 53840 4762 53892 4768
rect 53104 4140 53156 4146
rect 53104 4082 53156 4088
rect 53288 3732 53340 3738
rect 53288 3674 53340 3680
rect 52460 3528 52512 3534
rect 52460 3470 52512 3476
rect 53012 3528 53064 3534
rect 53012 3470 53064 3476
rect 52472 2990 52500 3470
rect 53300 3126 53328 3674
rect 53564 3460 53616 3466
rect 53564 3402 53616 3408
rect 53288 3120 53340 3126
rect 53288 3062 53340 3068
rect 52460 2984 52512 2990
rect 52460 2926 52512 2932
rect 53300 2582 53328 3062
rect 53288 2576 53340 2582
rect 53288 2518 53340 2524
rect 52196 2230 52408 2258
rect 52196 800 52224 2230
rect 53576 800 53604 3402
rect 53852 3126 53880 4762
rect 53944 3670 53972 35430
rect 54404 35018 54432 36518
rect 54772 36378 54800 36654
rect 54760 36372 54812 36378
rect 54760 36314 54812 36320
rect 54956 35834 54984 37198
rect 55140 37126 55168 39200
rect 55220 37664 55272 37670
rect 55220 37606 55272 37612
rect 55232 37466 55260 37606
rect 55220 37460 55272 37466
rect 55220 37402 55272 37408
rect 55678 37224 55734 37233
rect 55588 37188 55640 37194
rect 55678 37159 55680 37168
rect 55588 37130 55640 37136
rect 55732 37159 55734 37168
rect 55680 37130 55732 37136
rect 55128 37120 55180 37126
rect 55128 37062 55180 37068
rect 55600 36786 55628 37130
rect 56060 36786 56088 39200
rect 56140 37664 56192 37670
rect 56140 37606 56192 37612
rect 56152 37262 56180 37606
rect 56140 37256 56192 37262
rect 56140 37198 56192 37204
rect 56508 37120 56560 37126
rect 56612 37108 56640 39222
rect 56888 39114 56916 39222
rect 56966 39200 57022 40000
rect 57886 39200 57942 40000
rect 58806 39200 58862 40000
rect 59726 39200 59782 40000
rect 60646 39200 60702 40000
rect 61566 39200 61622 40000
rect 61672 39222 62068 39250
rect 56980 39114 57008 39200
rect 56888 39086 57008 39114
rect 57520 37460 57572 37466
rect 57520 37402 57572 37408
rect 56692 37256 56744 37262
rect 56692 37198 56744 37204
rect 56560 37080 56640 37108
rect 56508 37062 56560 37068
rect 55588 36780 55640 36786
rect 55588 36722 55640 36728
rect 56048 36780 56100 36786
rect 56048 36722 56100 36728
rect 55128 36576 55180 36582
rect 55128 36518 55180 36524
rect 55140 36310 55168 36518
rect 56060 36378 56088 36722
rect 56600 36712 56652 36718
rect 56600 36654 56652 36660
rect 56048 36372 56100 36378
rect 56048 36314 56100 36320
rect 56140 36372 56192 36378
rect 56140 36314 56192 36320
rect 55128 36304 55180 36310
rect 55128 36246 55180 36252
rect 56152 36009 56180 36314
rect 56612 36038 56640 36654
rect 56704 36582 56732 37198
rect 57532 37126 57560 37402
rect 56784 37120 56836 37126
rect 56784 37062 56836 37068
rect 57152 37120 57204 37126
rect 57152 37062 57204 37068
rect 57520 37120 57572 37126
rect 57520 37062 57572 37068
rect 56692 36576 56744 36582
rect 56692 36518 56744 36524
rect 56600 36032 56652 36038
rect 56138 36000 56194 36009
rect 56600 35974 56652 35980
rect 56138 35935 56194 35944
rect 54944 35828 54996 35834
rect 54944 35770 54996 35776
rect 56612 35494 56640 35974
rect 56600 35488 56652 35494
rect 56600 35430 56652 35436
rect 54392 35012 54444 35018
rect 54392 34954 54444 34960
rect 55864 33108 55916 33114
rect 55864 33050 55916 33056
rect 54300 4480 54352 4486
rect 54300 4422 54352 4428
rect 54312 4282 54340 4422
rect 54300 4276 54352 4282
rect 54300 4218 54352 4224
rect 54024 3936 54076 3942
rect 54024 3878 54076 3884
rect 53932 3664 53984 3670
rect 53932 3606 53984 3612
rect 54036 3194 54064 3878
rect 54208 3596 54260 3602
rect 54208 3538 54260 3544
rect 54024 3188 54076 3194
rect 54024 3130 54076 3136
rect 53840 3120 53892 3126
rect 53840 3062 53892 3068
rect 54220 2990 54248 3538
rect 54312 3398 54340 4218
rect 55876 4146 55904 33050
rect 56324 4480 56376 4486
rect 56324 4422 56376 4428
rect 56416 4480 56468 4486
rect 56416 4422 56468 4428
rect 56336 4214 56364 4422
rect 56324 4208 56376 4214
rect 56324 4150 56376 4156
rect 55864 4140 55916 4146
rect 55864 4082 55916 4088
rect 55220 3936 55272 3942
rect 55220 3878 55272 3884
rect 55128 3528 55180 3534
rect 55128 3470 55180 3476
rect 54300 3392 54352 3398
rect 54300 3334 54352 3340
rect 54576 3392 54628 3398
rect 54576 3334 54628 3340
rect 54208 2984 54260 2990
rect 54208 2926 54260 2932
rect 54220 2514 54248 2926
rect 54208 2508 54260 2514
rect 54208 2450 54260 2456
rect 54312 2446 54340 3334
rect 54588 3126 54616 3334
rect 54576 3120 54628 3126
rect 54576 3062 54628 3068
rect 54944 2576 54996 2582
rect 54944 2518 54996 2524
rect 54300 2440 54352 2446
rect 54300 2382 54352 2388
rect 54956 800 54984 2518
rect 55140 2514 55168 3470
rect 55232 3126 55260 3878
rect 55876 3602 55904 4082
rect 55864 3596 55916 3602
rect 55864 3538 55916 3544
rect 56048 3392 56100 3398
rect 56048 3334 56100 3340
rect 55220 3120 55272 3126
rect 55220 3062 55272 3068
rect 56060 2854 56088 3334
rect 55680 2848 55732 2854
rect 55680 2790 55732 2796
rect 56048 2848 56100 2854
rect 56048 2790 56100 2796
rect 55692 2514 55720 2790
rect 55128 2508 55180 2514
rect 55128 2450 55180 2456
rect 55680 2508 55732 2514
rect 55680 2450 55732 2456
rect 56060 2038 56088 2790
rect 56048 2032 56100 2038
rect 56048 1974 56100 1980
rect 56336 800 56364 4150
rect 56428 3398 56456 4422
rect 56612 4146 56640 35430
rect 56796 33114 56824 37062
rect 57164 36689 57192 37062
rect 57336 36780 57388 36786
rect 57336 36722 57388 36728
rect 57428 36780 57480 36786
rect 57428 36722 57480 36728
rect 57150 36680 57206 36689
rect 57150 36615 57206 36624
rect 57060 36576 57112 36582
rect 57060 36518 57112 36524
rect 57072 35154 57100 36518
rect 57152 36100 57204 36106
rect 57152 36042 57204 36048
rect 57060 35148 57112 35154
rect 57060 35090 57112 35096
rect 56784 33108 56836 33114
rect 56784 33050 56836 33056
rect 57164 32366 57192 36042
rect 57348 35494 57376 36722
rect 57440 35698 57468 36722
rect 57428 35692 57480 35698
rect 57428 35634 57480 35640
rect 57336 35488 57388 35494
rect 57336 35430 57388 35436
rect 57152 32360 57204 32366
rect 57152 32302 57204 32308
rect 56600 4140 56652 4146
rect 56600 4082 56652 4088
rect 57152 4072 57204 4078
rect 57152 4014 57204 4020
rect 56508 4004 56560 4010
rect 56508 3946 56560 3952
rect 56416 3392 56468 3398
rect 56416 3334 56468 3340
rect 56520 3058 56548 3946
rect 56600 3936 56652 3942
rect 56600 3878 56652 3884
rect 56508 3052 56560 3058
rect 56508 2994 56560 3000
rect 56612 2310 56640 3878
rect 57164 3534 57192 4014
rect 57152 3528 57204 3534
rect 57152 3470 57204 3476
rect 57348 3194 57376 35430
rect 57532 34474 57560 37062
rect 57900 36700 57928 39200
rect 58532 38208 58584 38214
rect 58532 38150 58584 38156
rect 58346 37496 58402 37505
rect 58164 37460 58216 37466
rect 58346 37431 58402 37440
rect 58164 37402 58216 37408
rect 57980 37120 58032 37126
rect 58032 37080 58112 37108
rect 57980 37062 58032 37068
rect 57900 36672 58020 36700
rect 57992 36174 58020 36672
rect 57980 36168 58032 36174
rect 57980 36110 58032 36116
rect 57992 35834 58020 36110
rect 58084 36106 58112 37080
rect 58072 36100 58124 36106
rect 58072 36042 58124 36048
rect 57980 35828 58032 35834
rect 57980 35770 58032 35776
rect 57520 34468 57572 34474
rect 57520 34410 57572 34416
rect 58176 28994 58204 37402
rect 58360 37398 58388 37431
rect 58348 37392 58400 37398
rect 58254 37360 58310 37369
rect 58348 37334 58400 37340
rect 58254 37295 58256 37304
rect 58308 37295 58310 37304
rect 58256 37266 58308 37272
rect 58268 36718 58296 37266
rect 58348 37256 58400 37262
rect 58346 37224 58348 37233
rect 58400 37224 58402 37233
rect 58346 37159 58402 37168
rect 58544 36718 58572 38150
rect 58716 38072 58768 38078
rect 58716 38014 58768 38020
rect 58622 37360 58678 37369
rect 58622 37295 58624 37304
rect 58676 37295 58678 37304
rect 58624 37266 58676 37272
rect 58728 37210 58756 38014
rect 58636 37182 58756 37210
rect 58636 37126 58664 37182
rect 58624 37120 58676 37126
rect 58624 37062 58676 37068
rect 58716 37120 58768 37126
rect 58716 37062 58768 37068
rect 58256 36712 58308 36718
rect 58256 36654 58308 36660
rect 58532 36712 58584 36718
rect 58532 36654 58584 36660
rect 58544 35154 58572 36654
rect 58636 35834 58664 37062
rect 58728 36378 58756 37062
rect 58820 36378 58848 39200
rect 59084 36576 59136 36582
rect 59084 36518 59136 36524
rect 58716 36372 58768 36378
rect 58716 36314 58768 36320
rect 58808 36372 58860 36378
rect 58808 36314 58860 36320
rect 58900 36100 58952 36106
rect 58900 36042 58952 36048
rect 58624 35828 58676 35834
rect 58624 35770 58676 35776
rect 58912 35494 58940 36042
rect 58900 35488 58952 35494
rect 58900 35430 58952 35436
rect 58532 35148 58584 35154
rect 58532 35090 58584 35096
rect 58176 28966 58388 28994
rect 58360 26234 58388 28966
rect 58360 26206 58756 26234
rect 58728 6914 58756 26206
rect 58636 6886 58756 6914
rect 58072 5024 58124 5030
rect 58072 4966 58124 4972
rect 57980 4820 58032 4826
rect 57980 4762 58032 4768
rect 57796 4548 57848 4554
rect 57796 4490 57848 4496
rect 57428 4140 57480 4146
rect 57428 4082 57480 4088
rect 57440 3738 57468 4082
rect 57428 3732 57480 3738
rect 57428 3674 57480 3680
rect 57704 3732 57756 3738
rect 57704 3674 57756 3680
rect 57716 3466 57744 3674
rect 57704 3460 57756 3466
rect 57704 3402 57756 3408
rect 57808 3398 57836 4490
rect 57992 3466 58020 4762
rect 57980 3460 58032 3466
rect 57980 3402 58032 3408
rect 57428 3392 57480 3398
rect 57428 3334 57480 3340
rect 57796 3392 57848 3398
rect 57796 3334 57848 3340
rect 57336 3188 57388 3194
rect 57336 3130 57388 3136
rect 56692 2848 56744 2854
rect 56692 2790 56744 2796
rect 56704 2378 56732 2790
rect 56692 2372 56744 2378
rect 56692 2314 56744 2320
rect 57440 2310 57468 3334
rect 58084 3126 58112 4966
rect 58636 4826 58664 6886
rect 58716 5024 58768 5030
rect 58716 4966 58768 4972
rect 58624 4820 58676 4826
rect 58624 4762 58676 4768
rect 58164 4616 58216 4622
rect 58164 4558 58216 4564
rect 57704 3120 57756 3126
rect 57704 3062 57756 3068
rect 58072 3120 58124 3126
rect 58072 3062 58124 3068
rect 56600 2304 56652 2310
rect 56600 2246 56652 2252
rect 57428 2304 57480 2310
rect 57428 2246 57480 2252
rect 57440 2106 57468 2246
rect 57428 2100 57480 2106
rect 57428 2042 57480 2048
rect 57716 800 57744 3062
rect 58176 2922 58204 4558
rect 58348 4480 58400 4486
rect 58348 4422 58400 4428
rect 58164 2916 58216 2922
rect 58164 2858 58216 2864
rect 58360 2378 58388 4422
rect 58624 3596 58676 3602
rect 58624 3538 58676 3544
rect 58636 2990 58664 3538
rect 58728 3398 58756 4966
rect 59096 4826 59124 36518
rect 59740 36242 59768 39200
rect 59912 38684 59964 38690
rect 59912 38626 59964 38632
rect 59818 37496 59874 37505
rect 59818 37431 59874 37440
rect 59832 37398 59860 37431
rect 59820 37392 59872 37398
rect 59820 37334 59872 37340
rect 59820 37188 59872 37194
rect 59820 37130 59872 37136
rect 59832 36378 59860 37130
rect 59820 36372 59872 36378
rect 59820 36314 59872 36320
rect 59728 36236 59780 36242
rect 59728 36178 59780 36184
rect 59924 36174 59952 38626
rect 60096 38616 60148 38622
rect 60096 38558 60148 38564
rect 60108 36786 60136 38558
rect 60660 36922 60688 39200
rect 61580 39114 61608 39200
rect 61672 39114 61700 39222
rect 61580 39086 61700 39114
rect 61292 38548 61344 38554
rect 61292 38490 61344 38496
rect 61108 37392 61160 37398
rect 61108 37334 61160 37340
rect 61016 37256 61068 37262
rect 60752 37216 61016 37244
rect 60752 37126 60780 37216
rect 61016 37198 61068 37204
rect 60740 37120 60792 37126
rect 60740 37062 60792 37068
rect 60648 36916 60700 36922
rect 60648 36858 60700 36864
rect 60096 36780 60148 36786
rect 60096 36722 60148 36728
rect 60740 36780 60792 36786
rect 60740 36722 60792 36728
rect 59912 36168 59964 36174
rect 59912 36110 59964 36116
rect 59268 36100 59320 36106
rect 59268 36042 59320 36048
rect 59280 34746 59308 36042
rect 59924 35154 59952 36110
rect 60108 35834 60136 36722
rect 60372 36168 60424 36174
rect 60372 36110 60424 36116
rect 60384 35834 60412 36110
rect 60096 35828 60148 35834
rect 60096 35770 60148 35776
rect 60372 35828 60424 35834
rect 60372 35770 60424 35776
rect 60752 35494 60780 36722
rect 61016 36576 61068 36582
rect 61016 36518 61068 36524
rect 60740 35488 60792 35494
rect 60740 35430 60792 35436
rect 59912 35148 59964 35154
rect 59912 35090 59964 35096
rect 60752 34950 60780 35430
rect 60740 34944 60792 34950
rect 60740 34886 60792 34892
rect 59268 34740 59320 34746
rect 59268 34682 59320 34688
rect 59084 4820 59136 4826
rect 59084 4762 59136 4768
rect 59096 3482 59124 4762
rect 60752 4146 60780 34886
rect 61028 34066 61056 36518
rect 61016 34060 61068 34066
rect 61016 34002 61068 34008
rect 60832 5092 60884 5098
rect 60832 5034 60884 5040
rect 60464 4140 60516 4146
rect 60464 4082 60516 4088
rect 60740 4140 60792 4146
rect 60740 4082 60792 4088
rect 59360 4004 59412 4010
rect 59360 3946 59412 3952
rect 59004 3454 59124 3482
rect 58716 3392 58768 3398
rect 58716 3334 58768 3340
rect 58728 3194 58756 3334
rect 58716 3188 58768 3194
rect 58716 3130 58768 3136
rect 58624 2984 58676 2990
rect 58624 2926 58676 2932
rect 58728 2514 58756 3130
rect 59004 3126 59032 3454
rect 59084 3392 59136 3398
rect 59084 3334 59136 3340
rect 58992 3120 59044 3126
rect 58992 3062 59044 3068
rect 58716 2508 58768 2514
rect 58716 2450 58768 2456
rect 58348 2372 58400 2378
rect 58348 2314 58400 2320
rect 59096 800 59124 3334
rect 59372 2378 59400 3946
rect 59636 3936 59688 3942
rect 59636 3878 59688 3884
rect 59648 3058 59676 3878
rect 60004 3392 60056 3398
rect 60004 3334 60056 3340
rect 60016 3126 60044 3334
rect 60004 3120 60056 3126
rect 60004 3062 60056 3068
rect 59636 3052 59688 3058
rect 59636 2994 59688 3000
rect 59648 2938 59676 2994
rect 59648 2910 59860 2938
rect 59360 2372 59412 2378
rect 59360 2314 59412 2320
rect 59832 2310 59860 2910
rect 59820 2304 59872 2310
rect 59820 2246 59872 2252
rect 59832 1630 59860 2246
rect 59820 1624 59872 1630
rect 59820 1566 59872 1572
rect 60476 800 60504 4082
rect 60844 2650 60872 5034
rect 61120 4826 61148 37334
rect 61304 37330 61332 38490
rect 61382 37360 61438 37369
rect 61292 37324 61344 37330
rect 61382 37295 61384 37304
rect 61292 37266 61344 37272
rect 61436 37295 61438 37304
rect 61384 37266 61436 37272
rect 61304 35834 61332 37266
rect 61396 36174 61424 37266
rect 61752 37256 61804 37262
rect 61752 37198 61804 37204
rect 61660 36780 61712 36786
rect 61660 36722 61712 36728
rect 61672 36378 61700 36722
rect 61660 36372 61712 36378
rect 61660 36314 61712 36320
rect 61384 36168 61436 36174
rect 61384 36110 61436 36116
rect 61672 36106 61700 36314
rect 61660 36100 61712 36106
rect 61660 36042 61712 36048
rect 61764 36009 61792 37198
rect 62040 36768 62068 39222
rect 62486 39200 62542 40000
rect 63406 39200 63462 40000
rect 64326 39200 64382 40000
rect 65246 39200 65302 40000
rect 66166 39200 66222 40000
rect 67086 39200 67142 40000
rect 68006 39200 68062 40000
rect 68652 39296 68704 39302
rect 68652 39238 68704 39244
rect 62396 37460 62448 37466
rect 62396 37402 62448 37408
rect 62408 37194 62436 37402
rect 62396 37188 62448 37194
rect 62396 37130 62448 37136
rect 62120 36780 62172 36786
rect 62040 36740 62120 36768
rect 62120 36722 62172 36728
rect 62028 36100 62080 36106
rect 62028 36042 62080 36048
rect 61750 36000 61806 36009
rect 61750 35935 61806 35944
rect 61292 35828 61344 35834
rect 61292 35770 61344 35776
rect 61764 34950 61792 35935
rect 62040 35494 62068 36042
rect 62028 35488 62080 35494
rect 62028 35430 62080 35436
rect 62040 34950 62068 35430
rect 62132 35154 62160 36722
rect 62408 36718 62436 37130
rect 62396 36712 62448 36718
rect 62396 36654 62448 36660
rect 62500 36378 62528 39200
rect 62856 38480 62908 38486
rect 62856 38422 62908 38428
rect 62672 37800 62724 37806
rect 62672 37742 62724 37748
rect 62580 37188 62632 37194
rect 62580 37130 62632 37136
rect 62488 36372 62540 36378
rect 62488 36314 62540 36320
rect 62592 36310 62620 37130
rect 62580 36304 62632 36310
rect 62580 36246 62632 36252
rect 62580 36168 62632 36174
rect 62580 36110 62632 36116
rect 62120 35148 62172 35154
rect 62120 35090 62172 35096
rect 62592 34950 62620 36110
rect 61200 34944 61252 34950
rect 61200 34886 61252 34892
rect 61752 34944 61804 34950
rect 61752 34886 61804 34892
rect 62028 34944 62080 34950
rect 62028 34886 62080 34892
rect 62580 34944 62632 34950
rect 62580 34886 62632 34892
rect 61212 29646 61240 34886
rect 62040 31634 62068 34886
rect 62684 31754 62712 37742
rect 62868 36174 62896 38422
rect 63420 36786 63448 39200
rect 63500 39092 63552 39098
rect 63500 39034 63552 39040
rect 63512 37262 63540 39034
rect 63500 37256 63552 37262
rect 63500 37198 63552 37204
rect 64144 37256 64196 37262
rect 64144 37198 64196 37204
rect 63592 37120 63644 37126
rect 63592 37062 63644 37068
rect 64052 37120 64104 37126
rect 64052 37062 64104 37068
rect 63408 36780 63460 36786
rect 63408 36722 63460 36728
rect 63316 36576 63368 36582
rect 63316 36518 63368 36524
rect 63328 36310 63356 36518
rect 63316 36304 63368 36310
rect 63316 36246 63368 36252
rect 62856 36168 62908 36174
rect 62856 36110 62908 36116
rect 62868 35154 62896 36110
rect 63420 35834 63448 36722
rect 63500 36576 63552 36582
rect 63500 36518 63552 36524
rect 63408 35828 63460 35834
rect 63408 35770 63460 35776
rect 62856 35148 62908 35154
rect 62856 35090 62908 35096
rect 62672 31748 62724 31754
rect 62672 31690 62724 31696
rect 62040 31606 62160 31634
rect 61200 29640 61252 29646
rect 61200 29582 61252 29588
rect 61844 5024 61896 5030
rect 61844 4966 61896 4972
rect 61108 4820 61160 4826
rect 61108 4762 61160 4768
rect 61120 3602 61148 4762
rect 61476 4480 61528 4486
rect 61476 4422 61528 4428
rect 61384 3936 61436 3942
rect 61384 3878 61436 3884
rect 61108 3596 61160 3602
rect 61108 3538 61160 3544
rect 61200 3392 61252 3398
rect 61200 3334 61252 3340
rect 60832 2644 60884 2650
rect 60832 2586 60884 2592
rect 61212 2378 61240 3334
rect 61396 3126 61424 3878
rect 61488 3466 61516 4422
rect 61476 3460 61528 3466
rect 61476 3402 61528 3408
rect 61384 3120 61436 3126
rect 61384 3062 61436 3068
rect 61488 2990 61516 3402
rect 61856 3058 61884 4966
rect 62028 3528 62080 3534
rect 62028 3470 62080 3476
rect 61844 3052 61896 3058
rect 61844 2994 61896 3000
rect 61476 2984 61528 2990
rect 61476 2926 61528 2932
rect 61200 2372 61252 2378
rect 61200 2314 61252 2320
rect 61488 2310 61516 2926
rect 61476 2304 61528 2310
rect 61476 2246 61528 2252
rect 61856 800 61884 2994
rect 62040 2922 62068 3470
rect 62132 3126 62160 31606
rect 63512 5370 63540 36518
rect 63604 35766 63632 37062
rect 63960 36712 64012 36718
rect 63960 36654 64012 36660
rect 63972 36582 64000 36654
rect 63960 36576 64012 36582
rect 63960 36518 64012 36524
rect 63684 36100 63736 36106
rect 63684 36042 63736 36048
rect 63868 36100 63920 36106
rect 63868 36042 63920 36048
rect 63592 35760 63644 35766
rect 63592 35702 63644 35708
rect 63696 35086 63724 36042
rect 63880 35698 63908 36042
rect 63868 35692 63920 35698
rect 63868 35634 63920 35640
rect 63684 35080 63736 35086
rect 63684 35022 63736 35028
rect 64064 5914 64092 37062
rect 64156 35154 64184 37198
rect 64236 36780 64288 36786
rect 64236 36722 64288 36728
rect 64144 35148 64196 35154
rect 64144 35090 64196 35096
rect 64248 34950 64276 36722
rect 64340 36378 64368 39200
rect 64696 38344 64748 38350
rect 64696 38286 64748 38292
rect 64420 37800 64472 37806
rect 64420 37742 64472 37748
rect 64432 36786 64460 37742
rect 64420 36780 64472 36786
rect 64420 36722 64472 36728
rect 64604 36780 64656 36786
rect 64604 36722 64656 36728
rect 64328 36372 64380 36378
rect 64328 36314 64380 36320
rect 64432 35834 64460 36722
rect 64616 36242 64644 36722
rect 64604 36236 64656 36242
rect 64604 36178 64656 36184
rect 64708 36174 64736 38286
rect 65064 37392 65116 37398
rect 65064 37334 65116 37340
rect 64788 37256 64840 37262
rect 64786 37224 64788 37233
rect 64880 37256 64932 37262
rect 64840 37224 64842 37233
rect 64880 37198 64932 37204
rect 64970 37224 65026 37233
rect 64786 37159 64842 37168
rect 64788 36916 64840 36922
rect 64788 36858 64840 36864
rect 64800 36666 64828 36858
rect 64892 36854 64920 37198
rect 64970 37159 65026 37168
rect 64880 36848 64932 36854
rect 64880 36790 64932 36796
rect 64800 36638 64920 36666
rect 64984 36650 65012 37159
rect 65076 36718 65104 37334
rect 65156 37324 65208 37330
rect 65156 37266 65208 37272
rect 65064 36712 65116 36718
rect 65064 36654 65116 36660
rect 64892 36582 64920 36638
rect 64972 36644 65024 36650
rect 64972 36586 65024 36592
rect 64788 36576 64840 36582
rect 64788 36518 64840 36524
rect 64880 36576 64932 36582
rect 64880 36518 64932 36524
rect 64800 36378 64828 36518
rect 64788 36372 64840 36378
rect 64788 36314 64840 36320
rect 64696 36168 64748 36174
rect 64696 36110 64748 36116
rect 64708 35834 64736 36110
rect 64788 36032 64840 36038
rect 64788 35974 64840 35980
rect 64420 35828 64472 35834
rect 64420 35770 64472 35776
rect 64696 35828 64748 35834
rect 64696 35770 64748 35776
rect 64800 35698 64828 35974
rect 64788 35692 64840 35698
rect 64788 35634 64840 35640
rect 64236 34944 64288 34950
rect 64236 34886 64288 34892
rect 64052 5908 64104 5914
rect 64052 5850 64104 5856
rect 63500 5364 63552 5370
rect 63500 5306 63552 5312
rect 63316 4684 63368 4690
rect 63316 4626 63368 4632
rect 62212 4616 62264 4622
rect 62212 4558 62264 4564
rect 62224 4146 62252 4558
rect 62304 4480 62356 4486
rect 62304 4422 62356 4428
rect 62212 4140 62264 4146
rect 62212 4082 62264 4088
rect 62120 3120 62172 3126
rect 62120 3062 62172 3068
rect 62028 2916 62080 2922
rect 62028 2858 62080 2864
rect 62316 2446 62344 4422
rect 63328 4146 63356 4626
rect 63408 4480 63460 4486
rect 63408 4422 63460 4428
rect 63420 4282 63448 4422
rect 63408 4276 63460 4282
rect 63408 4218 63460 4224
rect 63316 4140 63368 4146
rect 63316 4082 63368 4088
rect 63224 3936 63276 3942
rect 63224 3878 63276 3884
rect 62580 3596 62632 3602
rect 62580 3538 62632 3544
rect 62592 3398 62620 3538
rect 62580 3392 62632 3398
rect 62580 3334 62632 3340
rect 62304 2440 62356 2446
rect 62304 2382 62356 2388
rect 63236 800 63264 3878
rect 63512 3602 63540 5306
rect 63868 4072 63920 4078
rect 63868 4014 63920 4020
rect 63880 3602 63908 4014
rect 63960 4004 64012 4010
rect 63960 3946 64012 3952
rect 63500 3596 63552 3602
rect 63500 3538 63552 3544
rect 63868 3596 63920 3602
rect 63868 3538 63920 3544
rect 63500 3392 63552 3398
rect 63500 3334 63552 3340
rect 63512 2378 63540 3334
rect 63592 3052 63644 3058
rect 63592 2994 63644 3000
rect 63604 2650 63632 2994
rect 63880 2990 63908 3538
rect 63868 2984 63920 2990
rect 63868 2926 63920 2932
rect 63592 2644 63644 2650
rect 63592 2586 63644 2592
rect 63972 2378 64000 3946
rect 64064 3126 64092 5850
rect 64328 5024 64380 5030
rect 64328 4966 64380 4972
rect 64340 3126 64368 4966
rect 64420 4480 64472 4486
rect 64420 4422 64472 4428
rect 64432 4282 64460 4422
rect 64420 4276 64472 4282
rect 64420 4218 64472 4224
rect 64800 3126 64828 35634
rect 65168 35578 65196 37266
rect 65260 35698 65288 39200
rect 65654 37564 65962 37573
rect 65654 37562 65660 37564
rect 65716 37562 65740 37564
rect 65796 37562 65820 37564
rect 65876 37562 65900 37564
rect 65956 37562 65962 37564
rect 65716 37510 65718 37562
rect 65898 37510 65900 37562
rect 65654 37508 65660 37510
rect 65716 37508 65740 37510
rect 65796 37508 65820 37510
rect 65876 37508 65900 37510
rect 65956 37508 65962 37510
rect 65654 37499 65962 37508
rect 65432 37324 65484 37330
rect 65432 37266 65484 37272
rect 65340 36848 65392 36854
rect 65340 36790 65392 36796
rect 65352 36174 65380 36790
rect 65340 36168 65392 36174
rect 65340 36110 65392 36116
rect 65248 35692 65300 35698
rect 65248 35634 65300 35640
rect 65168 35550 65288 35578
rect 65260 35086 65288 35550
rect 65352 35154 65380 36110
rect 65444 36106 65472 37266
rect 65524 37256 65576 37262
rect 65524 37198 65576 37204
rect 65798 37224 65854 37233
rect 65536 36854 65564 37198
rect 65798 37159 65854 37168
rect 65524 36848 65576 36854
rect 65524 36790 65576 36796
rect 65812 36718 65840 37159
rect 65984 37120 66036 37126
rect 65984 37062 66036 37068
rect 65800 36712 65852 36718
rect 65536 36638 65748 36666
rect 65800 36654 65852 36660
rect 65432 36100 65484 36106
rect 65432 36042 65484 36048
rect 65340 35148 65392 35154
rect 65340 35090 65392 35096
rect 65248 35080 65300 35086
rect 65246 35048 65248 35057
rect 65300 35048 65302 35057
rect 65246 34983 65302 34992
rect 65536 5914 65564 36638
rect 65720 36582 65748 36638
rect 65708 36576 65760 36582
rect 65708 36518 65760 36524
rect 65654 36476 65962 36485
rect 65654 36474 65660 36476
rect 65716 36474 65740 36476
rect 65796 36474 65820 36476
rect 65876 36474 65900 36476
rect 65956 36474 65962 36476
rect 65716 36422 65718 36474
rect 65898 36422 65900 36474
rect 65654 36420 65660 36422
rect 65716 36420 65740 36422
rect 65796 36420 65820 36422
rect 65876 36420 65900 36422
rect 65956 36420 65962 36422
rect 65654 36411 65962 36420
rect 65654 35388 65962 35397
rect 65654 35386 65660 35388
rect 65716 35386 65740 35388
rect 65796 35386 65820 35388
rect 65876 35386 65900 35388
rect 65956 35386 65962 35388
rect 65716 35334 65718 35386
rect 65898 35334 65900 35386
rect 65654 35332 65660 35334
rect 65716 35332 65740 35334
rect 65796 35332 65820 35334
rect 65876 35332 65900 35334
rect 65956 35332 65962 35334
rect 65654 35323 65962 35332
rect 65654 34300 65962 34309
rect 65654 34298 65660 34300
rect 65716 34298 65740 34300
rect 65796 34298 65820 34300
rect 65876 34298 65900 34300
rect 65956 34298 65962 34300
rect 65716 34246 65718 34298
rect 65898 34246 65900 34298
rect 65654 34244 65660 34246
rect 65716 34244 65740 34246
rect 65796 34244 65820 34246
rect 65876 34244 65900 34246
rect 65956 34244 65962 34246
rect 65654 34235 65962 34244
rect 65654 33212 65962 33221
rect 65654 33210 65660 33212
rect 65716 33210 65740 33212
rect 65796 33210 65820 33212
rect 65876 33210 65900 33212
rect 65956 33210 65962 33212
rect 65716 33158 65718 33210
rect 65898 33158 65900 33210
rect 65654 33156 65660 33158
rect 65716 33156 65740 33158
rect 65796 33156 65820 33158
rect 65876 33156 65900 33158
rect 65956 33156 65962 33158
rect 65654 33147 65962 33156
rect 65654 32124 65962 32133
rect 65654 32122 65660 32124
rect 65716 32122 65740 32124
rect 65796 32122 65820 32124
rect 65876 32122 65900 32124
rect 65956 32122 65962 32124
rect 65716 32070 65718 32122
rect 65898 32070 65900 32122
rect 65654 32068 65660 32070
rect 65716 32068 65740 32070
rect 65796 32068 65820 32070
rect 65876 32068 65900 32070
rect 65956 32068 65962 32070
rect 65654 32059 65962 32068
rect 65996 31754 66024 37062
rect 66180 36904 66208 39200
rect 66536 38140 66588 38146
rect 66536 38082 66588 38088
rect 66260 37392 66312 37398
rect 66260 37334 66312 37340
rect 66272 37194 66300 37334
rect 66260 37188 66312 37194
rect 66260 37130 66312 37136
rect 66260 36916 66312 36922
rect 66180 36876 66260 36904
rect 66260 36858 66312 36864
rect 66548 36786 66576 38082
rect 66812 37120 66864 37126
rect 66812 37062 66864 37068
rect 66536 36780 66588 36786
rect 66536 36722 66588 36728
rect 66260 36576 66312 36582
rect 66260 36518 66312 36524
rect 66272 36378 66300 36518
rect 66260 36372 66312 36378
rect 66260 36314 66312 36320
rect 66076 36100 66128 36106
rect 66076 36042 66128 36048
rect 66088 33998 66116 36042
rect 66444 36032 66496 36038
rect 66442 36000 66444 36009
rect 66496 36000 66498 36009
rect 66442 35935 66498 35944
rect 66548 35834 66576 36722
rect 66536 35828 66588 35834
rect 66536 35770 66588 35776
rect 66076 33992 66128 33998
rect 66076 33934 66128 33940
rect 65996 31726 66116 31754
rect 65654 31036 65962 31045
rect 65654 31034 65660 31036
rect 65716 31034 65740 31036
rect 65796 31034 65820 31036
rect 65876 31034 65900 31036
rect 65956 31034 65962 31036
rect 65716 30982 65718 31034
rect 65898 30982 65900 31034
rect 65654 30980 65660 30982
rect 65716 30980 65740 30982
rect 65796 30980 65820 30982
rect 65876 30980 65900 30982
rect 65956 30980 65962 30982
rect 65654 30971 65962 30980
rect 65654 29948 65962 29957
rect 65654 29946 65660 29948
rect 65716 29946 65740 29948
rect 65796 29946 65820 29948
rect 65876 29946 65900 29948
rect 65956 29946 65962 29948
rect 65716 29894 65718 29946
rect 65898 29894 65900 29946
rect 65654 29892 65660 29894
rect 65716 29892 65740 29894
rect 65796 29892 65820 29894
rect 65876 29892 65900 29894
rect 65956 29892 65962 29894
rect 65654 29883 65962 29892
rect 65654 28860 65962 28869
rect 65654 28858 65660 28860
rect 65716 28858 65740 28860
rect 65796 28858 65820 28860
rect 65876 28858 65900 28860
rect 65956 28858 65962 28860
rect 65716 28806 65718 28858
rect 65898 28806 65900 28858
rect 65654 28804 65660 28806
rect 65716 28804 65740 28806
rect 65796 28804 65820 28806
rect 65876 28804 65900 28806
rect 65956 28804 65962 28806
rect 65654 28795 65962 28804
rect 65654 27772 65962 27781
rect 65654 27770 65660 27772
rect 65716 27770 65740 27772
rect 65796 27770 65820 27772
rect 65876 27770 65900 27772
rect 65956 27770 65962 27772
rect 65716 27718 65718 27770
rect 65898 27718 65900 27770
rect 65654 27716 65660 27718
rect 65716 27716 65740 27718
rect 65796 27716 65820 27718
rect 65876 27716 65900 27718
rect 65956 27716 65962 27718
rect 65654 27707 65962 27716
rect 65654 26684 65962 26693
rect 65654 26682 65660 26684
rect 65716 26682 65740 26684
rect 65796 26682 65820 26684
rect 65876 26682 65900 26684
rect 65956 26682 65962 26684
rect 65716 26630 65718 26682
rect 65898 26630 65900 26682
rect 65654 26628 65660 26630
rect 65716 26628 65740 26630
rect 65796 26628 65820 26630
rect 65876 26628 65900 26630
rect 65956 26628 65962 26630
rect 65654 26619 65962 26628
rect 65654 25596 65962 25605
rect 65654 25594 65660 25596
rect 65716 25594 65740 25596
rect 65796 25594 65820 25596
rect 65876 25594 65900 25596
rect 65956 25594 65962 25596
rect 65716 25542 65718 25594
rect 65898 25542 65900 25594
rect 65654 25540 65660 25542
rect 65716 25540 65740 25542
rect 65796 25540 65820 25542
rect 65876 25540 65900 25542
rect 65956 25540 65962 25542
rect 65654 25531 65962 25540
rect 65654 24508 65962 24517
rect 65654 24506 65660 24508
rect 65716 24506 65740 24508
rect 65796 24506 65820 24508
rect 65876 24506 65900 24508
rect 65956 24506 65962 24508
rect 65716 24454 65718 24506
rect 65898 24454 65900 24506
rect 65654 24452 65660 24454
rect 65716 24452 65740 24454
rect 65796 24452 65820 24454
rect 65876 24452 65900 24454
rect 65956 24452 65962 24454
rect 65654 24443 65962 24452
rect 65654 23420 65962 23429
rect 65654 23418 65660 23420
rect 65716 23418 65740 23420
rect 65796 23418 65820 23420
rect 65876 23418 65900 23420
rect 65956 23418 65962 23420
rect 65716 23366 65718 23418
rect 65898 23366 65900 23418
rect 65654 23364 65660 23366
rect 65716 23364 65740 23366
rect 65796 23364 65820 23366
rect 65876 23364 65900 23366
rect 65956 23364 65962 23366
rect 65654 23355 65962 23364
rect 65654 22332 65962 22341
rect 65654 22330 65660 22332
rect 65716 22330 65740 22332
rect 65796 22330 65820 22332
rect 65876 22330 65900 22332
rect 65956 22330 65962 22332
rect 65716 22278 65718 22330
rect 65898 22278 65900 22330
rect 65654 22276 65660 22278
rect 65716 22276 65740 22278
rect 65796 22276 65820 22278
rect 65876 22276 65900 22278
rect 65956 22276 65962 22278
rect 65654 22267 65962 22276
rect 65654 21244 65962 21253
rect 65654 21242 65660 21244
rect 65716 21242 65740 21244
rect 65796 21242 65820 21244
rect 65876 21242 65900 21244
rect 65956 21242 65962 21244
rect 65716 21190 65718 21242
rect 65898 21190 65900 21242
rect 65654 21188 65660 21190
rect 65716 21188 65740 21190
rect 65796 21188 65820 21190
rect 65876 21188 65900 21190
rect 65956 21188 65962 21190
rect 65654 21179 65962 21188
rect 65654 20156 65962 20165
rect 65654 20154 65660 20156
rect 65716 20154 65740 20156
rect 65796 20154 65820 20156
rect 65876 20154 65900 20156
rect 65956 20154 65962 20156
rect 65716 20102 65718 20154
rect 65898 20102 65900 20154
rect 65654 20100 65660 20102
rect 65716 20100 65740 20102
rect 65796 20100 65820 20102
rect 65876 20100 65900 20102
rect 65956 20100 65962 20102
rect 65654 20091 65962 20100
rect 65654 19068 65962 19077
rect 65654 19066 65660 19068
rect 65716 19066 65740 19068
rect 65796 19066 65820 19068
rect 65876 19066 65900 19068
rect 65956 19066 65962 19068
rect 65716 19014 65718 19066
rect 65898 19014 65900 19066
rect 65654 19012 65660 19014
rect 65716 19012 65740 19014
rect 65796 19012 65820 19014
rect 65876 19012 65900 19014
rect 65956 19012 65962 19014
rect 65654 19003 65962 19012
rect 65654 17980 65962 17989
rect 65654 17978 65660 17980
rect 65716 17978 65740 17980
rect 65796 17978 65820 17980
rect 65876 17978 65900 17980
rect 65956 17978 65962 17980
rect 65716 17926 65718 17978
rect 65898 17926 65900 17978
rect 65654 17924 65660 17926
rect 65716 17924 65740 17926
rect 65796 17924 65820 17926
rect 65876 17924 65900 17926
rect 65956 17924 65962 17926
rect 65654 17915 65962 17924
rect 65654 16892 65962 16901
rect 65654 16890 65660 16892
rect 65716 16890 65740 16892
rect 65796 16890 65820 16892
rect 65876 16890 65900 16892
rect 65956 16890 65962 16892
rect 65716 16838 65718 16890
rect 65898 16838 65900 16890
rect 65654 16836 65660 16838
rect 65716 16836 65740 16838
rect 65796 16836 65820 16838
rect 65876 16836 65900 16838
rect 65956 16836 65962 16838
rect 65654 16827 65962 16836
rect 65654 15804 65962 15813
rect 65654 15802 65660 15804
rect 65716 15802 65740 15804
rect 65796 15802 65820 15804
rect 65876 15802 65900 15804
rect 65956 15802 65962 15804
rect 65716 15750 65718 15802
rect 65898 15750 65900 15802
rect 65654 15748 65660 15750
rect 65716 15748 65740 15750
rect 65796 15748 65820 15750
rect 65876 15748 65900 15750
rect 65956 15748 65962 15750
rect 65654 15739 65962 15748
rect 65654 14716 65962 14725
rect 65654 14714 65660 14716
rect 65716 14714 65740 14716
rect 65796 14714 65820 14716
rect 65876 14714 65900 14716
rect 65956 14714 65962 14716
rect 65716 14662 65718 14714
rect 65898 14662 65900 14714
rect 65654 14660 65660 14662
rect 65716 14660 65740 14662
rect 65796 14660 65820 14662
rect 65876 14660 65900 14662
rect 65956 14660 65962 14662
rect 65654 14651 65962 14660
rect 65654 13628 65962 13637
rect 65654 13626 65660 13628
rect 65716 13626 65740 13628
rect 65796 13626 65820 13628
rect 65876 13626 65900 13628
rect 65956 13626 65962 13628
rect 65716 13574 65718 13626
rect 65898 13574 65900 13626
rect 65654 13572 65660 13574
rect 65716 13572 65740 13574
rect 65796 13572 65820 13574
rect 65876 13572 65900 13574
rect 65956 13572 65962 13574
rect 65654 13563 65962 13572
rect 65654 12540 65962 12549
rect 65654 12538 65660 12540
rect 65716 12538 65740 12540
rect 65796 12538 65820 12540
rect 65876 12538 65900 12540
rect 65956 12538 65962 12540
rect 65716 12486 65718 12538
rect 65898 12486 65900 12538
rect 65654 12484 65660 12486
rect 65716 12484 65740 12486
rect 65796 12484 65820 12486
rect 65876 12484 65900 12486
rect 65956 12484 65962 12486
rect 65654 12475 65962 12484
rect 65654 11452 65962 11461
rect 65654 11450 65660 11452
rect 65716 11450 65740 11452
rect 65796 11450 65820 11452
rect 65876 11450 65900 11452
rect 65956 11450 65962 11452
rect 65716 11398 65718 11450
rect 65898 11398 65900 11450
rect 65654 11396 65660 11398
rect 65716 11396 65740 11398
rect 65796 11396 65820 11398
rect 65876 11396 65900 11398
rect 65956 11396 65962 11398
rect 65654 11387 65962 11396
rect 65654 10364 65962 10373
rect 65654 10362 65660 10364
rect 65716 10362 65740 10364
rect 65796 10362 65820 10364
rect 65876 10362 65900 10364
rect 65956 10362 65962 10364
rect 65716 10310 65718 10362
rect 65898 10310 65900 10362
rect 65654 10308 65660 10310
rect 65716 10308 65740 10310
rect 65796 10308 65820 10310
rect 65876 10308 65900 10310
rect 65956 10308 65962 10310
rect 65654 10299 65962 10308
rect 65654 9276 65962 9285
rect 65654 9274 65660 9276
rect 65716 9274 65740 9276
rect 65796 9274 65820 9276
rect 65876 9274 65900 9276
rect 65956 9274 65962 9276
rect 65716 9222 65718 9274
rect 65898 9222 65900 9274
rect 65654 9220 65660 9222
rect 65716 9220 65740 9222
rect 65796 9220 65820 9222
rect 65876 9220 65900 9222
rect 65956 9220 65962 9222
rect 65654 9211 65962 9220
rect 65654 8188 65962 8197
rect 65654 8186 65660 8188
rect 65716 8186 65740 8188
rect 65796 8186 65820 8188
rect 65876 8186 65900 8188
rect 65956 8186 65962 8188
rect 65716 8134 65718 8186
rect 65898 8134 65900 8186
rect 65654 8132 65660 8134
rect 65716 8132 65740 8134
rect 65796 8132 65820 8134
rect 65876 8132 65900 8134
rect 65956 8132 65962 8134
rect 65654 8123 65962 8132
rect 65654 7100 65962 7109
rect 65654 7098 65660 7100
rect 65716 7098 65740 7100
rect 65796 7098 65820 7100
rect 65876 7098 65900 7100
rect 65956 7098 65962 7100
rect 65716 7046 65718 7098
rect 65898 7046 65900 7098
rect 65654 7044 65660 7046
rect 65716 7044 65740 7046
rect 65796 7044 65820 7046
rect 65876 7044 65900 7046
rect 65956 7044 65962 7046
rect 65654 7035 65962 7044
rect 65654 6012 65962 6021
rect 65654 6010 65660 6012
rect 65716 6010 65740 6012
rect 65796 6010 65820 6012
rect 65876 6010 65900 6012
rect 65956 6010 65962 6012
rect 65716 5958 65718 6010
rect 65898 5958 65900 6010
rect 65654 5956 65660 5958
rect 65716 5956 65740 5958
rect 65796 5956 65820 5958
rect 65876 5956 65900 5958
rect 65956 5956 65962 5958
rect 65654 5947 65962 5956
rect 65524 5908 65576 5914
rect 65524 5850 65576 5856
rect 65156 5568 65208 5574
rect 65156 5510 65208 5516
rect 64880 5024 64932 5030
rect 64880 4966 64932 4972
rect 64892 3534 64920 4966
rect 65064 4616 65116 4622
rect 65064 4558 65116 4564
rect 65076 3738 65104 4558
rect 65168 4078 65196 5510
rect 65340 5024 65392 5030
rect 65340 4966 65392 4972
rect 65248 4480 65300 4486
rect 65248 4422 65300 4428
rect 65156 4072 65208 4078
rect 65156 4014 65208 4020
rect 65064 3732 65116 3738
rect 65064 3674 65116 3680
rect 64880 3528 64932 3534
rect 64880 3470 64932 3476
rect 64052 3120 64104 3126
rect 64052 3062 64104 3068
rect 64328 3120 64380 3126
rect 64328 3062 64380 3068
rect 64604 3120 64656 3126
rect 64604 3062 64656 3068
rect 64788 3120 64840 3126
rect 64788 3062 64840 3068
rect 63500 2372 63552 2378
rect 63500 2314 63552 2320
rect 63960 2372 64012 2378
rect 63960 2314 64012 2320
rect 64616 800 64644 3062
rect 64892 1970 64920 3470
rect 65064 3460 65116 3466
rect 65064 3402 65116 3408
rect 65076 2990 65104 3402
rect 65168 3194 65196 4014
rect 65156 3188 65208 3194
rect 65156 3130 65208 3136
rect 65064 2984 65116 2990
rect 65064 2926 65116 2932
rect 65076 2650 65104 2926
rect 65064 2644 65116 2650
rect 65064 2586 65116 2592
rect 65260 2378 65288 4422
rect 65352 4010 65380 4966
rect 65536 4026 65564 5850
rect 66088 5370 66116 31726
rect 66824 8362 66852 37062
rect 67100 36786 67128 39200
rect 67548 37732 67600 37738
rect 67548 37674 67600 37680
rect 67560 37398 67588 37674
rect 67548 37392 67600 37398
rect 67548 37334 67600 37340
rect 67824 37392 67876 37398
rect 67824 37334 67876 37340
rect 67272 37256 67324 37262
rect 67272 37198 67324 37204
rect 67088 36780 67140 36786
rect 67088 36722 67140 36728
rect 67100 36378 67128 36722
rect 67088 36372 67140 36378
rect 67088 36314 67140 36320
rect 67284 35834 67312 37198
rect 67732 37188 67784 37194
rect 67732 37130 67784 37136
rect 67744 36242 67772 37130
rect 67836 36310 67864 37334
rect 68020 36378 68048 39200
rect 68376 37732 68428 37738
rect 68376 37674 68428 37680
rect 68008 36372 68060 36378
rect 68008 36314 68060 36320
rect 67824 36304 67876 36310
rect 67824 36246 67876 36252
rect 67732 36236 67784 36242
rect 67732 36178 67784 36184
rect 68388 36174 68416 37674
rect 68558 37224 68614 37233
rect 68558 37159 68560 37168
rect 68612 37159 68614 37168
rect 68560 37130 68612 37136
rect 68192 36168 68244 36174
rect 68192 36110 68244 36116
rect 68376 36168 68428 36174
rect 68376 36110 68428 36116
rect 68204 36009 68232 36110
rect 68190 36000 68246 36009
rect 68190 35935 68246 35944
rect 68388 35834 68416 36110
rect 67272 35828 67324 35834
rect 67272 35770 67324 35776
rect 68376 35828 68428 35834
rect 68376 35770 68428 35776
rect 68572 35154 68600 37130
rect 68664 36786 68692 39238
rect 68926 39200 68982 40000
rect 69846 39200 69902 40000
rect 70766 39200 70822 40000
rect 71686 39200 71742 40000
rect 72606 39200 72662 40000
rect 73526 39200 73582 40000
rect 73620 39364 73672 39370
rect 73620 39306 73672 39312
rect 68652 36780 68704 36786
rect 68652 36722 68704 36728
rect 68940 36174 68968 39200
rect 69860 37126 69888 39200
rect 70492 37256 70544 37262
rect 70492 37198 70544 37204
rect 69020 37120 69072 37126
rect 69020 37062 69072 37068
rect 69848 37120 69900 37126
rect 69848 37062 69900 37068
rect 68928 36168 68980 36174
rect 68928 36110 68980 36116
rect 68560 35148 68612 35154
rect 68560 35090 68612 35096
rect 69032 34626 69060 37062
rect 69204 36780 69256 36786
rect 69204 36722 69256 36728
rect 69664 36780 69716 36786
rect 69664 36722 69716 36728
rect 69216 35494 69244 36722
rect 69204 35488 69256 35494
rect 69204 35430 69256 35436
rect 69032 34598 69152 34626
rect 69020 34536 69072 34542
rect 69020 34478 69072 34484
rect 66812 8356 66864 8362
rect 66812 8298 66864 8304
rect 67640 8356 67692 8362
rect 67640 8298 67692 8304
rect 66076 5364 66128 5370
rect 66076 5306 66128 5312
rect 65654 4924 65962 4933
rect 65654 4922 65660 4924
rect 65716 4922 65740 4924
rect 65796 4922 65820 4924
rect 65876 4922 65900 4924
rect 65956 4922 65962 4924
rect 65716 4870 65718 4922
rect 65898 4870 65900 4922
rect 65654 4868 65660 4870
rect 65716 4868 65740 4870
rect 65796 4868 65820 4870
rect 65876 4868 65900 4870
rect 65956 4868 65962 4870
rect 65654 4859 65962 4868
rect 66088 4214 66116 5306
rect 67652 4826 67680 8298
rect 68192 5296 68244 5302
rect 68192 5238 68244 5244
rect 68204 4826 68232 5238
rect 68928 5024 68980 5030
rect 68928 4966 68980 4972
rect 67640 4820 67692 4826
rect 67640 4762 67692 4768
rect 68192 4820 68244 4826
rect 68192 4762 68244 4768
rect 66168 4752 66220 4758
rect 66168 4694 66220 4700
rect 66536 4752 66588 4758
rect 66536 4694 66588 4700
rect 66076 4208 66128 4214
rect 66076 4150 66128 4156
rect 65340 4004 65392 4010
rect 65340 3946 65392 3952
rect 65444 3998 65564 4026
rect 65444 3602 65472 3998
rect 65524 3936 65576 3942
rect 65524 3878 65576 3884
rect 65432 3596 65484 3602
rect 65432 3538 65484 3544
rect 65536 3126 65564 3878
rect 65654 3836 65962 3845
rect 65654 3834 65660 3836
rect 65716 3834 65740 3836
rect 65796 3834 65820 3836
rect 65876 3834 65900 3836
rect 65956 3834 65962 3836
rect 65716 3782 65718 3834
rect 65898 3782 65900 3834
rect 65654 3780 65660 3782
rect 65716 3780 65740 3782
rect 65796 3780 65820 3782
rect 65876 3780 65900 3782
rect 65956 3780 65962 3782
rect 65654 3771 65962 3780
rect 66180 3534 66208 4694
rect 66548 4146 66576 4694
rect 66536 4140 66588 4146
rect 66456 4100 66536 4128
rect 66456 3738 66484 4100
rect 66536 4082 66588 4088
rect 67364 4004 67416 4010
rect 67364 3946 67416 3952
rect 66536 3936 66588 3942
rect 66536 3878 66588 3884
rect 66444 3732 66496 3738
rect 66444 3674 66496 3680
rect 66456 3602 66484 3674
rect 66444 3596 66496 3602
rect 66444 3538 66496 3544
rect 66168 3528 66220 3534
rect 66168 3470 66220 3476
rect 66180 3194 66208 3470
rect 66168 3188 66220 3194
rect 66168 3130 66220 3136
rect 65524 3120 65576 3126
rect 65524 3062 65576 3068
rect 65654 2748 65962 2757
rect 65654 2746 65660 2748
rect 65716 2746 65740 2748
rect 65796 2746 65820 2748
rect 65876 2746 65900 2748
rect 65956 2746 65962 2748
rect 65716 2694 65718 2746
rect 65898 2694 65900 2746
rect 65654 2692 65660 2694
rect 65716 2692 65740 2694
rect 65796 2692 65820 2694
rect 65876 2692 65900 2694
rect 65956 2692 65962 2694
rect 65654 2683 65962 2692
rect 66548 2378 66576 3878
rect 67376 3398 67404 3946
rect 67652 3534 67680 4762
rect 68652 4480 68704 4486
rect 68652 4422 68704 4428
rect 68664 4282 68692 4422
rect 68284 4276 68336 4282
rect 68284 4218 68336 4224
rect 68652 4276 68704 4282
rect 68652 4218 68704 4224
rect 68296 3602 68324 4218
rect 68836 4140 68888 4146
rect 68836 4082 68888 4088
rect 68468 3936 68520 3942
rect 68468 3878 68520 3884
rect 68008 3596 68060 3602
rect 68008 3538 68060 3544
rect 68284 3596 68336 3602
rect 68284 3538 68336 3544
rect 67640 3528 67692 3534
rect 67640 3470 67692 3476
rect 66812 3392 66864 3398
rect 66812 3334 66864 3340
rect 67272 3392 67324 3398
rect 67272 3334 67324 3340
rect 67364 3392 67416 3398
rect 67364 3334 67416 3340
rect 66824 3058 66852 3334
rect 67284 3126 67312 3334
rect 67272 3120 67324 3126
rect 67272 3062 67324 3068
rect 66812 3052 66864 3058
rect 66812 2994 66864 3000
rect 67376 2938 67404 3334
rect 68020 3058 68048 3538
rect 68480 3534 68508 3878
rect 68848 3738 68876 4082
rect 68836 3732 68888 3738
rect 68836 3674 68888 3680
rect 68468 3528 68520 3534
rect 68466 3496 68468 3505
rect 68520 3496 68522 3505
rect 68466 3431 68522 3440
rect 68008 3052 68060 3058
rect 68008 2994 68060 3000
rect 68836 3052 68888 3058
rect 68836 2994 68888 3000
rect 67284 2910 67404 2938
rect 67284 2854 67312 2910
rect 67272 2848 67324 2854
rect 67272 2790 67324 2796
rect 67364 2848 67416 2854
rect 67364 2790 67416 2796
rect 65248 2372 65300 2378
rect 65248 2314 65300 2320
rect 66536 2372 66588 2378
rect 66536 2314 66588 2320
rect 64880 1964 64932 1970
rect 64880 1906 64932 1912
rect 67376 800 67404 2790
rect 68848 2582 68876 2994
rect 68836 2576 68888 2582
rect 68836 2518 68888 2524
rect 68940 2378 68968 4966
rect 69032 2650 69060 34478
rect 69124 5370 69152 34598
rect 69216 34542 69244 35430
rect 69204 34536 69256 34542
rect 69204 34478 69256 34484
rect 69676 33930 69704 36722
rect 70504 36394 70532 37198
rect 70780 36786 70808 39200
rect 70860 37324 70912 37330
rect 70860 37266 70912 37272
rect 70768 36780 70820 36786
rect 70768 36722 70820 36728
rect 70872 36582 70900 37266
rect 71136 37188 71188 37194
rect 71136 37130 71188 37136
rect 71596 37188 71648 37194
rect 71596 37130 71648 37136
rect 70860 36576 70912 36582
rect 70860 36518 70912 36524
rect 71044 36576 71096 36582
rect 71044 36518 71096 36524
rect 70412 36378 70532 36394
rect 70400 36372 70532 36378
rect 70452 36366 70532 36372
rect 70400 36314 70452 36320
rect 70504 35766 70532 36366
rect 70872 36310 70900 36518
rect 70860 36304 70912 36310
rect 70860 36246 70912 36252
rect 71056 36242 71084 36518
rect 71148 36310 71176 37130
rect 71320 37120 71372 37126
rect 71320 37062 71372 37068
rect 71504 37120 71556 37126
rect 71504 37062 71556 37068
rect 71332 36650 71360 37062
rect 71320 36644 71372 36650
rect 71320 36586 71372 36592
rect 71136 36304 71188 36310
rect 71136 36246 71188 36252
rect 71044 36236 71096 36242
rect 71044 36178 71096 36184
rect 70492 35760 70544 35766
rect 70492 35702 70544 35708
rect 69664 33924 69716 33930
rect 69664 33866 69716 33872
rect 71516 31754 71544 37062
rect 71608 36938 71636 37130
rect 71700 37108 71728 39200
rect 72332 37460 72384 37466
rect 72332 37402 72384 37408
rect 71780 37120 71832 37126
rect 71700 37080 71780 37108
rect 71780 37062 71832 37068
rect 71608 36910 71728 36938
rect 71700 36582 71728 36910
rect 71688 36576 71740 36582
rect 71688 36518 71740 36524
rect 71700 35193 71728 36518
rect 72344 36378 72372 37402
rect 72516 37256 72568 37262
rect 72516 37198 72568 37204
rect 72528 36666 72556 37198
rect 72620 36786 72648 39200
rect 73158 37360 73214 37369
rect 73158 37295 73214 37304
rect 72792 36916 72844 36922
rect 73172 36904 73200 37295
rect 73540 37126 73568 39200
rect 73632 37194 73660 39306
rect 74446 39200 74502 40000
rect 75366 39200 75422 40000
rect 76286 39200 76342 40000
rect 77206 39200 77262 40000
rect 78126 39200 78182 40000
rect 78232 39222 78628 39250
rect 73620 37188 73672 37194
rect 73620 37130 73672 37136
rect 73804 37188 73856 37194
rect 73804 37130 73856 37136
rect 73528 37120 73580 37126
rect 73528 37062 73580 37068
rect 72844 36876 73200 36904
rect 72792 36858 72844 36864
rect 72608 36780 72660 36786
rect 72608 36722 72660 36728
rect 72528 36638 72648 36666
rect 73816 36650 73844 37130
rect 72620 36378 72648 36638
rect 73804 36644 73856 36650
rect 73804 36586 73856 36592
rect 73988 36576 74040 36582
rect 73988 36518 74040 36524
rect 72332 36372 72384 36378
rect 72332 36314 72384 36320
rect 72608 36372 72660 36378
rect 72608 36314 72660 36320
rect 71686 35184 71742 35193
rect 71686 35119 71742 35128
rect 72620 33862 72648 36314
rect 74000 36106 74028 36518
rect 74460 36378 74488 39200
rect 75184 39160 75236 39166
rect 75184 39102 75236 39108
rect 75196 37874 75224 39102
rect 75184 37868 75236 37874
rect 75184 37810 75236 37816
rect 74540 37256 74592 37262
rect 74540 37198 74592 37204
rect 74724 37256 74776 37262
rect 74724 37198 74776 37204
rect 74552 36786 74580 37198
rect 74736 36922 74764 37198
rect 75092 37188 75144 37194
rect 75092 37130 75144 37136
rect 74906 36952 74962 36961
rect 74724 36916 74776 36922
rect 74906 36887 74962 36896
rect 74724 36858 74776 36864
rect 74540 36780 74592 36786
rect 74540 36722 74592 36728
rect 74632 36644 74684 36650
rect 74632 36586 74684 36592
rect 74448 36372 74500 36378
rect 74448 36314 74500 36320
rect 74460 36174 74488 36314
rect 74644 36174 74672 36586
rect 74920 36417 74948 36887
rect 74998 36816 75054 36825
rect 74998 36751 75054 36760
rect 75012 36553 75040 36751
rect 74998 36544 75054 36553
rect 74998 36479 75054 36488
rect 74906 36408 74962 36417
rect 74906 36343 74962 36352
rect 74448 36168 74500 36174
rect 74448 36110 74500 36116
rect 74632 36168 74684 36174
rect 74632 36110 74684 36116
rect 75104 36106 75132 37130
rect 75184 36780 75236 36786
rect 75184 36722 75236 36728
rect 73988 36100 74040 36106
rect 73988 36042 74040 36048
rect 75092 36100 75144 36106
rect 75092 36042 75144 36048
rect 75104 35494 75132 36042
rect 75196 36038 75224 36722
rect 75380 36666 75408 39200
rect 75920 37868 75972 37874
rect 75920 37810 75972 37816
rect 75828 37324 75880 37330
rect 75828 37266 75880 37272
rect 75552 37188 75604 37194
rect 75552 37130 75604 37136
rect 75458 36952 75514 36961
rect 75458 36887 75514 36896
rect 75472 36718 75500 36887
rect 75288 36650 75408 36666
rect 75460 36712 75512 36718
rect 75460 36654 75512 36660
rect 75276 36644 75408 36650
rect 75328 36638 75408 36644
rect 75276 36586 75328 36592
rect 75564 36378 75592 37130
rect 75736 37120 75788 37126
rect 75736 37062 75788 37068
rect 75552 36372 75604 36378
rect 75552 36314 75604 36320
rect 75748 36038 75776 37062
rect 75184 36032 75236 36038
rect 75184 35974 75236 35980
rect 75736 36032 75788 36038
rect 75736 35974 75788 35980
rect 75092 35488 75144 35494
rect 75092 35430 75144 35436
rect 72608 33856 72660 33862
rect 72608 33798 72660 33804
rect 71424 31726 71544 31754
rect 69480 5568 69532 5574
rect 69480 5510 69532 5516
rect 69492 5370 69520 5510
rect 69112 5364 69164 5370
rect 69112 5306 69164 5312
rect 69480 5364 69532 5370
rect 69480 5306 69532 5312
rect 69124 3534 69152 5306
rect 69664 5024 69716 5030
rect 69664 4966 69716 4972
rect 70308 5024 70360 5030
rect 70308 4966 70360 4972
rect 69204 4480 69256 4486
rect 69204 4422 69256 4428
rect 69216 4078 69244 4422
rect 69296 4208 69348 4214
rect 69296 4150 69348 4156
rect 69204 4072 69256 4078
rect 69204 4014 69256 4020
rect 69216 3942 69244 4014
rect 69204 3936 69256 3942
rect 69204 3878 69256 3884
rect 69112 3528 69164 3534
rect 69112 3470 69164 3476
rect 69308 3194 69336 4150
rect 69676 3534 69704 4966
rect 69848 4616 69900 4622
rect 69848 4558 69900 4564
rect 69756 4072 69808 4078
rect 69756 4014 69808 4020
rect 69664 3528 69716 3534
rect 69664 3470 69716 3476
rect 69676 3194 69704 3470
rect 69768 3466 69796 4014
rect 69860 3738 69888 4558
rect 70320 4554 70348 4966
rect 70308 4548 70360 4554
rect 70308 4490 70360 4496
rect 69952 3738 70164 3754
rect 69848 3732 69900 3738
rect 69848 3674 69900 3680
rect 69952 3732 70176 3738
rect 69952 3726 70124 3732
rect 69952 3534 69980 3726
rect 70124 3674 70176 3680
rect 69940 3528 69992 3534
rect 69940 3470 69992 3476
rect 70032 3528 70084 3534
rect 70032 3470 70084 3476
rect 69756 3460 69808 3466
rect 69756 3402 69808 3408
rect 69940 3392 69992 3398
rect 69768 3340 69940 3346
rect 69768 3334 69992 3340
rect 69768 3318 69980 3334
rect 69296 3188 69348 3194
rect 69296 3130 69348 3136
rect 69664 3188 69716 3194
rect 69664 3130 69716 3136
rect 69768 3058 69796 3318
rect 70044 3210 70072 3470
rect 70124 3460 70176 3466
rect 70124 3402 70176 3408
rect 69860 3182 70072 3210
rect 69860 3126 69888 3182
rect 69848 3120 69900 3126
rect 70136 3108 70164 3402
rect 69848 3062 69900 3068
rect 70044 3080 70164 3108
rect 69756 3052 69808 3058
rect 69756 2994 69808 3000
rect 69940 2984 69992 2990
rect 69938 2952 69940 2961
rect 69992 2952 69994 2961
rect 70044 2922 70072 3080
rect 69938 2887 69994 2896
rect 70032 2916 70084 2922
rect 70032 2858 70084 2864
rect 70124 2916 70176 2922
rect 70124 2858 70176 2864
rect 70136 2802 70164 2858
rect 70320 2802 70348 4490
rect 70400 4480 70452 4486
rect 70400 4422 70452 4428
rect 70412 3126 70440 4422
rect 71424 4146 71452 31726
rect 75104 24206 75132 35430
rect 75840 34202 75868 37266
rect 75932 35290 75960 37810
rect 76196 37324 76248 37330
rect 76196 37266 76248 37272
rect 76208 36786 76236 37266
rect 76300 36922 76328 39200
rect 77024 37324 77076 37330
rect 77024 37266 77076 37272
rect 76472 37120 76524 37126
rect 76472 37062 76524 37068
rect 76288 36916 76340 36922
rect 76288 36858 76340 36864
rect 76196 36780 76248 36786
rect 76196 36722 76248 36728
rect 76288 36780 76340 36786
rect 76288 36722 76340 36728
rect 76104 36576 76156 36582
rect 76104 36518 76156 36524
rect 76116 36174 76144 36518
rect 76300 36378 76328 36722
rect 76288 36372 76340 36378
rect 76288 36314 76340 36320
rect 76104 36168 76156 36174
rect 76104 36110 76156 36116
rect 75920 35284 75972 35290
rect 75920 35226 75972 35232
rect 75828 34196 75880 34202
rect 75828 34138 75880 34144
rect 73712 24200 73764 24206
rect 73712 24142 73764 24148
rect 75092 24200 75144 24206
rect 75092 24142 75144 24148
rect 71596 4616 71648 4622
rect 71596 4558 71648 4564
rect 71412 4140 71464 4146
rect 71412 4082 71464 4088
rect 71228 3936 71280 3942
rect 71228 3878 71280 3884
rect 71240 3505 71268 3878
rect 71424 3602 71452 4082
rect 71608 3942 71636 4558
rect 72424 4072 72476 4078
rect 72424 4014 72476 4020
rect 72516 4072 72568 4078
rect 72516 4014 72568 4020
rect 71596 3936 71648 3942
rect 71596 3878 71648 3884
rect 71608 3602 71636 3878
rect 71412 3596 71464 3602
rect 71412 3538 71464 3544
rect 71596 3596 71648 3602
rect 71596 3538 71648 3544
rect 71226 3496 71282 3505
rect 71226 3431 71282 3440
rect 70400 3120 70452 3126
rect 70400 3062 70452 3068
rect 70492 3120 70544 3126
rect 70492 3062 70544 3068
rect 70136 2774 70348 2802
rect 70136 2650 70164 2774
rect 69020 2644 69072 2650
rect 69020 2586 69072 2592
rect 69112 2644 69164 2650
rect 69112 2586 69164 2592
rect 70124 2644 70176 2650
rect 70124 2586 70176 2592
rect 69124 2514 69152 2586
rect 70504 2582 70532 3062
rect 71136 2848 71188 2854
rect 71136 2790 71188 2796
rect 70952 2644 71004 2650
rect 70952 2586 71004 2592
rect 70492 2576 70544 2582
rect 70492 2518 70544 2524
rect 70964 2514 70992 2586
rect 69112 2508 69164 2514
rect 69112 2450 69164 2456
rect 70952 2508 71004 2514
rect 70952 2450 71004 2456
rect 71148 2378 71176 2790
rect 68928 2372 68980 2378
rect 68756 2332 68928 2360
rect 67548 2304 67600 2310
rect 67548 2246 67600 2252
rect 67560 1970 67588 2246
rect 67548 1964 67600 1970
rect 67548 1906 67600 1912
rect 68756 800 68784 2332
rect 68928 2314 68980 2320
rect 71136 2372 71188 2378
rect 71136 2314 71188 2320
rect 70952 2304 71004 2310
rect 70952 2246 71004 2252
rect 70964 1902 70992 2246
rect 70952 1896 71004 1902
rect 70952 1838 71004 1844
rect 71240 1766 71268 3431
rect 72436 3058 72464 4014
rect 72528 3194 72556 4014
rect 73528 4004 73580 4010
rect 73528 3946 73580 3952
rect 72700 3392 72752 3398
rect 72700 3334 72752 3340
rect 72884 3392 72936 3398
rect 72884 3334 72936 3340
rect 72516 3188 72568 3194
rect 72516 3130 72568 3136
rect 72424 3052 72476 3058
rect 72424 2994 72476 3000
rect 71504 2916 71556 2922
rect 71504 2858 71556 2864
rect 71228 1760 71280 1766
rect 71228 1702 71280 1708
rect 71516 800 71544 2858
rect 71688 2372 71740 2378
rect 71688 2314 71740 2320
rect 71700 1902 71728 2314
rect 72712 2310 72740 3334
rect 72896 3058 72924 3334
rect 72884 3052 72936 3058
rect 72884 2994 72936 3000
rect 72700 2304 72752 2310
rect 72700 2246 72752 2252
rect 71688 1896 71740 1902
rect 71688 1838 71740 1844
rect 72712 1834 72740 2246
rect 72700 1828 72752 1834
rect 72700 1770 72752 1776
rect 72896 800 72924 2994
rect 73540 2514 73568 3946
rect 73724 3194 73752 24142
rect 76484 5574 76512 37062
rect 76654 36952 76710 36961
rect 77036 36922 77064 37266
rect 77116 37120 77168 37126
rect 77220 37108 77248 39200
rect 78140 39114 78168 39200
rect 78232 39114 78260 39222
rect 78140 39086 78260 39114
rect 77392 37256 77444 37262
rect 77392 37198 77444 37204
rect 77300 37120 77352 37126
rect 77220 37080 77300 37108
rect 77116 37062 77168 37068
rect 77300 37062 77352 37068
rect 77128 36938 77156 37062
rect 76654 36887 76710 36896
rect 77024 36916 77076 36922
rect 76668 36718 76696 36887
rect 77128 36910 77340 36938
rect 77024 36858 77076 36864
rect 76656 36712 76708 36718
rect 76656 36654 76708 36660
rect 76564 36644 76616 36650
rect 76564 36586 76616 36592
rect 76576 36009 76604 36586
rect 77312 36582 77340 36910
rect 77300 36576 77352 36582
rect 77300 36518 77352 36524
rect 77300 36168 77352 36174
rect 77404 36156 77432 37198
rect 78600 36904 78628 39222
rect 79046 39200 79102 40000
rect 79966 39200 80022 40000
rect 80886 39200 80942 40000
rect 81806 39200 81862 40000
rect 81912 39222 82216 39250
rect 79060 37505 79088 39200
rect 79980 38026 80008 39200
rect 79980 37998 80192 38026
rect 79324 37868 79376 37874
rect 79324 37810 79376 37816
rect 79046 37496 79102 37505
rect 79336 37466 79364 37810
rect 79506 37632 79562 37641
rect 79506 37567 79562 37576
rect 79046 37431 79102 37440
rect 79324 37460 79376 37466
rect 79324 37402 79376 37408
rect 79140 37392 79192 37398
rect 79140 37334 79192 37340
rect 79048 37120 79100 37126
rect 79048 37062 79100 37068
rect 78680 36916 78732 36922
rect 78600 36876 78680 36904
rect 78680 36858 78732 36864
rect 78956 36780 79008 36786
rect 78956 36722 79008 36728
rect 77760 36576 77812 36582
rect 77760 36518 77812 36524
rect 77352 36128 77432 36156
rect 77300 36110 77352 36116
rect 76562 36000 76618 36009
rect 76562 35935 76618 35944
rect 77312 35873 77340 36110
rect 77298 35864 77354 35873
rect 77298 35799 77354 35808
rect 77772 33114 77800 36518
rect 78496 36100 78548 36106
rect 78496 36042 78548 36048
rect 77760 33108 77812 33114
rect 77760 33050 77812 33056
rect 78220 5704 78272 5710
rect 78220 5646 78272 5652
rect 75736 5568 75788 5574
rect 75736 5510 75788 5516
rect 76472 5568 76524 5574
rect 76472 5510 76524 5516
rect 77208 5568 77260 5574
rect 77208 5510 77260 5516
rect 75092 4480 75144 4486
rect 75092 4422 75144 4428
rect 74080 3528 74132 3534
rect 74080 3470 74132 3476
rect 74540 3528 74592 3534
rect 74540 3470 74592 3476
rect 73712 3188 73764 3194
rect 73712 3130 73764 3136
rect 74092 2990 74120 3470
rect 74448 3392 74500 3398
rect 74448 3334 74500 3340
rect 74460 3058 74488 3334
rect 74448 3052 74500 3058
rect 74448 2994 74500 3000
rect 74080 2984 74132 2990
rect 74080 2926 74132 2932
rect 73804 2848 73856 2854
rect 73804 2790 73856 2796
rect 73528 2508 73580 2514
rect 73528 2450 73580 2456
rect 73816 2378 73844 2790
rect 74552 2378 74580 3470
rect 75104 3058 75132 4422
rect 75748 4146 75776 5510
rect 75736 4140 75788 4146
rect 75736 4082 75788 4088
rect 75368 3936 75420 3942
rect 75368 3878 75420 3884
rect 75380 3602 75408 3878
rect 75368 3596 75420 3602
rect 75368 3538 75420 3544
rect 75748 3534 75776 4082
rect 77116 4004 77168 4010
rect 77116 3946 77168 3952
rect 76472 3936 76524 3942
rect 76472 3878 76524 3884
rect 76484 3670 76512 3878
rect 76472 3664 76524 3670
rect 76472 3606 76524 3612
rect 75736 3528 75788 3534
rect 75736 3470 75788 3476
rect 75828 3528 75880 3534
rect 75828 3470 75880 3476
rect 75840 3398 75868 3470
rect 76196 3460 76248 3466
rect 76196 3402 76248 3408
rect 75828 3392 75880 3398
rect 75828 3334 75880 3340
rect 75092 3052 75144 3058
rect 75092 2994 75144 3000
rect 75736 3052 75788 3058
rect 75736 2994 75788 3000
rect 75748 2961 75776 2994
rect 75734 2952 75790 2961
rect 75734 2887 75790 2896
rect 75644 2848 75696 2854
rect 75644 2790 75696 2796
rect 73804 2372 73856 2378
rect 73804 2314 73856 2320
rect 74540 2372 74592 2378
rect 74540 2314 74592 2320
rect 75656 800 75684 2790
rect 75840 2446 75868 3334
rect 76208 2990 76236 3402
rect 76380 3392 76432 3398
rect 76380 3334 76432 3340
rect 76196 2984 76248 2990
rect 76196 2926 76248 2932
rect 75828 2440 75880 2446
rect 75828 2382 75880 2388
rect 76392 2378 76420 3334
rect 76484 2854 76512 3606
rect 77128 3602 77156 3946
rect 77116 3596 77168 3602
rect 77116 3538 77168 3544
rect 76564 3528 76616 3534
rect 76564 3470 76616 3476
rect 76576 2854 76604 3470
rect 77220 3194 77248 5510
rect 78232 4826 78260 5646
rect 78508 5574 78536 36042
rect 78968 36038 78996 36722
rect 78956 36032 79008 36038
rect 78956 35974 79008 35980
rect 79060 5710 79088 37062
rect 79152 36786 79180 37334
rect 79520 37330 79548 37567
rect 79508 37324 79560 37330
rect 79560 37284 79640 37312
rect 79508 37266 79560 37272
rect 79140 36780 79192 36786
rect 79140 36722 79192 36728
rect 79140 36032 79192 36038
rect 79140 35974 79192 35980
rect 79152 33658 79180 35974
rect 79508 35624 79560 35630
rect 79508 35566 79560 35572
rect 79520 35290 79548 35566
rect 79612 35290 79640 37284
rect 79966 36952 80022 36961
rect 79966 36887 80022 36896
rect 79784 36576 79836 36582
rect 79784 36518 79836 36524
rect 79508 35284 79560 35290
rect 79508 35226 79560 35232
rect 79600 35284 79652 35290
rect 79600 35226 79652 35232
rect 79140 33652 79192 33658
rect 79140 33594 79192 33600
rect 79796 31770 79824 36518
rect 79980 36378 80008 36887
rect 80164 36378 80192 37998
rect 80244 37868 80296 37874
rect 80244 37810 80296 37816
rect 80256 36922 80284 37810
rect 80426 37496 80482 37505
rect 80426 37431 80482 37440
rect 80440 37262 80468 37431
rect 80796 37324 80848 37330
rect 80796 37266 80848 37272
rect 80428 37256 80480 37262
rect 80428 37198 80480 37204
rect 80334 36952 80390 36961
rect 80244 36916 80296 36922
rect 80334 36887 80336 36896
rect 80244 36858 80296 36864
rect 80388 36887 80390 36896
rect 80336 36858 80388 36864
rect 79968 36372 80020 36378
rect 79968 36314 80020 36320
rect 80152 36372 80204 36378
rect 80152 36314 80204 36320
rect 80060 36168 80112 36174
rect 80060 36110 80112 36116
rect 80072 35494 80100 36110
rect 80060 35488 80112 35494
rect 80060 35430 80112 35436
rect 80072 35154 80100 35430
rect 80256 35290 80284 36858
rect 80440 36174 80468 37198
rect 80808 37126 80836 37266
rect 80796 37120 80848 37126
rect 80796 37062 80848 37068
rect 80520 36780 80572 36786
rect 80520 36722 80572 36728
rect 80612 36780 80664 36786
rect 80612 36722 80664 36728
rect 80532 36378 80560 36722
rect 80520 36372 80572 36378
rect 80520 36314 80572 36320
rect 80624 36242 80652 36722
rect 80808 36718 80836 37062
rect 80796 36712 80848 36718
rect 80796 36654 80848 36660
rect 80612 36236 80664 36242
rect 80612 36178 80664 36184
rect 80428 36168 80480 36174
rect 80428 36110 80480 36116
rect 80900 35834 80928 39200
rect 81820 39114 81848 39200
rect 81912 39114 81940 39222
rect 81820 39086 81940 39114
rect 82084 39024 82136 39030
rect 82084 38966 82136 38972
rect 81348 37460 81400 37466
rect 81348 37402 81400 37408
rect 81360 37330 81388 37402
rect 81624 37392 81676 37398
rect 81624 37334 81676 37340
rect 81348 37324 81400 37330
rect 81348 37266 81400 37272
rect 81014 37020 81322 37029
rect 81014 37018 81020 37020
rect 81076 37018 81100 37020
rect 81156 37018 81180 37020
rect 81236 37018 81260 37020
rect 81316 37018 81322 37020
rect 81076 36966 81078 37018
rect 81258 36966 81260 37018
rect 81014 36964 81020 36966
rect 81076 36964 81100 36966
rect 81156 36964 81180 36966
rect 81236 36964 81260 36966
rect 81316 36964 81322 36966
rect 81014 36955 81322 36964
rect 81360 36242 81388 37266
rect 81440 37188 81492 37194
rect 81440 37130 81492 37136
rect 81348 36236 81400 36242
rect 81348 36178 81400 36184
rect 81014 35932 81322 35941
rect 81014 35930 81020 35932
rect 81076 35930 81100 35932
rect 81156 35930 81180 35932
rect 81236 35930 81260 35932
rect 81316 35930 81322 35932
rect 81076 35878 81078 35930
rect 81258 35878 81260 35930
rect 81014 35876 81020 35878
rect 81076 35876 81100 35878
rect 81156 35876 81180 35878
rect 81236 35876 81260 35878
rect 81316 35876 81322 35878
rect 81014 35867 81322 35876
rect 81360 35834 81388 36178
rect 80888 35828 80940 35834
rect 80888 35770 80940 35776
rect 81348 35828 81400 35834
rect 81348 35770 81400 35776
rect 80426 35728 80482 35737
rect 80426 35663 80428 35672
rect 80480 35663 80482 35672
rect 80428 35634 80480 35640
rect 81360 35630 81388 35770
rect 81348 35624 81400 35630
rect 81348 35566 81400 35572
rect 81360 35290 81388 35566
rect 81452 35562 81480 37130
rect 81636 36174 81664 37334
rect 81808 37120 81860 37126
rect 81808 37062 81860 37068
rect 81624 36168 81676 36174
rect 81624 36110 81676 36116
rect 81716 36168 81768 36174
rect 81716 36110 81768 36116
rect 81728 36038 81756 36110
rect 81716 36032 81768 36038
rect 81716 35974 81768 35980
rect 81440 35556 81492 35562
rect 81440 35498 81492 35504
rect 80244 35284 80296 35290
rect 80244 35226 80296 35232
rect 81348 35284 81400 35290
rect 81348 35226 81400 35232
rect 80060 35148 80112 35154
rect 80060 35090 80112 35096
rect 81014 34844 81322 34853
rect 81014 34842 81020 34844
rect 81076 34842 81100 34844
rect 81156 34842 81180 34844
rect 81236 34842 81260 34844
rect 81316 34842 81322 34844
rect 81076 34790 81078 34842
rect 81258 34790 81260 34842
rect 81014 34788 81020 34790
rect 81076 34788 81100 34790
rect 81156 34788 81180 34790
rect 81236 34788 81260 34790
rect 81316 34788 81322 34790
rect 81014 34779 81322 34788
rect 81014 33756 81322 33765
rect 81014 33754 81020 33756
rect 81076 33754 81100 33756
rect 81156 33754 81180 33756
rect 81236 33754 81260 33756
rect 81316 33754 81322 33756
rect 81076 33702 81078 33754
rect 81258 33702 81260 33754
rect 81014 33700 81020 33702
rect 81076 33700 81100 33702
rect 81156 33700 81180 33702
rect 81236 33700 81260 33702
rect 81316 33700 81322 33702
rect 81014 33691 81322 33700
rect 81014 32668 81322 32677
rect 81014 32666 81020 32668
rect 81076 32666 81100 32668
rect 81156 32666 81180 32668
rect 81236 32666 81260 32668
rect 81316 32666 81322 32668
rect 81076 32614 81078 32666
rect 81258 32614 81260 32666
rect 81014 32612 81020 32614
rect 81076 32612 81100 32614
rect 81156 32612 81180 32614
rect 81236 32612 81260 32614
rect 81316 32612 81322 32614
rect 81014 32603 81322 32612
rect 79796 31742 80100 31770
rect 80072 5914 80100 31742
rect 81014 31580 81322 31589
rect 81014 31578 81020 31580
rect 81076 31578 81100 31580
rect 81156 31578 81180 31580
rect 81236 31578 81260 31580
rect 81316 31578 81322 31580
rect 81076 31526 81078 31578
rect 81258 31526 81260 31578
rect 81014 31524 81020 31526
rect 81076 31524 81100 31526
rect 81156 31524 81180 31526
rect 81236 31524 81260 31526
rect 81316 31524 81322 31526
rect 81014 31515 81322 31524
rect 81014 30492 81322 30501
rect 81014 30490 81020 30492
rect 81076 30490 81100 30492
rect 81156 30490 81180 30492
rect 81236 30490 81260 30492
rect 81316 30490 81322 30492
rect 81076 30438 81078 30490
rect 81258 30438 81260 30490
rect 81014 30436 81020 30438
rect 81076 30436 81100 30438
rect 81156 30436 81180 30438
rect 81236 30436 81260 30438
rect 81316 30436 81322 30438
rect 81014 30427 81322 30436
rect 81014 29404 81322 29413
rect 81014 29402 81020 29404
rect 81076 29402 81100 29404
rect 81156 29402 81180 29404
rect 81236 29402 81260 29404
rect 81316 29402 81322 29404
rect 81076 29350 81078 29402
rect 81258 29350 81260 29402
rect 81014 29348 81020 29350
rect 81076 29348 81100 29350
rect 81156 29348 81180 29350
rect 81236 29348 81260 29350
rect 81316 29348 81322 29350
rect 81014 29339 81322 29348
rect 81014 28316 81322 28325
rect 81014 28314 81020 28316
rect 81076 28314 81100 28316
rect 81156 28314 81180 28316
rect 81236 28314 81260 28316
rect 81316 28314 81322 28316
rect 81076 28262 81078 28314
rect 81258 28262 81260 28314
rect 81014 28260 81020 28262
rect 81076 28260 81100 28262
rect 81156 28260 81180 28262
rect 81236 28260 81260 28262
rect 81316 28260 81322 28262
rect 81014 28251 81322 28260
rect 81014 27228 81322 27237
rect 81014 27226 81020 27228
rect 81076 27226 81100 27228
rect 81156 27226 81180 27228
rect 81236 27226 81260 27228
rect 81316 27226 81322 27228
rect 81076 27174 81078 27226
rect 81258 27174 81260 27226
rect 81014 27172 81020 27174
rect 81076 27172 81100 27174
rect 81156 27172 81180 27174
rect 81236 27172 81260 27174
rect 81316 27172 81322 27174
rect 81014 27163 81322 27172
rect 81820 26234 81848 37062
rect 82096 36786 82124 38966
rect 82084 36780 82136 36786
rect 82084 36722 82136 36728
rect 81900 36712 81952 36718
rect 81900 36654 81952 36660
rect 81912 35698 81940 36654
rect 82084 36576 82136 36582
rect 82188 36564 82216 39222
rect 82726 39200 82782 40000
rect 83646 39200 83702 40000
rect 83832 39228 83884 39234
rect 82740 37330 82768 39200
rect 83188 37868 83240 37874
rect 83188 37810 83240 37816
rect 83200 37398 83228 37810
rect 83188 37392 83240 37398
rect 82818 37360 82874 37369
rect 82728 37324 82780 37330
rect 83188 37334 83240 37340
rect 82818 37295 82874 37304
rect 83096 37324 83148 37330
rect 82728 37266 82780 37272
rect 82832 37262 82860 37295
rect 83096 37266 83148 37272
rect 82636 37256 82688 37262
rect 82636 37198 82688 37204
rect 82820 37256 82872 37262
rect 82820 37198 82872 37204
rect 82268 37188 82320 37194
rect 82268 37130 82320 37136
rect 82280 36786 82308 37130
rect 82452 37120 82504 37126
rect 82452 37062 82504 37068
rect 82648 37074 82676 37198
rect 83108 37126 83136 37266
rect 83096 37120 83148 37126
rect 82268 36780 82320 36786
rect 82268 36722 82320 36728
rect 82268 36576 82320 36582
rect 82188 36536 82268 36564
rect 82084 36518 82136 36524
rect 82268 36518 82320 36524
rect 81992 36032 82044 36038
rect 81992 35974 82044 35980
rect 81900 35692 81952 35698
rect 81900 35634 81952 35640
rect 82004 34134 82032 35974
rect 81900 34128 81952 34134
rect 81900 34070 81952 34076
rect 81992 34128 82044 34134
rect 81992 34070 82044 34076
rect 81912 33658 81940 34070
rect 81900 33652 81952 33658
rect 81900 33594 81952 33600
rect 82096 31754 82124 36518
rect 82360 36168 82412 36174
rect 82360 36110 82412 36116
rect 82372 35834 82400 36110
rect 82360 35828 82412 35834
rect 82360 35770 82412 35776
rect 82096 31726 82400 31754
rect 81728 26206 81848 26234
rect 81014 26140 81322 26149
rect 81014 26138 81020 26140
rect 81076 26138 81100 26140
rect 81156 26138 81180 26140
rect 81236 26138 81260 26140
rect 81316 26138 81322 26140
rect 81076 26086 81078 26138
rect 81258 26086 81260 26138
rect 81014 26084 81020 26086
rect 81076 26084 81100 26086
rect 81156 26084 81180 26086
rect 81236 26084 81260 26086
rect 81316 26084 81322 26086
rect 81014 26075 81322 26084
rect 81014 25052 81322 25061
rect 81014 25050 81020 25052
rect 81076 25050 81100 25052
rect 81156 25050 81180 25052
rect 81236 25050 81260 25052
rect 81316 25050 81322 25052
rect 81076 24998 81078 25050
rect 81258 24998 81260 25050
rect 81014 24996 81020 24998
rect 81076 24996 81100 24998
rect 81156 24996 81180 24998
rect 81236 24996 81260 24998
rect 81316 24996 81322 24998
rect 81014 24987 81322 24996
rect 81014 23964 81322 23973
rect 81014 23962 81020 23964
rect 81076 23962 81100 23964
rect 81156 23962 81180 23964
rect 81236 23962 81260 23964
rect 81316 23962 81322 23964
rect 81076 23910 81078 23962
rect 81258 23910 81260 23962
rect 81014 23908 81020 23910
rect 81076 23908 81100 23910
rect 81156 23908 81180 23910
rect 81236 23908 81260 23910
rect 81316 23908 81322 23910
rect 81014 23899 81322 23908
rect 81014 22876 81322 22885
rect 81014 22874 81020 22876
rect 81076 22874 81100 22876
rect 81156 22874 81180 22876
rect 81236 22874 81260 22876
rect 81316 22874 81322 22876
rect 81076 22822 81078 22874
rect 81258 22822 81260 22874
rect 81014 22820 81020 22822
rect 81076 22820 81100 22822
rect 81156 22820 81180 22822
rect 81236 22820 81260 22822
rect 81316 22820 81322 22822
rect 81014 22811 81322 22820
rect 81014 21788 81322 21797
rect 81014 21786 81020 21788
rect 81076 21786 81100 21788
rect 81156 21786 81180 21788
rect 81236 21786 81260 21788
rect 81316 21786 81322 21788
rect 81076 21734 81078 21786
rect 81258 21734 81260 21786
rect 81014 21732 81020 21734
rect 81076 21732 81100 21734
rect 81156 21732 81180 21734
rect 81236 21732 81260 21734
rect 81316 21732 81322 21734
rect 81014 21723 81322 21732
rect 81014 20700 81322 20709
rect 81014 20698 81020 20700
rect 81076 20698 81100 20700
rect 81156 20698 81180 20700
rect 81236 20698 81260 20700
rect 81316 20698 81322 20700
rect 81076 20646 81078 20698
rect 81258 20646 81260 20698
rect 81014 20644 81020 20646
rect 81076 20644 81100 20646
rect 81156 20644 81180 20646
rect 81236 20644 81260 20646
rect 81316 20644 81322 20646
rect 81014 20635 81322 20644
rect 81014 19612 81322 19621
rect 81014 19610 81020 19612
rect 81076 19610 81100 19612
rect 81156 19610 81180 19612
rect 81236 19610 81260 19612
rect 81316 19610 81322 19612
rect 81076 19558 81078 19610
rect 81258 19558 81260 19610
rect 81014 19556 81020 19558
rect 81076 19556 81100 19558
rect 81156 19556 81180 19558
rect 81236 19556 81260 19558
rect 81316 19556 81322 19558
rect 81014 19547 81322 19556
rect 81014 18524 81322 18533
rect 81014 18522 81020 18524
rect 81076 18522 81100 18524
rect 81156 18522 81180 18524
rect 81236 18522 81260 18524
rect 81316 18522 81322 18524
rect 81076 18470 81078 18522
rect 81258 18470 81260 18522
rect 81014 18468 81020 18470
rect 81076 18468 81100 18470
rect 81156 18468 81180 18470
rect 81236 18468 81260 18470
rect 81316 18468 81322 18470
rect 81014 18459 81322 18468
rect 81014 17436 81322 17445
rect 81014 17434 81020 17436
rect 81076 17434 81100 17436
rect 81156 17434 81180 17436
rect 81236 17434 81260 17436
rect 81316 17434 81322 17436
rect 81076 17382 81078 17434
rect 81258 17382 81260 17434
rect 81014 17380 81020 17382
rect 81076 17380 81100 17382
rect 81156 17380 81180 17382
rect 81236 17380 81260 17382
rect 81316 17380 81322 17382
rect 81014 17371 81322 17380
rect 81728 16574 81756 26206
rect 81728 16546 81848 16574
rect 81014 16348 81322 16357
rect 81014 16346 81020 16348
rect 81076 16346 81100 16348
rect 81156 16346 81180 16348
rect 81236 16346 81260 16348
rect 81316 16346 81322 16348
rect 81076 16294 81078 16346
rect 81258 16294 81260 16346
rect 81014 16292 81020 16294
rect 81076 16292 81100 16294
rect 81156 16292 81180 16294
rect 81236 16292 81260 16294
rect 81316 16292 81322 16294
rect 81014 16283 81322 16292
rect 81014 15260 81322 15269
rect 81014 15258 81020 15260
rect 81076 15258 81100 15260
rect 81156 15258 81180 15260
rect 81236 15258 81260 15260
rect 81316 15258 81322 15260
rect 81076 15206 81078 15258
rect 81258 15206 81260 15258
rect 81014 15204 81020 15206
rect 81076 15204 81100 15206
rect 81156 15204 81180 15206
rect 81236 15204 81260 15206
rect 81316 15204 81322 15206
rect 81014 15195 81322 15204
rect 81014 14172 81322 14181
rect 81014 14170 81020 14172
rect 81076 14170 81100 14172
rect 81156 14170 81180 14172
rect 81236 14170 81260 14172
rect 81316 14170 81322 14172
rect 81076 14118 81078 14170
rect 81258 14118 81260 14170
rect 81014 14116 81020 14118
rect 81076 14116 81100 14118
rect 81156 14116 81180 14118
rect 81236 14116 81260 14118
rect 81316 14116 81322 14118
rect 81014 14107 81322 14116
rect 81014 13084 81322 13093
rect 81014 13082 81020 13084
rect 81076 13082 81100 13084
rect 81156 13082 81180 13084
rect 81236 13082 81260 13084
rect 81316 13082 81322 13084
rect 81076 13030 81078 13082
rect 81258 13030 81260 13082
rect 81014 13028 81020 13030
rect 81076 13028 81100 13030
rect 81156 13028 81180 13030
rect 81236 13028 81260 13030
rect 81316 13028 81322 13030
rect 81014 13019 81322 13028
rect 81014 11996 81322 12005
rect 81014 11994 81020 11996
rect 81076 11994 81100 11996
rect 81156 11994 81180 11996
rect 81236 11994 81260 11996
rect 81316 11994 81322 11996
rect 81076 11942 81078 11994
rect 81258 11942 81260 11994
rect 81014 11940 81020 11942
rect 81076 11940 81100 11942
rect 81156 11940 81180 11942
rect 81236 11940 81260 11942
rect 81316 11940 81322 11942
rect 81014 11931 81322 11940
rect 81014 10908 81322 10917
rect 81014 10906 81020 10908
rect 81076 10906 81100 10908
rect 81156 10906 81180 10908
rect 81236 10906 81260 10908
rect 81316 10906 81322 10908
rect 81076 10854 81078 10906
rect 81258 10854 81260 10906
rect 81014 10852 81020 10854
rect 81076 10852 81100 10854
rect 81156 10852 81180 10854
rect 81236 10852 81260 10854
rect 81316 10852 81322 10854
rect 81014 10843 81322 10852
rect 81014 9820 81322 9829
rect 81014 9818 81020 9820
rect 81076 9818 81100 9820
rect 81156 9818 81180 9820
rect 81236 9818 81260 9820
rect 81316 9818 81322 9820
rect 81076 9766 81078 9818
rect 81258 9766 81260 9818
rect 81014 9764 81020 9766
rect 81076 9764 81100 9766
rect 81156 9764 81180 9766
rect 81236 9764 81260 9766
rect 81316 9764 81322 9766
rect 81014 9755 81322 9764
rect 81014 8732 81322 8741
rect 81014 8730 81020 8732
rect 81076 8730 81100 8732
rect 81156 8730 81180 8732
rect 81236 8730 81260 8732
rect 81316 8730 81322 8732
rect 81076 8678 81078 8730
rect 81258 8678 81260 8730
rect 81014 8676 81020 8678
rect 81076 8676 81100 8678
rect 81156 8676 81180 8678
rect 81236 8676 81260 8678
rect 81316 8676 81322 8678
rect 81014 8667 81322 8676
rect 81014 7644 81322 7653
rect 81014 7642 81020 7644
rect 81076 7642 81100 7644
rect 81156 7642 81180 7644
rect 81236 7642 81260 7644
rect 81316 7642 81322 7644
rect 81076 7590 81078 7642
rect 81258 7590 81260 7642
rect 81014 7588 81020 7590
rect 81076 7588 81100 7590
rect 81156 7588 81180 7590
rect 81236 7588 81260 7590
rect 81316 7588 81322 7590
rect 81014 7579 81322 7588
rect 81014 6556 81322 6565
rect 81014 6554 81020 6556
rect 81076 6554 81100 6556
rect 81156 6554 81180 6556
rect 81236 6554 81260 6556
rect 81316 6554 81322 6556
rect 81076 6502 81078 6554
rect 81258 6502 81260 6554
rect 81014 6500 81020 6502
rect 81076 6500 81100 6502
rect 81156 6500 81180 6502
rect 81236 6500 81260 6502
rect 81316 6500 81322 6502
rect 81014 6491 81322 6500
rect 80060 5908 80112 5914
rect 80060 5850 80112 5856
rect 79048 5704 79100 5710
rect 79048 5646 79100 5652
rect 78496 5568 78548 5574
rect 78496 5510 78548 5516
rect 79140 5568 79192 5574
rect 79140 5510 79192 5516
rect 79152 5098 79180 5510
rect 79140 5092 79192 5098
rect 79140 5034 79192 5040
rect 78220 4820 78272 4826
rect 78220 4762 78272 4768
rect 77668 4480 77720 4486
rect 77668 4422 77720 4428
rect 77680 3398 77708 4422
rect 78232 3534 78260 4762
rect 78680 4684 78732 4690
rect 78680 4626 78732 4632
rect 78692 4486 78720 4626
rect 78680 4480 78732 4486
rect 78680 4422 78732 4428
rect 78772 4480 78824 4486
rect 78772 4422 78824 4428
rect 78692 4010 78720 4422
rect 78784 4146 78812 4422
rect 78772 4140 78824 4146
rect 78772 4082 78824 4088
rect 79152 4078 79180 5034
rect 79416 5024 79468 5030
rect 79416 4966 79468 4972
rect 79508 5024 79560 5030
rect 79508 4966 79560 4972
rect 79140 4072 79192 4078
rect 79140 4014 79192 4020
rect 78680 4004 78732 4010
rect 78680 3946 78732 3952
rect 78772 3936 78824 3942
rect 78772 3878 78824 3884
rect 78784 3602 78812 3878
rect 78772 3596 78824 3602
rect 78772 3538 78824 3544
rect 78220 3528 78272 3534
rect 78220 3470 78272 3476
rect 77668 3392 77720 3398
rect 77668 3334 77720 3340
rect 78128 3392 78180 3398
rect 78128 3334 78180 3340
rect 77208 3188 77260 3194
rect 77208 3130 77260 3136
rect 77024 3052 77076 3058
rect 77024 2994 77076 3000
rect 76840 2916 76892 2922
rect 76840 2858 76892 2864
rect 76472 2848 76524 2854
rect 76472 2790 76524 2796
rect 76564 2848 76616 2854
rect 76564 2790 76616 2796
rect 76484 2514 76512 2790
rect 76472 2508 76524 2514
rect 76472 2450 76524 2456
rect 76852 2378 76880 2858
rect 76380 2372 76432 2378
rect 76380 2314 76432 2320
rect 76840 2372 76892 2378
rect 76840 2314 76892 2320
rect 77036 800 77064 2994
rect 78140 2378 78168 3334
rect 79152 2990 79180 4014
rect 79428 3466 79456 4966
rect 79520 4214 79548 4966
rect 79784 4684 79836 4690
rect 79784 4626 79836 4632
rect 79508 4208 79560 4214
rect 79508 4150 79560 4156
rect 79796 4078 79824 4626
rect 80072 4622 80100 5850
rect 80152 5568 80204 5574
rect 80152 5510 80204 5516
rect 80060 4616 80112 4622
rect 80060 4558 80112 4564
rect 80164 4486 80192 5510
rect 81014 5468 81322 5477
rect 81014 5466 81020 5468
rect 81076 5466 81100 5468
rect 81156 5466 81180 5468
rect 81236 5466 81260 5468
rect 81316 5466 81322 5468
rect 81076 5414 81078 5466
rect 81258 5414 81260 5466
rect 81014 5412 81020 5414
rect 81076 5412 81100 5414
rect 81156 5412 81180 5414
rect 81236 5412 81260 5414
rect 81316 5412 81322 5414
rect 81014 5403 81322 5412
rect 81716 5160 81768 5166
rect 81716 5102 81768 5108
rect 81440 5092 81492 5098
rect 81440 5034 81492 5040
rect 80244 5024 80296 5030
rect 80244 4966 80296 4972
rect 80796 5024 80848 5030
rect 80796 4966 80848 4972
rect 80152 4480 80204 4486
rect 80152 4422 80204 4428
rect 79784 4072 79836 4078
rect 79784 4014 79836 4020
rect 80164 3602 80192 4422
rect 80152 3596 80204 3602
rect 80152 3538 80204 3544
rect 79416 3460 79468 3466
rect 79416 3402 79468 3408
rect 79784 3188 79836 3194
rect 79784 3130 79836 3136
rect 78680 2984 78732 2990
rect 78680 2926 78732 2932
rect 79140 2984 79192 2990
rect 79140 2926 79192 2932
rect 78692 2514 78720 2926
rect 78680 2508 78732 2514
rect 78680 2450 78732 2456
rect 78128 2372 78180 2378
rect 78128 2314 78180 2320
rect 78140 1698 78168 2314
rect 78128 1692 78180 1698
rect 78128 1634 78180 1640
rect 79796 800 79824 3130
rect 80256 2990 80284 4966
rect 80428 4616 80480 4622
rect 80428 4558 80480 4564
rect 80336 4548 80388 4554
rect 80336 4490 80388 4496
rect 80244 2984 80296 2990
rect 80244 2926 80296 2932
rect 80348 2774 80376 4490
rect 80440 3738 80468 4558
rect 80428 3732 80480 3738
rect 80428 3674 80480 3680
rect 80256 2746 80376 2774
rect 80256 2514 80284 2746
rect 80244 2508 80296 2514
rect 80244 2450 80296 2456
rect 80808 2446 80836 4966
rect 81348 4480 81400 4486
rect 81348 4422 81400 4428
rect 81014 4380 81322 4389
rect 81014 4378 81020 4380
rect 81076 4378 81100 4380
rect 81156 4378 81180 4380
rect 81236 4378 81260 4380
rect 81316 4378 81322 4380
rect 81076 4326 81078 4378
rect 81258 4326 81260 4378
rect 81014 4324 81020 4326
rect 81076 4324 81100 4326
rect 81156 4324 81180 4326
rect 81236 4324 81260 4326
rect 81316 4324 81322 4326
rect 81014 4315 81322 4324
rect 81360 4214 81388 4422
rect 81452 4282 81480 5034
rect 81532 4752 81584 4758
rect 81532 4694 81584 4700
rect 81440 4276 81492 4282
rect 81440 4218 81492 4224
rect 81348 4208 81400 4214
rect 81348 4150 81400 4156
rect 81440 3936 81492 3942
rect 81440 3878 81492 3884
rect 81346 3632 81402 3641
rect 81346 3567 81348 3576
rect 81400 3567 81402 3576
rect 81348 3538 81400 3544
rect 81014 3292 81322 3301
rect 81014 3290 81020 3292
rect 81076 3290 81100 3292
rect 81156 3290 81180 3292
rect 81236 3290 81260 3292
rect 81316 3290 81322 3292
rect 81076 3238 81078 3290
rect 81258 3238 81260 3290
rect 81014 3236 81020 3238
rect 81076 3236 81100 3238
rect 81156 3236 81180 3238
rect 81236 3236 81260 3238
rect 81316 3236 81322 3238
rect 81014 3227 81322 3236
rect 81348 2644 81400 2650
rect 81348 2586 81400 2592
rect 80796 2440 80848 2446
rect 80796 2382 80848 2388
rect 81360 2310 81388 2586
rect 81348 2304 81400 2310
rect 81348 2246 81400 2252
rect 81014 2204 81322 2213
rect 81014 2202 81020 2204
rect 81076 2202 81100 2204
rect 81156 2202 81180 2204
rect 81236 2202 81260 2204
rect 81316 2202 81322 2204
rect 81076 2150 81078 2202
rect 81258 2150 81260 2202
rect 81014 2148 81020 2150
rect 81076 2148 81100 2150
rect 81156 2148 81180 2150
rect 81236 2148 81260 2150
rect 81316 2148 81322 2150
rect 81014 2139 81322 2148
rect 81164 1896 81216 1902
rect 81164 1838 81216 1844
rect 81176 800 81204 1838
rect 81452 1494 81480 3878
rect 81544 2394 81572 4694
rect 81728 3194 81756 5102
rect 81820 3466 81848 16546
rect 81992 5024 82044 5030
rect 81992 4966 82044 4972
rect 82004 4690 82032 4966
rect 81992 4684 82044 4690
rect 81992 4626 82044 4632
rect 82084 4616 82136 4622
rect 82084 4558 82136 4564
rect 81992 4072 82044 4078
rect 81992 4014 82044 4020
rect 82004 3602 82032 4014
rect 82096 3738 82124 4558
rect 82084 3732 82136 3738
rect 82084 3674 82136 3680
rect 81992 3596 82044 3602
rect 81992 3538 82044 3544
rect 81808 3460 81860 3466
rect 81808 3402 81860 3408
rect 81716 3188 81768 3194
rect 81716 3130 81768 3136
rect 82004 2990 82032 3538
rect 82372 3466 82400 31726
rect 82464 6866 82492 37062
rect 82648 37046 82860 37074
rect 83096 37062 83148 37068
rect 82832 36242 82860 37046
rect 83188 36780 83240 36786
rect 83188 36722 83240 36728
rect 82820 36236 82872 36242
rect 82820 36178 82872 36184
rect 83096 36032 83148 36038
rect 83096 35974 83148 35980
rect 83108 35698 83136 35974
rect 83096 35692 83148 35698
rect 83096 35634 83148 35640
rect 82912 35488 82964 35494
rect 82912 35430 82964 35436
rect 82924 26234 82952 35430
rect 83108 34406 83136 35634
rect 83096 34400 83148 34406
rect 83096 34342 83148 34348
rect 83200 33522 83228 36722
rect 83660 36582 83688 39200
rect 84566 39200 84622 40000
rect 84936 39296 84988 39302
rect 84936 39238 84988 39244
rect 83832 39170 83884 39176
rect 83844 36786 83872 39170
rect 84200 37324 84252 37330
rect 84200 37266 84252 37272
rect 83924 37188 83976 37194
rect 83924 37130 83976 37136
rect 83740 36780 83792 36786
rect 83740 36722 83792 36728
rect 83832 36780 83884 36786
rect 83832 36722 83884 36728
rect 83648 36576 83700 36582
rect 83648 36518 83700 36524
rect 83648 36236 83700 36242
rect 83648 36178 83700 36184
rect 83660 36038 83688 36178
rect 83752 36038 83780 36722
rect 83648 36032 83700 36038
rect 83648 35974 83700 35980
rect 83740 36032 83792 36038
rect 83740 35974 83792 35980
rect 83660 35630 83688 35974
rect 83844 35834 83872 36722
rect 83832 35828 83884 35834
rect 83832 35770 83884 35776
rect 83648 35624 83700 35630
rect 83648 35566 83700 35572
rect 83936 35494 83964 37130
rect 84212 36038 84240 37266
rect 84580 37194 84608 39200
rect 84844 37256 84896 37262
rect 84844 37198 84896 37204
rect 84568 37188 84620 37194
rect 84568 37130 84620 37136
rect 84660 37120 84712 37126
rect 84660 37062 84712 37068
rect 84672 36417 84700 37062
rect 84750 36816 84806 36825
rect 84750 36751 84806 36760
rect 84764 36553 84792 36751
rect 84856 36718 84884 37198
rect 84948 36786 84976 39238
rect 85486 39200 85542 40000
rect 86406 39200 86462 40000
rect 86512 39222 86908 39250
rect 85304 39160 85356 39166
rect 85304 39102 85356 39108
rect 85316 37262 85344 39102
rect 85304 37256 85356 37262
rect 85304 37198 85356 37204
rect 84936 36780 84988 36786
rect 84936 36722 84988 36728
rect 84844 36712 84896 36718
rect 84844 36654 84896 36660
rect 84750 36544 84806 36553
rect 84750 36479 84806 36488
rect 84658 36408 84714 36417
rect 84658 36343 84714 36352
rect 84200 36032 84252 36038
rect 84200 35974 84252 35980
rect 84752 36032 84804 36038
rect 84752 35974 84804 35980
rect 83924 35488 83976 35494
rect 83924 35430 83976 35436
rect 84764 35290 84792 35974
rect 85316 35834 85344 37198
rect 85500 37074 85528 39200
rect 86420 39114 86448 39200
rect 86512 39114 86540 39222
rect 86420 39086 86540 39114
rect 85762 37632 85818 37641
rect 85762 37567 85818 37576
rect 85580 37120 85632 37126
rect 85500 37068 85580 37074
rect 85500 37062 85632 37068
rect 85500 37046 85620 37062
rect 85488 36780 85540 36786
rect 85488 36722 85540 36728
rect 85500 36038 85528 36722
rect 85776 36718 85804 37567
rect 86776 37256 86828 37262
rect 86880 37244 86908 39222
rect 87326 39200 87382 40000
rect 88246 39200 88302 40000
rect 89166 39200 89222 40000
rect 90086 39200 90142 40000
rect 91006 39200 91062 40000
rect 91926 39200 91982 40000
rect 92846 39200 92902 40000
rect 93766 39200 93822 40000
rect 94686 39200 94742 40000
rect 94792 39222 95188 39250
rect 86960 37256 87012 37262
rect 86880 37216 86960 37244
rect 86776 37198 86828 37204
rect 86960 37198 87012 37204
rect 85764 36712 85816 36718
rect 85764 36654 85816 36660
rect 86408 36576 86460 36582
rect 86788 36564 86816 37198
rect 87340 37126 87368 39200
rect 87512 37256 87564 37262
rect 87512 37198 87564 37204
rect 88064 37256 88116 37262
rect 88064 37198 88116 37204
rect 87236 37120 87288 37126
rect 87236 37062 87288 37068
rect 87328 37120 87380 37126
rect 87328 37062 87380 37068
rect 87248 36854 87276 37062
rect 87524 36854 87552 37198
rect 87236 36848 87288 36854
rect 87236 36790 87288 36796
rect 87512 36848 87564 36854
rect 87512 36790 87564 36796
rect 87604 36848 87656 36854
rect 87604 36790 87656 36796
rect 86868 36576 86920 36582
rect 86788 36536 86868 36564
rect 86408 36518 86460 36524
rect 86868 36518 86920 36524
rect 86420 36310 86448 36518
rect 86408 36304 86460 36310
rect 86408 36246 86460 36252
rect 85488 36032 85540 36038
rect 85488 35974 85540 35980
rect 85304 35828 85356 35834
rect 85304 35770 85356 35776
rect 84752 35284 84804 35290
rect 84752 35226 84804 35232
rect 83832 34128 83884 34134
rect 83832 34070 83884 34076
rect 83188 33516 83240 33522
rect 83188 33458 83240 33464
rect 82924 26206 83228 26234
rect 82452 6860 82504 6866
rect 82452 6802 82504 6808
rect 83096 6860 83148 6866
rect 83096 6802 83148 6808
rect 83004 5024 83056 5030
rect 83004 4966 83056 4972
rect 82820 4480 82872 4486
rect 82820 4422 82872 4428
rect 82728 4276 82780 4282
rect 82728 4218 82780 4224
rect 82740 4010 82768 4218
rect 82728 4004 82780 4010
rect 82728 3946 82780 3952
rect 82728 3732 82780 3738
rect 82728 3674 82780 3680
rect 82360 3460 82412 3466
rect 82360 3402 82412 3408
rect 82372 3194 82400 3402
rect 82740 3398 82768 3674
rect 82832 3534 82860 4422
rect 83016 4078 83044 4966
rect 83108 4826 83136 6802
rect 83096 4820 83148 4826
rect 83096 4762 83148 4768
rect 83108 4146 83136 4762
rect 83096 4140 83148 4146
rect 83096 4082 83148 4088
rect 83004 4072 83056 4078
rect 83004 4014 83056 4020
rect 82820 3528 82872 3534
rect 82872 3476 83044 3482
rect 82820 3470 83044 3476
rect 82832 3454 83044 3470
rect 82728 3392 82780 3398
rect 82728 3334 82780 3340
rect 82360 3188 82412 3194
rect 82360 3130 82412 3136
rect 82820 3120 82872 3126
rect 82820 3062 82872 3068
rect 81992 2984 82044 2990
rect 81992 2926 82044 2932
rect 82832 2446 82860 3062
rect 82912 2576 82964 2582
rect 82912 2518 82964 2524
rect 82820 2440 82872 2446
rect 81544 2378 81664 2394
rect 82820 2382 82872 2388
rect 81544 2372 81676 2378
rect 81544 2366 81624 2372
rect 81624 2314 81676 2320
rect 82820 2304 82872 2310
rect 82924 2258 82952 2518
rect 83016 2310 83044 3454
rect 83200 3194 83228 26206
rect 83372 5092 83424 5098
rect 83372 5034 83424 5040
rect 83278 3632 83334 3641
rect 83278 3567 83280 3576
rect 83332 3567 83334 3576
rect 83280 3538 83332 3544
rect 83384 3398 83412 5034
rect 83844 4146 83872 34070
rect 84200 4548 84252 4554
rect 84200 4490 84252 4496
rect 83832 4140 83884 4146
rect 83832 4082 83884 4088
rect 83648 4072 83700 4078
rect 83648 4014 83700 4020
rect 83464 3936 83516 3942
rect 83464 3878 83516 3884
rect 83372 3392 83424 3398
rect 83372 3334 83424 3340
rect 83384 3194 83412 3334
rect 83188 3188 83240 3194
rect 83188 3130 83240 3136
rect 83372 3188 83424 3194
rect 83372 3130 83424 3136
rect 83280 3052 83332 3058
rect 83476 3040 83504 3878
rect 83660 3398 83688 4014
rect 83844 3534 83872 4082
rect 83832 3528 83884 3534
rect 83832 3470 83884 3476
rect 83648 3392 83700 3398
rect 83648 3334 83700 3340
rect 83332 3012 83504 3040
rect 83280 2994 83332 3000
rect 83188 2848 83240 2854
rect 83108 2796 83188 2802
rect 83108 2790 83240 2796
rect 83108 2774 83228 2790
rect 83108 2378 83136 2774
rect 83096 2372 83148 2378
rect 83096 2314 83148 2320
rect 82872 2252 82952 2258
rect 82820 2246 82952 2252
rect 83004 2304 83056 2310
rect 83004 2246 83056 2252
rect 82832 2230 82952 2246
rect 83016 1562 83044 2246
rect 83292 1902 83320 2994
rect 83660 2990 83688 3334
rect 84108 3188 84160 3194
rect 84108 3130 84160 3136
rect 83648 2984 83700 2990
rect 83648 2926 83700 2932
rect 84120 2582 84148 3130
rect 84212 3058 84240 4490
rect 84844 3732 84896 3738
rect 84844 3674 84896 3680
rect 84200 3052 84252 3058
rect 84200 2994 84252 3000
rect 84856 2922 84884 3674
rect 85396 3392 85448 3398
rect 85396 3334 85448 3340
rect 85408 3058 85436 3334
rect 84936 3052 84988 3058
rect 84936 2994 84988 3000
rect 85396 3052 85448 3058
rect 85396 2994 85448 3000
rect 84844 2916 84896 2922
rect 84844 2858 84896 2864
rect 84108 2576 84160 2582
rect 84108 2518 84160 2524
rect 84200 2508 84252 2514
rect 84200 2450 84252 2456
rect 84212 2310 84240 2450
rect 84948 2446 84976 2994
rect 85500 2650 85528 35974
rect 86880 33590 86908 36518
rect 87616 36174 87644 36790
rect 88076 36582 88104 37198
rect 88260 37074 88288 39200
rect 88340 37120 88392 37126
rect 88260 37068 88340 37074
rect 88260 37062 88392 37068
rect 88260 37046 88380 37062
rect 89076 36780 89128 36786
rect 89076 36722 89128 36728
rect 88064 36576 88116 36582
rect 88064 36518 88116 36524
rect 87604 36168 87656 36174
rect 87604 36110 87656 36116
rect 86868 33584 86920 33590
rect 86868 33526 86920 33532
rect 88076 32978 88104 36518
rect 89088 36038 89116 36722
rect 89180 36582 89208 39200
rect 89812 38956 89864 38962
rect 89812 38898 89864 38904
rect 89824 37466 89852 38898
rect 89720 37460 89772 37466
rect 89720 37402 89772 37408
rect 89812 37460 89864 37466
rect 89812 37402 89864 37408
rect 89732 37330 89760 37402
rect 89720 37324 89772 37330
rect 89720 37266 89772 37272
rect 90100 37262 90128 39200
rect 89628 37256 89680 37262
rect 89628 37198 89680 37204
rect 90088 37256 90140 37262
rect 90088 37198 90140 37204
rect 90732 37256 90784 37262
rect 90732 37198 90784 37204
rect 89260 37120 89312 37126
rect 89260 37062 89312 37068
rect 89168 36576 89220 36582
rect 89168 36518 89220 36524
rect 89272 36378 89300 37062
rect 89260 36372 89312 36378
rect 89260 36314 89312 36320
rect 89640 36038 89668 37198
rect 90364 37188 90416 37194
rect 90364 37130 90416 37136
rect 90376 36786 90404 37130
rect 90364 36780 90416 36786
rect 90364 36722 90416 36728
rect 90376 36038 90404 36722
rect 90456 36576 90508 36582
rect 90456 36518 90508 36524
rect 89076 36032 89128 36038
rect 89076 35974 89128 35980
rect 89628 36032 89680 36038
rect 89628 35974 89680 35980
rect 89720 36032 89772 36038
rect 89720 35974 89772 35980
rect 90364 36032 90416 36038
rect 90364 35974 90416 35980
rect 89088 33969 89116 35974
rect 89074 33960 89130 33969
rect 89074 33895 89130 33904
rect 89640 33658 89668 35974
rect 89628 33652 89680 33658
rect 89628 33594 89680 33600
rect 88064 32972 88116 32978
rect 88064 32914 88116 32920
rect 85672 2848 85724 2854
rect 85672 2790 85724 2796
rect 85488 2644 85540 2650
rect 85488 2586 85540 2592
rect 84936 2440 84988 2446
rect 84936 2382 84988 2388
rect 85304 2372 85356 2378
rect 85304 2314 85356 2320
rect 83924 2304 83976 2310
rect 83924 2246 83976 2252
rect 84200 2304 84252 2310
rect 84200 2246 84252 2252
rect 83280 1896 83332 1902
rect 83280 1838 83332 1844
rect 83004 1556 83056 1562
rect 83004 1498 83056 1504
rect 81440 1488 81492 1494
rect 81440 1430 81492 1436
rect 83936 800 83964 2246
rect 85316 800 85344 2314
rect 85684 2310 85712 2790
rect 89732 2650 89760 35974
rect 90468 35562 90496 36518
rect 90744 36378 90772 37198
rect 91020 37074 91048 39200
rect 91560 37256 91612 37262
rect 91560 37198 91612 37204
rect 91100 37120 91152 37126
rect 91020 37068 91100 37074
rect 91020 37062 91152 37068
rect 91020 37046 91140 37062
rect 91572 36582 91600 37198
rect 91940 37126 91968 39200
rect 92112 37256 92164 37262
rect 92112 37198 92164 37204
rect 91928 37120 91980 37126
rect 91928 37062 91980 37068
rect 92124 36582 92152 37198
rect 92860 37126 92888 39200
rect 93032 38888 93084 38894
rect 93032 38830 93084 38836
rect 92940 37256 92992 37262
rect 92940 37198 92992 37204
rect 92848 37120 92900 37126
rect 92848 37062 92900 37068
rect 92952 36938 92980 37198
rect 92860 36910 92980 36938
rect 91560 36576 91612 36582
rect 91560 36518 91612 36524
rect 92112 36576 92164 36582
rect 92112 36518 92164 36524
rect 90732 36372 90784 36378
rect 90732 36314 90784 36320
rect 90456 35556 90508 35562
rect 90456 35498 90508 35504
rect 91572 32842 91600 36518
rect 92124 34105 92152 36518
rect 92388 36100 92440 36106
rect 92388 36042 92440 36048
rect 92400 35018 92428 36042
rect 92860 36038 92888 36910
rect 93044 36786 93072 38830
rect 93780 37244 93808 39200
rect 94700 39114 94728 39200
rect 94792 39114 94820 39222
rect 94700 39086 94820 39114
rect 95056 38888 95108 38894
rect 95056 38830 95108 38836
rect 94228 38820 94280 38826
rect 94228 38762 94280 38768
rect 94240 37466 94268 38762
rect 95068 37466 95096 38830
rect 94228 37460 94280 37466
rect 94228 37402 94280 37408
rect 95056 37460 95108 37466
rect 95056 37402 95108 37408
rect 93860 37256 93912 37262
rect 93780 37216 93860 37244
rect 93860 37198 93912 37204
rect 93032 36780 93084 36786
rect 93032 36722 93084 36728
rect 93872 36378 93900 37198
rect 94320 37120 94372 37126
rect 94320 37062 94372 37068
rect 95160 37074 95188 39222
rect 95606 39200 95662 40000
rect 96526 39200 96582 40000
rect 97446 39200 97502 40000
rect 97552 39222 97948 39250
rect 95240 37120 95292 37126
rect 95160 37068 95240 37074
rect 95160 37062 95292 37068
rect 94332 36786 94360 37062
rect 95160 37046 95280 37062
rect 94320 36780 94372 36786
rect 94320 36722 94372 36728
rect 95240 36780 95292 36786
rect 95240 36722 95292 36728
rect 94332 36582 94360 36722
rect 94320 36576 94372 36582
rect 94320 36518 94372 36524
rect 95056 36576 95108 36582
rect 95056 36518 95108 36524
rect 93860 36372 93912 36378
rect 93860 36314 93912 36320
rect 94332 36038 94360 36518
rect 95068 36174 95096 36518
rect 95056 36168 95108 36174
rect 95056 36110 95108 36116
rect 95252 36106 95280 36722
rect 95620 36582 95648 39200
rect 96540 37754 96568 39200
rect 97460 39114 97488 39200
rect 97552 39114 97580 39222
rect 97460 39086 97580 39114
rect 97540 38004 97592 38010
rect 97540 37946 97592 37952
rect 96540 37726 96752 37754
rect 96374 37564 96682 37573
rect 96374 37562 96380 37564
rect 96436 37562 96460 37564
rect 96516 37562 96540 37564
rect 96596 37562 96620 37564
rect 96676 37562 96682 37564
rect 96436 37510 96438 37562
rect 96618 37510 96620 37562
rect 96374 37508 96380 37510
rect 96436 37508 96460 37510
rect 96516 37508 96540 37510
rect 96596 37508 96620 37510
rect 96676 37508 96682 37510
rect 96374 37499 96682 37508
rect 96724 37262 96752 37726
rect 97552 37466 97580 37946
rect 97540 37460 97592 37466
rect 97540 37402 97592 37408
rect 96160 37256 96212 37262
rect 96160 37198 96212 37204
rect 96712 37256 96764 37262
rect 96712 37198 96764 37204
rect 95884 36780 95936 36786
rect 95884 36722 95936 36728
rect 95608 36576 95660 36582
rect 95608 36518 95660 36524
rect 95240 36100 95292 36106
rect 95240 36042 95292 36048
rect 95896 36038 95924 36722
rect 96172 36582 96200 37198
rect 96724 36854 96752 37198
rect 97816 37188 97868 37194
rect 97816 37130 97868 37136
rect 96804 37120 96856 37126
rect 96802 37088 96804 37097
rect 96856 37088 96858 37097
rect 96802 37023 96858 37032
rect 96712 36848 96764 36854
rect 96712 36790 96764 36796
rect 96160 36576 96212 36582
rect 96160 36518 96212 36524
rect 92848 36032 92900 36038
rect 92848 35974 92900 35980
rect 94320 36032 94372 36038
rect 94320 35974 94372 35980
rect 95884 36032 95936 36038
rect 95884 35974 95936 35980
rect 92388 35012 92440 35018
rect 92388 34954 92440 34960
rect 92860 34513 92888 35974
rect 92846 34504 92902 34513
rect 92846 34439 92902 34448
rect 92110 34096 92166 34105
rect 92110 34031 92166 34040
rect 91560 32836 91612 32842
rect 91560 32778 91612 32784
rect 94332 2650 94360 35974
rect 95896 33561 95924 35974
rect 95882 33552 95938 33561
rect 95882 33487 95938 33496
rect 96172 31754 96200 36518
rect 96374 36476 96682 36485
rect 96374 36474 96380 36476
rect 96436 36474 96460 36476
rect 96516 36474 96540 36476
rect 96596 36474 96620 36476
rect 96676 36474 96682 36476
rect 96436 36422 96438 36474
rect 96618 36422 96620 36474
rect 96374 36420 96380 36422
rect 96436 36420 96460 36422
rect 96516 36420 96540 36422
rect 96596 36420 96620 36422
rect 96676 36420 96682 36422
rect 96374 36411 96682 36420
rect 97828 36038 97856 37130
rect 97920 37074 97948 39222
rect 98366 39200 98422 40000
rect 98472 39222 98684 39250
rect 98380 39114 98408 39200
rect 98472 39114 98500 39222
rect 98380 39086 98500 39114
rect 98460 37256 98512 37262
rect 98460 37198 98512 37204
rect 98000 37120 98052 37126
rect 97920 37068 98000 37074
rect 97920 37062 98052 37068
rect 97920 37046 98040 37062
rect 98000 36780 98052 36786
rect 98000 36722 98052 36728
rect 98012 36582 98040 36722
rect 98000 36576 98052 36582
rect 98000 36518 98052 36524
rect 97816 36032 97868 36038
rect 97816 35974 97868 35980
rect 96374 35388 96682 35397
rect 96374 35386 96380 35388
rect 96436 35386 96460 35388
rect 96516 35386 96540 35388
rect 96596 35386 96620 35388
rect 96676 35386 96682 35388
rect 96436 35334 96438 35386
rect 96618 35334 96620 35386
rect 96374 35332 96380 35334
rect 96436 35332 96460 35334
rect 96516 35332 96540 35334
rect 96596 35332 96620 35334
rect 96676 35332 96682 35334
rect 96374 35323 96682 35332
rect 96374 34300 96682 34309
rect 96374 34298 96380 34300
rect 96436 34298 96460 34300
rect 96516 34298 96540 34300
rect 96596 34298 96620 34300
rect 96676 34298 96682 34300
rect 96436 34246 96438 34298
rect 96618 34246 96620 34298
rect 96374 34244 96380 34246
rect 96436 34244 96460 34246
rect 96516 34244 96540 34246
rect 96596 34244 96620 34246
rect 96676 34244 96682 34246
rect 96374 34235 96682 34244
rect 96374 33212 96682 33221
rect 96374 33210 96380 33212
rect 96436 33210 96460 33212
rect 96516 33210 96540 33212
rect 96596 33210 96620 33212
rect 96676 33210 96682 33212
rect 96436 33158 96438 33210
rect 96618 33158 96620 33210
rect 96374 33156 96380 33158
rect 96436 33156 96460 33158
rect 96516 33156 96540 33158
rect 96596 33156 96620 33158
rect 96676 33156 96682 33158
rect 96374 33147 96682 33156
rect 96374 32124 96682 32133
rect 96374 32122 96380 32124
rect 96436 32122 96460 32124
rect 96516 32122 96540 32124
rect 96596 32122 96620 32124
rect 96676 32122 96682 32124
rect 96436 32070 96438 32122
rect 96618 32070 96620 32122
rect 96374 32068 96380 32070
rect 96436 32068 96460 32070
rect 96516 32068 96540 32070
rect 96596 32068 96620 32070
rect 96676 32068 96682 32070
rect 96374 32059 96682 32068
rect 96160 31748 96212 31754
rect 96160 31690 96212 31696
rect 96374 31036 96682 31045
rect 96374 31034 96380 31036
rect 96436 31034 96460 31036
rect 96516 31034 96540 31036
rect 96596 31034 96620 31036
rect 96676 31034 96682 31036
rect 96436 30982 96438 31034
rect 96618 30982 96620 31034
rect 96374 30980 96380 30982
rect 96436 30980 96460 30982
rect 96516 30980 96540 30982
rect 96596 30980 96620 30982
rect 96676 30980 96682 30982
rect 96374 30971 96682 30980
rect 96374 29948 96682 29957
rect 96374 29946 96380 29948
rect 96436 29946 96460 29948
rect 96516 29946 96540 29948
rect 96596 29946 96620 29948
rect 96676 29946 96682 29948
rect 96436 29894 96438 29946
rect 96618 29894 96620 29946
rect 96374 29892 96380 29894
rect 96436 29892 96460 29894
rect 96516 29892 96540 29894
rect 96596 29892 96620 29894
rect 96676 29892 96682 29894
rect 96374 29883 96682 29892
rect 96374 28860 96682 28869
rect 96374 28858 96380 28860
rect 96436 28858 96460 28860
rect 96516 28858 96540 28860
rect 96596 28858 96620 28860
rect 96676 28858 96682 28860
rect 96436 28806 96438 28858
rect 96618 28806 96620 28858
rect 96374 28804 96380 28806
rect 96436 28804 96460 28806
rect 96516 28804 96540 28806
rect 96596 28804 96620 28806
rect 96676 28804 96682 28806
rect 96374 28795 96682 28804
rect 96374 27772 96682 27781
rect 96374 27770 96380 27772
rect 96436 27770 96460 27772
rect 96516 27770 96540 27772
rect 96596 27770 96620 27772
rect 96676 27770 96682 27772
rect 96436 27718 96438 27770
rect 96618 27718 96620 27770
rect 96374 27716 96380 27718
rect 96436 27716 96460 27718
rect 96516 27716 96540 27718
rect 96596 27716 96620 27718
rect 96676 27716 96682 27718
rect 96374 27707 96682 27716
rect 96374 26684 96682 26693
rect 96374 26682 96380 26684
rect 96436 26682 96460 26684
rect 96516 26682 96540 26684
rect 96596 26682 96620 26684
rect 96676 26682 96682 26684
rect 96436 26630 96438 26682
rect 96618 26630 96620 26682
rect 96374 26628 96380 26630
rect 96436 26628 96460 26630
rect 96516 26628 96540 26630
rect 96596 26628 96620 26630
rect 96676 26628 96682 26630
rect 96374 26619 96682 26628
rect 96374 25596 96682 25605
rect 96374 25594 96380 25596
rect 96436 25594 96460 25596
rect 96516 25594 96540 25596
rect 96596 25594 96620 25596
rect 96676 25594 96682 25596
rect 96436 25542 96438 25594
rect 96618 25542 96620 25594
rect 96374 25540 96380 25542
rect 96436 25540 96460 25542
rect 96516 25540 96540 25542
rect 96596 25540 96620 25542
rect 96676 25540 96682 25542
rect 96374 25531 96682 25540
rect 96374 24508 96682 24517
rect 96374 24506 96380 24508
rect 96436 24506 96460 24508
rect 96516 24506 96540 24508
rect 96596 24506 96620 24508
rect 96676 24506 96682 24508
rect 96436 24454 96438 24506
rect 96618 24454 96620 24506
rect 96374 24452 96380 24454
rect 96436 24452 96460 24454
rect 96516 24452 96540 24454
rect 96596 24452 96620 24454
rect 96676 24452 96682 24454
rect 96374 24443 96682 24452
rect 96374 23420 96682 23429
rect 96374 23418 96380 23420
rect 96436 23418 96460 23420
rect 96516 23418 96540 23420
rect 96596 23418 96620 23420
rect 96676 23418 96682 23420
rect 96436 23366 96438 23418
rect 96618 23366 96620 23418
rect 96374 23364 96380 23366
rect 96436 23364 96460 23366
rect 96516 23364 96540 23366
rect 96596 23364 96620 23366
rect 96676 23364 96682 23366
rect 96374 23355 96682 23364
rect 96374 22332 96682 22341
rect 96374 22330 96380 22332
rect 96436 22330 96460 22332
rect 96516 22330 96540 22332
rect 96596 22330 96620 22332
rect 96676 22330 96682 22332
rect 96436 22278 96438 22330
rect 96618 22278 96620 22330
rect 96374 22276 96380 22278
rect 96436 22276 96460 22278
rect 96516 22276 96540 22278
rect 96596 22276 96620 22278
rect 96676 22276 96682 22278
rect 96374 22267 96682 22276
rect 96374 21244 96682 21253
rect 96374 21242 96380 21244
rect 96436 21242 96460 21244
rect 96516 21242 96540 21244
rect 96596 21242 96620 21244
rect 96676 21242 96682 21244
rect 96436 21190 96438 21242
rect 96618 21190 96620 21242
rect 96374 21188 96380 21190
rect 96436 21188 96460 21190
rect 96516 21188 96540 21190
rect 96596 21188 96620 21190
rect 96676 21188 96682 21190
rect 96374 21179 96682 21188
rect 96374 20156 96682 20165
rect 96374 20154 96380 20156
rect 96436 20154 96460 20156
rect 96516 20154 96540 20156
rect 96596 20154 96620 20156
rect 96676 20154 96682 20156
rect 96436 20102 96438 20154
rect 96618 20102 96620 20154
rect 96374 20100 96380 20102
rect 96436 20100 96460 20102
rect 96516 20100 96540 20102
rect 96596 20100 96620 20102
rect 96676 20100 96682 20102
rect 96374 20091 96682 20100
rect 96374 19068 96682 19077
rect 96374 19066 96380 19068
rect 96436 19066 96460 19068
rect 96516 19066 96540 19068
rect 96596 19066 96620 19068
rect 96676 19066 96682 19068
rect 96436 19014 96438 19066
rect 96618 19014 96620 19066
rect 96374 19012 96380 19014
rect 96436 19012 96460 19014
rect 96516 19012 96540 19014
rect 96596 19012 96620 19014
rect 96676 19012 96682 19014
rect 96374 19003 96682 19012
rect 96374 17980 96682 17989
rect 96374 17978 96380 17980
rect 96436 17978 96460 17980
rect 96516 17978 96540 17980
rect 96596 17978 96620 17980
rect 96676 17978 96682 17980
rect 96436 17926 96438 17978
rect 96618 17926 96620 17978
rect 96374 17924 96380 17926
rect 96436 17924 96460 17926
rect 96516 17924 96540 17926
rect 96596 17924 96620 17926
rect 96676 17924 96682 17926
rect 96374 17915 96682 17924
rect 96374 16892 96682 16901
rect 96374 16890 96380 16892
rect 96436 16890 96460 16892
rect 96516 16890 96540 16892
rect 96596 16890 96620 16892
rect 96676 16890 96682 16892
rect 96436 16838 96438 16890
rect 96618 16838 96620 16890
rect 96374 16836 96380 16838
rect 96436 16836 96460 16838
rect 96516 16836 96540 16838
rect 96596 16836 96620 16838
rect 96676 16836 96682 16838
rect 96374 16827 96682 16836
rect 96374 15804 96682 15813
rect 96374 15802 96380 15804
rect 96436 15802 96460 15804
rect 96516 15802 96540 15804
rect 96596 15802 96620 15804
rect 96676 15802 96682 15804
rect 96436 15750 96438 15802
rect 96618 15750 96620 15802
rect 96374 15748 96380 15750
rect 96436 15748 96460 15750
rect 96516 15748 96540 15750
rect 96596 15748 96620 15750
rect 96676 15748 96682 15750
rect 96374 15739 96682 15748
rect 96374 14716 96682 14725
rect 96374 14714 96380 14716
rect 96436 14714 96460 14716
rect 96516 14714 96540 14716
rect 96596 14714 96620 14716
rect 96676 14714 96682 14716
rect 96436 14662 96438 14714
rect 96618 14662 96620 14714
rect 96374 14660 96380 14662
rect 96436 14660 96460 14662
rect 96516 14660 96540 14662
rect 96596 14660 96620 14662
rect 96676 14660 96682 14662
rect 96374 14651 96682 14660
rect 96374 13628 96682 13637
rect 96374 13626 96380 13628
rect 96436 13626 96460 13628
rect 96516 13626 96540 13628
rect 96596 13626 96620 13628
rect 96676 13626 96682 13628
rect 96436 13574 96438 13626
rect 96618 13574 96620 13626
rect 96374 13572 96380 13574
rect 96436 13572 96460 13574
rect 96516 13572 96540 13574
rect 96596 13572 96620 13574
rect 96676 13572 96682 13574
rect 96374 13563 96682 13572
rect 96374 12540 96682 12549
rect 96374 12538 96380 12540
rect 96436 12538 96460 12540
rect 96516 12538 96540 12540
rect 96596 12538 96620 12540
rect 96676 12538 96682 12540
rect 96436 12486 96438 12538
rect 96618 12486 96620 12538
rect 96374 12484 96380 12486
rect 96436 12484 96460 12486
rect 96516 12484 96540 12486
rect 96596 12484 96620 12486
rect 96676 12484 96682 12486
rect 96374 12475 96682 12484
rect 96374 11452 96682 11461
rect 96374 11450 96380 11452
rect 96436 11450 96460 11452
rect 96516 11450 96540 11452
rect 96596 11450 96620 11452
rect 96676 11450 96682 11452
rect 96436 11398 96438 11450
rect 96618 11398 96620 11450
rect 96374 11396 96380 11398
rect 96436 11396 96460 11398
rect 96516 11396 96540 11398
rect 96596 11396 96620 11398
rect 96676 11396 96682 11398
rect 96374 11387 96682 11396
rect 96374 10364 96682 10373
rect 96374 10362 96380 10364
rect 96436 10362 96460 10364
rect 96516 10362 96540 10364
rect 96596 10362 96620 10364
rect 96676 10362 96682 10364
rect 96436 10310 96438 10362
rect 96618 10310 96620 10362
rect 96374 10308 96380 10310
rect 96436 10308 96460 10310
rect 96516 10308 96540 10310
rect 96596 10308 96620 10310
rect 96676 10308 96682 10310
rect 96374 10299 96682 10308
rect 96374 9276 96682 9285
rect 96374 9274 96380 9276
rect 96436 9274 96460 9276
rect 96516 9274 96540 9276
rect 96596 9274 96620 9276
rect 96676 9274 96682 9276
rect 96436 9222 96438 9274
rect 96618 9222 96620 9274
rect 96374 9220 96380 9222
rect 96436 9220 96460 9222
rect 96516 9220 96540 9222
rect 96596 9220 96620 9222
rect 96676 9220 96682 9222
rect 96374 9211 96682 9220
rect 96374 8188 96682 8197
rect 96374 8186 96380 8188
rect 96436 8186 96460 8188
rect 96516 8186 96540 8188
rect 96596 8186 96620 8188
rect 96676 8186 96682 8188
rect 96436 8134 96438 8186
rect 96618 8134 96620 8186
rect 96374 8132 96380 8134
rect 96436 8132 96460 8134
rect 96516 8132 96540 8134
rect 96596 8132 96620 8134
rect 96676 8132 96682 8134
rect 96374 8123 96682 8132
rect 96374 7100 96682 7109
rect 96374 7098 96380 7100
rect 96436 7098 96460 7100
rect 96516 7098 96540 7100
rect 96596 7098 96620 7100
rect 96676 7098 96682 7100
rect 96436 7046 96438 7098
rect 96618 7046 96620 7098
rect 96374 7044 96380 7046
rect 96436 7044 96460 7046
rect 96516 7044 96540 7046
rect 96596 7044 96620 7046
rect 96676 7044 96682 7046
rect 96374 7035 96682 7044
rect 96374 6012 96682 6021
rect 96374 6010 96380 6012
rect 96436 6010 96460 6012
rect 96516 6010 96540 6012
rect 96596 6010 96620 6012
rect 96676 6010 96682 6012
rect 96436 5958 96438 6010
rect 96618 5958 96620 6010
rect 96374 5956 96380 5958
rect 96436 5956 96460 5958
rect 96516 5956 96540 5958
rect 96596 5956 96620 5958
rect 96676 5956 96682 5958
rect 96374 5947 96682 5956
rect 96374 4924 96682 4933
rect 96374 4922 96380 4924
rect 96436 4922 96460 4924
rect 96516 4922 96540 4924
rect 96596 4922 96620 4924
rect 96676 4922 96682 4924
rect 96436 4870 96438 4922
rect 96618 4870 96620 4922
rect 96374 4868 96380 4870
rect 96436 4868 96460 4870
rect 96516 4868 96540 4870
rect 96596 4868 96620 4870
rect 96676 4868 96682 4870
rect 96374 4859 96682 4868
rect 96374 3836 96682 3845
rect 96374 3834 96380 3836
rect 96436 3834 96460 3836
rect 96516 3834 96540 3836
rect 96596 3834 96620 3836
rect 96676 3834 96682 3836
rect 96436 3782 96438 3834
rect 96618 3782 96620 3834
rect 96374 3780 96380 3782
rect 96436 3780 96460 3782
rect 96516 3780 96540 3782
rect 96596 3780 96620 3782
rect 96676 3780 96682 3782
rect 96374 3771 96682 3780
rect 97724 2848 97776 2854
rect 97724 2790 97776 2796
rect 96374 2748 96682 2757
rect 96374 2746 96380 2748
rect 96436 2746 96460 2748
rect 96516 2746 96540 2748
rect 96596 2746 96620 2748
rect 96676 2746 96682 2748
rect 96436 2694 96438 2746
rect 96618 2694 96620 2746
rect 96374 2692 96380 2694
rect 96436 2692 96460 2694
rect 96516 2692 96540 2694
rect 96596 2692 96620 2694
rect 96676 2692 96682 2694
rect 96374 2683 96682 2692
rect 89720 2644 89772 2650
rect 89720 2586 89772 2592
rect 94320 2644 94372 2650
rect 94320 2586 94372 2592
rect 97736 2378 97764 2790
rect 97828 2650 97856 35974
rect 98012 32774 98040 36518
rect 98472 36258 98500 37198
rect 98552 37120 98604 37126
rect 98552 37062 98604 37068
rect 98564 36854 98592 37062
rect 98552 36848 98604 36854
rect 98552 36790 98604 36796
rect 98656 36582 98684 39222
rect 99286 39200 99342 40000
rect 100206 39200 100262 40000
rect 100312 39222 100708 39250
rect 99300 37262 99328 39200
rect 100220 39114 100248 39200
rect 100312 39114 100340 39222
rect 100220 39086 100340 39114
rect 99472 37868 99524 37874
rect 99472 37810 99524 37816
rect 99484 37466 99512 37810
rect 99472 37460 99524 37466
rect 99472 37402 99524 37408
rect 99472 37324 99524 37330
rect 99472 37266 99524 37272
rect 99288 37256 99340 37262
rect 99288 37198 99340 37204
rect 98736 37188 98788 37194
rect 98736 37130 98788 37136
rect 99380 37188 99432 37194
rect 99380 37130 99432 37136
rect 98748 36854 98776 37130
rect 99392 36854 99420 37130
rect 98736 36848 98788 36854
rect 98736 36790 98788 36796
rect 99380 36848 99432 36854
rect 99380 36790 99432 36796
rect 98644 36576 98696 36582
rect 98644 36518 98696 36524
rect 98380 36230 98500 36258
rect 98380 36038 98408 36230
rect 99484 36174 99512 37266
rect 99840 37256 99892 37262
rect 99840 37198 99892 37204
rect 100576 37256 100628 37262
rect 100576 37198 100628 37204
rect 99852 36854 99880 37198
rect 100208 37120 100260 37126
rect 100208 37062 100260 37068
rect 99840 36848 99892 36854
rect 99840 36790 99892 36796
rect 100220 36689 100248 37062
rect 100206 36680 100262 36689
rect 100206 36615 100262 36624
rect 99380 36168 99432 36174
rect 98472 36106 98684 36122
rect 99380 36110 99432 36116
rect 99472 36168 99524 36174
rect 99472 36110 99524 36116
rect 98460 36100 98696 36106
rect 98512 36094 98644 36100
rect 98460 36042 98512 36048
rect 98644 36042 98696 36048
rect 99392 36038 99420 36110
rect 100588 36038 100616 37198
rect 100680 37108 100708 39222
rect 101126 39200 101182 40000
rect 102046 39200 102102 40000
rect 102966 39200 103022 40000
rect 103886 39200 103942 40000
rect 104806 39200 104862 40000
rect 105726 39200 105782 40000
rect 106646 39200 106702 40000
rect 107566 39200 107622 40000
rect 108486 39200 108542 40000
rect 109406 39200 109462 40000
rect 110326 39200 110382 40000
rect 111246 39200 111302 40000
rect 111352 39222 111656 39250
rect 100760 37120 100812 37126
rect 100680 37080 100760 37108
rect 100760 37062 100812 37068
rect 100760 36780 100812 36786
rect 100760 36722 100812 36728
rect 100772 36582 100800 36722
rect 101140 36582 101168 39200
rect 101956 37936 102008 37942
rect 101956 37878 102008 37884
rect 101968 37466 101996 37878
rect 101956 37460 102008 37466
rect 101956 37402 102008 37408
rect 102060 37330 102088 39200
rect 102048 37324 102100 37330
rect 102048 37266 102100 37272
rect 102784 37256 102836 37262
rect 102784 37198 102836 37204
rect 102876 37256 102928 37262
rect 102876 37198 102928 37204
rect 102140 37188 102192 37194
rect 102140 37130 102192 37136
rect 102152 36582 102180 37130
rect 102796 37126 102824 37198
rect 102692 37120 102744 37126
rect 102692 37062 102744 37068
rect 102784 37120 102836 37126
rect 102784 37062 102836 37068
rect 100760 36576 100812 36582
rect 100760 36518 100812 36524
rect 101128 36576 101180 36582
rect 101128 36518 101180 36524
rect 102140 36576 102192 36582
rect 102140 36518 102192 36524
rect 98368 36032 98420 36038
rect 98368 35974 98420 35980
rect 99380 36032 99432 36038
rect 99380 35974 99432 35980
rect 100576 36032 100628 36038
rect 100576 35974 100628 35980
rect 98380 35601 98408 35974
rect 98366 35592 98422 35601
rect 98366 35527 98422 35536
rect 98000 32768 98052 32774
rect 98000 32710 98052 32716
rect 100772 32570 100800 36518
rect 100760 32564 100812 32570
rect 100760 32506 100812 32512
rect 101864 2848 101916 2854
rect 101864 2790 101916 2796
rect 97816 2644 97868 2650
rect 97816 2586 97868 2592
rect 101876 2378 101904 2790
rect 102152 2650 102180 36518
rect 102704 36145 102732 37062
rect 102888 36854 102916 37198
rect 102876 36848 102928 36854
rect 102876 36790 102928 36796
rect 102980 36582 103008 39200
rect 103428 37188 103480 37194
rect 103428 37130 103480 37136
rect 103060 36780 103112 36786
rect 103060 36722 103112 36728
rect 102968 36576 103020 36582
rect 102968 36518 103020 36524
rect 103072 36378 103100 36722
rect 103440 36378 103468 37130
rect 103900 37126 103928 39200
rect 104440 37256 104492 37262
rect 104440 37198 104492 37204
rect 104820 37210 104848 39200
rect 105268 38752 105320 38758
rect 105268 38694 105320 38700
rect 104900 37256 104952 37262
rect 104820 37204 104900 37210
rect 104820 37198 104952 37204
rect 103888 37120 103940 37126
rect 103888 37062 103940 37068
rect 104452 36582 104480 37198
rect 104820 37182 104940 37198
rect 104440 36576 104492 36582
rect 104440 36518 104492 36524
rect 102876 36372 102928 36378
rect 102876 36314 102928 36320
rect 103060 36372 103112 36378
rect 103060 36314 103112 36320
rect 103428 36372 103480 36378
rect 103428 36314 103480 36320
rect 102690 36136 102746 36145
rect 102690 36071 102746 36080
rect 102888 34746 102916 36314
rect 102876 34740 102928 34746
rect 102876 34682 102928 34688
rect 104452 32502 104480 36518
rect 104912 36378 104940 37182
rect 105280 36854 105308 38694
rect 105360 37120 105412 37126
rect 105360 37062 105412 37068
rect 105268 36848 105320 36854
rect 105268 36790 105320 36796
rect 104900 36372 104952 36378
rect 104900 36314 104952 36320
rect 105372 36281 105400 37062
rect 105740 36582 105768 39200
rect 105912 37324 105964 37330
rect 105912 37266 105964 37272
rect 105728 36576 105780 36582
rect 105728 36518 105780 36524
rect 105358 36272 105414 36281
rect 105358 36207 105414 36216
rect 105636 36168 105688 36174
rect 105688 36116 105860 36122
rect 105636 36110 105860 36116
rect 105648 36094 105860 36110
rect 105832 36038 105860 36094
rect 105820 36032 105872 36038
rect 105820 35974 105872 35980
rect 105924 33862 105952 37266
rect 106660 37262 106688 39200
rect 106648 37256 106700 37262
rect 106648 37198 106700 37204
rect 107292 37256 107344 37262
rect 107292 37198 107344 37204
rect 106556 37120 106608 37126
rect 106556 37062 106608 37068
rect 107108 37120 107160 37126
rect 107108 37062 107160 37068
rect 106464 36848 106516 36854
rect 106464 36790 106516 36796
rect 106372 36780 106424 36786
rect 106372 36722 106424 36728
rect 106384 36378 106412 36722
rect 106372 36372 106424 36378
rect 106292 36332 106372 36360
rect 105912 33856 105964 33862
rect 105912 33798 105964 33804
rect 104440 32496 104492 32502
rect 104440 32438 104492 32444
rect 106292 32434 106320 36332
rect 106372 36314 106424 36320
rect 106476 36242 106504 36790
rect 106568 36378 106596 37062
rect 107120 36825 107148 37062
rect 107304 36854 107332 37198
rect 107580 37108 107608 39200
rect 108500 37262 108528 39200
rect 107752 37256 107804 37262
rect 107752 37198 107804 37204
rect 108488 37256 108540 37262
rect 108488 37198 108540 37204
rect 107660 37120 107712 37126
rect 107580 37080 107660 37108
rect 107660 37062 107712 37068
rect 107292 36848 107344 36854
rect 107106 36816 107162 36825
rect 107292 36790 107344 36796
rect 107106 36751 107162 36760
rect 107568 36780 107620 36786
rect 107568 36722 107620 36728
rect 107580 36378 107608 36722
rect 107764 36378 107792 37198
rect 108500 36854 108528 37198
rect 109420 37126 109448 39200
rect 110236 37664 110288 37670
rect 110236 37606 110288 37612
rect 110248 37330 110276 37606
rect 110236 37324 110288 37330
rect 110236 37266 110288 37272
rect 109592 37256 109644 37262
rect 109592 37198 109644 37204
rect 110340 37210 110368 39200
rect 111260 39114 111288 39200
rect 111352 39114 111380 39222
rect 111260 39086 111380 39114
rect 111248 38276 111300 38282
rect 111248 38218 111300 38224
rect 110696 37256 110748 37262
rect 110340 37204 110696 37210
rect 110340 37198 110748 37204
rect 108764 37120 108816 37126
rect 108764 37062 108816 37068
rect 109408 37120 109460 37126
rect 109408 37062 109460 37068
rect 108488 36848 108540 36854
rect 108488 36790 108540 36796
rect 108304 36712 108356 36718
rect 108304 36654 108356 36660
rect 106556 36372 106608 36378
rect 106556 36314 106608 36320
rect 107568 36372 107620 36378
rect 107568 36314 107620 36320
rect 107752 36372 107804 36378
rect 107752 36314 107804 36320
rect 106464 36236 106516 36242
rect 106464 36178 106516 36184
rect 106280 32428 106332 32434
rect 106280 32370 106332 32376
rect 106476 26234 106504 36178
rect 107764 34066 107792 36314
rect 108316 36242 108344 36654
rect 108304 36236 108356 36242
rect 108304 36178 108356 36184
rect 107752 34060 107804 34066
rect 107752 34002 107804 34008
rect 108776 32910 108804 37062
rect 109406 36816 109462 36825
rect 109406 36751 109462 36760
rect 109420 36582 109448 36751
rect 109604 36582 109632 37198
rect 110340 37182 110736 37198
rect 110420 37120 110472 37126
rect 110420 37062 110472 37068
rect 110432 36768 110460 37062
rect 110512 36780 110564 36786
rect 110432 36740 110512 36768
rect 110512 36722 110564 36728
rect 110524 36582 110552 36722
rect 109408 36576 109460 36582
rect 109408 36518 109460 36524
rect 109592 36576 109644 36582
rect 109592 36518 109644 36524
rect 110512 36576 110564 36582
rect 110512 36518 110564 36524
rect 109604 33998 109632 36518
rect 110234 36408 110290 36417
rect 110234 36343 110290 36352
rect 110248 36038 110276 36343
rect 110236 36032 110288 36038
rect 110236 35974 110288 35980
rect 109592 33992 109644 33998
rect 109592 33934 109644 33940
rect 108764 32904 108816 32910
rect 108764 32846 108816 32852
rect 106292 26206 106504 26234
rect 104532 3664 104584 3670
rect 104532 3606 104584 3612
rect 104544 3058 104572 3606
rect 104532 3052 104584 3058
rect 104532 2994 104584 3000
rect 102140 2644 102192 2650
rect 102140 2586 102192 2592
rect 104544 2446 104572 2994
rect 106292 2650 106320 26206
rect 108304 3460 108356 3466
rect 108304 3402 108356 3408
rect 106280 2644 106332 2650
rect 106280 2586 106332 2592
rect 108316 2514 108344 3402
rect 110420 2848 110472 2854
rect 110420 2790 110472 2796
rect 108764 2576 108816 2582
rect 108764 2518 108816 2524
rect 108304 2508 108356 2514
rect 108304 2450 108356 2456
rect 104532 2440 104584 2446
rect 104532 2382 104584 2388
rect 89444 2372 89496 2378
rect 89444 2314 89496 2320
rect 97724 2372 97776 2378
rect 97724 2314 97776 2320
rect 101864 2372 101916 2378
rect 101864 2314 101916 2320
rect 106004 2372 106056 2378
rect 106004 2314 106056 2320
rect 85672 2304 85724 2310
rect 85672 2246 85724 2252
rect 87604 2304 87656 2310
rect 87604 2246 87656 2252
rect 88064 2304 88116 2310
rect 88064 2246 88116 2252
rect 87616 1630 87644 2246
rect 87604 1624 87656 1630
rect 87604 1566 87656 1572
rect 88076 800 88104 2246
rect 89456 800 89484 2314
rect 91744 2304 91796 2310
rect 91744 2246 91796 2252
rect 92204 2304 92256 2310
rect 92204 2246 92256 2252
rect 93584 2304 93636 2310
rect 93584 2246 93636 2252
rect 96068 2304 96120 2310
rect 96068 2246 96120 2252
rect 96344 2304 96396 2310
rect 96344 2246 96396 2252
rect 91756 2038 91784 2246
rect 91744 2032 91796 2038
rect 91744 1974 91796 1980
rect 92216 800 92244 2246
rect 93596 800 93624 2246
rect 96080 2106 96108 2246
rect 96068 2100 96120 2106
rect 96068 2042 96120 2048
rect 96356 800 96384 2246
rect 97736 800 97764 2314
rect 100024 2304 100076 2310
rect 100024 2246 100076 2252
rect 100484 2304 100536 2310
rect 100484 2246 100536 2252
rect 100036 1970 100064 2246
rect 100024 1964 100076 1970
rect 100024 1906 100076 1912
rect 100496 800 100524 2246
rect 101876 800 101904 2314
rect 104624 2304 104676 2310
rect 104624 2246 104676 2252
rect 104636 800 104664 2246
rect 106016 800 106044 2314
rect 108776 800 108804 2518
rect 110432 2378 110460 2790
rect 110524 2650 110552 36518
rect 110708 36378 110736 37182
rect 111260 37126 111288 38218
rect 111248 37120 111300 37126
rect 111628 37108 111656 39222
rect 112166 39200 112222 40000
rect 113086 39200 113142 40000
rect 114006 39200 114062 40000
rect 114926 39200 114982 40000
rect 115846 39200 115902 40000
rect 116766 39200 116822 40000
rect 116872 39222 117268 39250
rect 112180 37346 112208 39200
rect 112996 38412 113048 38418
rect 112996 38354 113048 38360
rect 112180 37318 112300 37346
rect 112272 37262 112300 37318
rect 112168 37256 112220 37262
rect 112168 37198 112220 37204
rect 112260 37256 112312 37262
rect 112260 37198 112312 37204
rect 112720 37256 112772 37262
rect 112720 37198 112772 37204
rect 111800 37120 111852 37126
rect 111628 37080 111800 37108
rect 111248 37062 111300 37068
rect 111800 37062 111852 37068
rect 111734 37020 112042 37029
rect 111734 37018 111740 37020
rect 111796 37018 111820 37020
rect 111876 37018 111900 37020
rect 111956 37018 111980 37020
rect 112036 37018 112042 37020
rect 111796 36966 111798 37018
rect 111978 36966 111980 37018
rect 111734 36964 111740 36966
rect 111796 36964 111820 36966
rect 111876 36964 111900 36966
rect 111956 36964 111980 36966
rect 112036 36964 112042 36966
rect 111734 36955 112042 36964
rect 112076 36780 112128 36786
rect 112076 36722 112128 36728
rect 111890 36680 111946 36689
rect 111890 36615 111946 36624
rect 111904 36582 111932 36615
rect 111892 36576 111944 36582
rect 111892 36518 111944 36524
rect 110696 36372 110748 36378
rect 110696 36314 110748 36320
rect 111734 35932 112042 35941
rect 111734 35930 111740 35932
rect 111796 35930 111820 35932
rect 111876 35930 111900 35932
rect 111956 35930 111980 35932
rect 112036 35930 112042 35932
rect 111796 35878 111798 35930
rect 111978 35878 111980 35930
rect 111734 35876 111740 35878
rect 111796 35876 111820 35878
rect 111876 35876 111900 35878
rect 111956 35876 111980 35878
rect 112036 35876 112042 35878
rect 111734 35867 112042 35876
rect 112088 35766 112116 36722
rect 112180 36038 112208 37198
rect 112536 36848 112588 36854
rect 112536 36790 112588 36796
rect 112352 36372 112404 36378
rect 112352 36314 112404 36320
rect 112364 36174 112392 36314
rect 112548 36174 112576 36790
rect 112352 36168 112404 36174
rect 112352 36110 112404 36116
rect 112536 36168 112588 36174
rect 112536 36110 112588 36116
rect 112732 36038 112760 37198
rect 113008 37126 113036 38354
rect 112996 37120 113048 37126
rect 113100 37108 113128 39200
rect 113732 38684 113784 38690
rect 113732 38626 113784 38632
rect 113456 37256 113508 37262
rect 113456 37198 113508 37204
rect 113180 37120 113232 37126
rect 113100 37080 113180 37108
rect 112996 37062 113048 37068
rect 113180 37062 113232 37068
rect 113468 36038 113496 37198
rect 113744 36786 113772 38626
rect 114020 37262 114048 39200
rect 114008 37256 114060 37262
rect 114008 37198 114060 37204
rect 114836 37256 114888 37262
rect 114836 37198 114888 37204
rect 114560 37120 114612 37126
rect 114560 37062 114612 37068
rect 113732 36780 113784 36786
rect 113732 36722 113784 36728
rect 112168 36032 112220 36038
rect 112168 35974 112220 35980
rect 112720 36032 112772 36038
rect 112720 35974 112772 35980
rect 113456 36032 113508 36038
rect 113456 35974 113508 35980
rect 112076 35760 112128 35766
rect 112076 35702 112128 35708
rect 111734 34844 112042 34853
rect 111734 34842 111740 34844
rect 111796 34842 111820 34844
rect 111876 34842 111900 34844
rect 111956 34842 111980 34844
rect 112036 34842 112042 34844
rect 111796 34790 111798 34842
rect 111978 34790 111980 34842
rect 111734 34788 111740 34790
rect 111796 34788 111820 34790
rect 111876 34788 111900 34790
rect 111956 34788 111980 34790
rect 112036 34788 112042 34790
rect 111734 34779 112042 34788
rect 112180 33930 112208 35974
rect 113468 34202 113496 35974
rect 113456 34196 113508 34202
rect 113456 34138 113508 34144
rect 112168 33924 112220 33930
rect 112168 33866 112220 33872
rect 111734 33756 112042 33765
rect 111734 33754 111740 33756
rect 111796 33754 111820 33756
rect 111876 33754 111900 33756
rect 111956 33754 111980 33756
rect 112036 33754 112042 33756
rect 111796 33702 111798 33754
rect 111978 33702 111980 33754
rect 111734 33700 111740 33702
rect 111796 33700 111820 33702
rect 111876 33700 111900 33702
rect 111956 33700 111980 33702
rect 112036 33700 112042 33702
rect 111734 33691 112042 33700
rect 114572 33046 114600 37062
rect 114848 36938 114876 37198
rect 114940 37108 114968 39200
rect 115480 37256 115532 37262
rect 115480 37198 115532 37204
rect 115860 37210 115888 39200
rect 116780 39114 116808 39200
rect 116872 39114 116900 39222
rect 116780 39086 116900 39114
rect 116216 37800 116268 37806
rect 116216 37742 116268 37748
rect 116228 37330 116256 37742
rect 116216 37324 116268 37330
rect 116216 37266 116268 37272
rect 115940 37256 115992 37262
rect 115860 37204 115940 37210
rect 115860 37198 115992 37204
rect 116124 37256 116176 37262
rect 116124 37198 116176 37204
rect 117136 37256 117188 37262
rect 117136 37198 117188 37204
rect 115020 37120 115072 37126
rect 114940 37080 115020 37108
rect 115020 37062 115072 37068
rect 114848 36910 114968 36938
rect 114652 36780 114704 36786
rect 114652 36722 114704 36728
rect 114664 36038 114692 36722
rect 114940 36038 114968 36910
rect 115492 36378 115520 37198
rect 115860 37182 115980 37198
rect 116136 36854 116164 37198
rect 116124 36848 116176 36854
rect 116124 36790 116176 36796
rect 116308 36848 116360 36854
rect 116308 36790 116360 36796
rect 116032 36780 116084 36786
rect 116032 36722 116084 36728
rect 116044 36666 116072 36722
rect 115860 36638 116072 36666
rect 115860 36417 115888 36638
rect 115846 36408 115902 36417
rect 115480 36372 115532 36378
rect 115846 36343 115902 36352
rect 115480 36314 115532 36320
rect 116320 36242 116348 36790
rect 117148 36786 117176 37198
rect 117240 37108 117268 39222
rect 117686 39200 117742 40000
rect 118606 39200 118662 40000
rect 119526 39200 119582 40000
rect 120446 39200 120502 40000
rect 121366 39200 121422 40000
rect 122286 39200 122342 40000
rect 122392 39222 122696 39250
rect 117700 37194 117728 39200
rect 118056 39092 118108 39098
rect 118056 39034 118108 39040
rect 117872 38616 117924 38622
rect 117872 38558 117924 38564
rect 117688 37188 117740 37194
rect 117688 37130 117740 37136
rect 117320 37120 117372 37126
rect 117240 37080 117320 37108
rect 117320 37062 117372 37068
rect 117136 36780 117188 36786
rect 117136 36722 117188 36728
rect 116952 36576 117004 36582
rect 116952 36518 117004 36524
rect 116308 36236 116360 36242
rect 116308 36178 116360 36184
rect 116964 36038 116992 36518
rect 117700 36378 117728 37130
rect 117884 36786 117912 38558
rect 118068 37330 118096 39034
rect 118056 37324 118108 37330
rect 118056 37266 118108 37272
rect 118620 37108 118648 39200
rect 119540 37262 119568 39200
rect 120080 38548 120132 38554
rect 120080 38490 120132 38496
rect 119896 37664 119948 37670
rect 119896 37606 119948 37612
rect 119908 37466 119936 37606
rect 120092 37466 120120 38490
rect 120460 37466 120488 39200
rect 120632 37732 120684 37738
rect 120632 37674 120684 37680
rect 119896 37460 119948 37466
rect 119896 37402 119948 37408
rect 120080 37460 120132 37466
rect 120080 37402 120132 37408
rect 120448 37460 120500 37466
rect 120448 37402 120500 37408
rect 120644 37330 120672 37674
rect 120632 37324 120684 37330
rect 120632 37266 120684 37272
rect 119160 37256 119212 37262
rect 119160 37198 119212 37204
rect 119528 37256 119580 37262
rect 119528 37198 119580 37204
rect 119896 37256 119948 37262
rect 119896 37198 119948 37204
rect 118700 37120 118752 37126
rect 118620 37080 118700 37108
rect 118700 37062 118752 37068
rect 117872 36780 117924 36786
rect 117872 36722 117924 36728
rect 118700 36780 118752 36786
rect 118700 36722 118752 36728
rect 117688 36372 117740 36378
rect 117688 36314 117740 36320
rect 114652 36032 114704 36038
rect 114652 35974 114704 35980
rect 114928 36032 114980 36038
rect 114928 35974 114980 35980
rect 116952 36032 117004 36038
rect 116952 35974 117004 35980
rect 114560 33040 114612 33046
rect 114560 32982 114612 32988
rect 111734 32668 112042 32677
rect 111734 32666 111740 32668
rect 111796 32666 111820 32668
rect 111876 32666 111900 32668
rect 111956 32666 111980 32668
rect 112036 32666 112042 32668
rect 111796 32614 111798 32666
rect 111978 32614 111980 32666
rect 111734 32612 111740 32614
rect 111796 32612 111820 32614
rect 111876 32612 111900 32614
rect 111956 32612 111980 32614
rect 112036 32612 112042 32614
rect 111734 32603 112042 32612
rect 114664 31754 114692 35974
rect 114664 31726 114876 31754
rect 111734 31580 112042 31589
rect 111734 31578 111740 31580
rect 111796 31578 111820 31580
rect 111876 31578 111900 31580
rect 111956 31578 111980 31580
rect 112036 31578 112042 31580
rect 111796 31526 111798 31578
rect 111978 31526 111980 31578
rect 111734 31524 111740 31526
rect 111796 31524 111820 31526
rect 111876 31524 111900 31526
rect 111956 31524 111980 31526
rect 112036 31524 112042 31526
rect 111734 31515 112042 31524
rect 111734 30492 112042 30501
rect 111734 30490 111740 30492
rect 111796 30490 111820 30492
rect 111876 30490 111900 30492
rect 111956 30490 111980 30492
rect 112036 30490 112042 30492
rect 111796 30438 111798 30490
rect 111978 30438 111980 30490
rect 111734 30436 111740 30438
rect 111796 30436 111820 30438
rect 111876 30436 111900 30438
rect 111956 30436 111980 30438
rect 112036 30436 112042 30438
rect 111734 30427 112042 30436
rect 111734 29404 112042 29413
rect 111734 29402 111740 29404
rect 111796 29402 111820 29404
rect 111876 29402 111900 29404
rect 111956 29402 111980 29404
rect 112036 29402 112042 29404
rect 111796 29350 111798 29402
rect 111978 29350 111980 29402
rect 111734 29348 111740 29350
rect 111796 29348 111820 29350
rect 111876 29348 111900 29350
rect 111956 29348 111980 29350
rect 112036 29348 112042 29350
rect 111734 29339 112042 29348
rect 111734 28316 112042 28325
rect 111734 28314 111740 28316
rect 111796 28314 111820 28316
rect 111876 28314 111900 28316
rect 111956 28314 111980 28316
rect 112036 28314 112042 28316
rect 111796 28262 111798 28314
rect 111978 28262 111980 28314
rect 111734 28260 111740 28262
rect 111796 28260 111820 28262
rect 111876 28260 111900 28262
rect 111956 28260 111980 28262
rect 112036 28260 112042 28262
rect 111734 28251 112042 28260
rect 111734 27228 112042 27237
rect 111734 27226 111740 27228
rect 111796 27226 111820 27228
rect 111876 27226 111900 27228
rect 111956 27226 111980 27228
rect 112036 27226 112042 27228
rect 111796 27174 111798 27226
rect 111978 27174 111980 27226
rect 111734 27172 111740 27174
rect 111796 27172 111820 27174
rect 111876 27172 111900 27174
rect 111956 27172 111980 27174
rect 112036 27172 112042 27174
rect 111734 27163 112042 27172
rect 111734 26140 112042 26149
rect 111734 26138 111740 26140
rect 111796 26138 111820 26140
rect 111876 26138 111900 26140
rect 111956 26138 111980 26140
rect 112036 26138 112042 26140
rect 111796 26086 111798 26138
rect 111978 26086 111980 26138
rect 111734 26084 111740 26086
rect 111796 26084 111820 26086
rect 111876 26084 111900 26086
rect 111956 26084 111980 26086
rect 112036 26084 112042 26086
rect 111734 26075 112042 26084
rect 111734 25052 112042 25061
rect 111734 25050 111740 25052
rect 111796 25050 111820 25052
rect 111876 25050 111900 25052
rect 111956 25050 111980 25052
rect 112036 25050 112042 25052
rect 111796 24998 111798 25050
rect 111978 24998 111980 25050
rect 111734 24996 111740 24998
rect 111796 24996 111820 24998
rect 111876 24996 111900 24998
rect 111956 24996 111980 24998
rect 112036 24996 112042 24998
rect 111734 24987 112042 24996
rect 111734 23964 112042 23973
rect 111734 23962 111740 23964
rect 111796 23962 111820 23964
rect 111876 23962 111900 23964
rect 111956 23962 111980 23964
rect 112036 23962 112042 23964
rect 111796 23910 111798 23962
rect 111978 23910 111980 23962
rect 111734 23908 111740 23910
rect 111796 23908 111820 23910
rect 111876 23908 111900 23910
rect 111956 23908 111980 23910
rect 112036 23908 112042 23910
rect 111734 23899 112042 23908
rect 111734 22876 112042 22885
rect 111734 22874 111740 22876
rect 111796 22874 111820 22876
rect 111876 22874 111900 22876
rect 111956 22874 111980 22876
rect 112036 22874 112042 22876
rect 111796 22822 111798 22874
rect 111978 22822 111980 22874
rect 111734 22820 111740 22822
rect 111796 22820 111820 22822
rect 111876 22820 111900 22822
rect 111956 22820 111980 22822
rect 112036 22820 112042 22822
rect 111734 22811 112042 22820
rect 111734 21788 112042 21797
rect 111734 21786 111740 21788
rect 111796 21786 111820 21788
rect 111876 21786 111900 21788
rect 111956 21786 111980 21788
rect 112036 21786 112042 21788
rect 111796 21734 111798 21786
rect 111978 21734 111980 21786
rect 111734 21732 111740 21734
rect 111796 21732 111820 21734
rect 111876 21732 111900 21734
rect 111956 21732 111980 21734
rect 112036 21732 112042 21734
rect 111734 21723 112042 21732
rect 111734 20700 112042 20709
rect 111734 20698 111740 20700
rect 111796 20698 111820 20700
rect 111876 20698 111900 20700
rect 111956 20698 111980 20700
rect 112036 20698 112042 20700
rect 111796 20646 111798 20698
rect 111978 20646 111980 20698
rect 111734 20644 111740 20646
rect 111796 20644 111820 20646
rect 111876 20644 111900 20646
rect 111956 20644 111980 20646
rect 112036 20644 112042 20646
rect 111734 20635 112042 20644
rect 111734 19612 112042 19621
rect 111734 19610 111740 19612
rect 111796 19610 111820 19612
rect 111876 19610 111900 19612
rect 111956 19610 111980 19612
rect 112036 19610 112042 19612
rect 111796 19558 111798 19610
rect 111978 19558 111980 19610
rect 111734 19556 111740 19558
rect 111796 19556 111820 19558
rect 111876 19556 111900 19558
rect 111956 19556 111980 19558
rect 112036 19556 112042 19558
rect 111734 19547 112042 19556
rect 111734 18524 112042 18533
rect 111734 18522 111740 18524
rect 111796 18522 111820 18524
rect 111876 18522 111900 18524
rect 111956 18522 111980 18524
rect 112036 18522 112042 18524
rect 111796 18470 111798 18522
rect 111978 18470 111980 18522
rect 111734 18468 111740 18470
rect 111796 18468 111820 18470
rect 111876 18468 111900 18470
rect 111956 18468 111980 18470
rect 112036 18468 112042 18470
rect 111734 18459 112042 18468
rect 111734 17436 112042 17445
rect 111734 17434 111740 17436
rect 111796 17434 111820 17436
rect 111876 17434 111900 17436
rect 111956 17434 111980 17436
rect 112036 17434 112042 17436
rect 111796 17382 111798 17434
rect 111978 17382 111980 17434
rect 111734 17380 111740 17382
rect 111796 17380 111820 17382
rect 111876 17380 111900 17382
rect 111956 17380 111980 17382
rect 112036 17380 112042 17382
rect 111734 17371 112042 17380
rect 111734 16348 112042 16357
rect 111734 16346 111740 16348
rect 111796 16346 111820 16348
rect 111876 16346 111900 16348
rect 111956 16346 111980 16348
rect 112036 16346 112042 16348
rect 111796 16294 111798 16346
rect 111978 16294 111980 16346
rect 111734 16292 111740 16294
rect 111796 16292 111820 16294
rect 111876 16292 111900 16294
rect 111956 16292 111980 16294
rect 112036 16292 112042 16294
rect 111734 16283 112042 16292
rect 111734 15260 112042 15269
rect 111734 15258 111740 15260
rect 111796 15258 111820 15260
rect 111876 15258 111900 15260
rect 111956 15258 111980 15260
rect 112036 15258 112042 15260
rect 111796 15206 111798 15258
rect 111978 15206 111980 15258
rect 111734 15204 111740 15206
rect 111796 15204 111820 15206
rect 111876 15204 111900 15206
rect 111956 15204 111980 15206
rect 112036 15204 112042 15206
rect 111734 15195 112042 15204
rect 111734 14172 112042 14181
rect 111734 14170 111740 14172
rect 111796 14170 111820 14172
rect 111876 14170 111900 14172
rect 111956 14170 111980 14172
rect 112036 14170 112042 14172
rect 111796 14118 111798 14170
rect 111978 14118 111980 14170
rect 111734 14116 111740 14118
rect 111796 14116 111820 14118
rect 111876 14116 111900 14118
rect 111956 14116 111980 14118
rect 112036 14116 112042 14118
rect 111734 14107 112042 14116
rect 111734 13084 112042 13093
rect 111734 13082 111740 13084
rect 111796 13082 111820 13084
rect 111876 13082 111900 13084
rect 111956 13082 111980 13084
rect 112036 13082 112042 13084
rect 111796 13030 111798 13082
rect 111978 13030 111980 13082
rect 111734 13028 111740 13030
rect 111796 13028 111820 13030
rect 111876 13028 111900 13030
rect 111956 13028 111980 13030
rect 112036 13028 112042 13030
rect 111734 13019 112042 13028
rect 111734 11996 112042 12005
rect 111734 11994 111740 11996
rect 111796 11994 111820 11996
rect 111876 11994 111900 11996
rect 111956 11994 111980 11996
rect 112036 11994 112042 11996
rect 111796 11942 111798 11994
rect 111978 11942 111980 11994
rect 111734 11940 111740 11942
rect 111796 11940 111820 11942
rect 111876 11940 111900 11942
rect 111956 11940 111980 11942
rect 112036 11940 112042 11942
rect 111734 11931 112042 11940
rect 111734 10908 112042 10917
rect 111734 10906 111740 10908
rect 111796 10906 111820 10908
rect 111876 10906 111900 10908
rect 111956 10906 111980 10908
rect 112036 10906 112042 10908
rect 111796 10854 111798 10906
rect 111978 10854 111980 10906
rect 111734 10852 111740 10854
rect 111796 10852 111820 10854
rect 111876 10852 111900 10854
rect 111956 10852 111980 10854
rect 112036 10852 112042 10854
rect 111734 10843 112042 10852
rect 111734 9820 112042 9829
rect 111734 9818 111740 9820
rect 111796 9818 111820 9820
rect 111876 9818 111900 9820
rect 111956 9818 111980 9820
rect 112036 9818 112042 9820
rect 111796 9766 111798 9818
rect 111978 9766 111980 9818
rect 111734 9764 111740 9766
rect 111796 9764 111820 9766
rect 111876 9764 111900 9766
rect 111956 9764 111980 9766
rect 112036 9764 112042 9766
rect 111734 9755 112042 9764
rect 111734 8732 112042 8741
rect 111734 8730 111740 8732
rect 111796 8730 111820 8732
rect 111876 8730 111900 8732
rect 111956 8730 111980 8732
rect 112036 8730 112042 8732
rect 111796 8678 111798 8730
rect 111978 8678 111980 8730
rect 111734 8676 111740 8678
rect 111796 8676 111820 8678
rect 111876 8676 111900 8678
rect 111956 8676 111980 8678
rect 112036 8676 112042 8678
rect 111734 8667 112042 8676
rect 111734 7644 112042 7653
rect 111734 7642 111740 7644
rect 111796 7642 111820 7644
rect 111876 7642 111900 7644
rect 111956 7642 111980 7644
rect 112036 7642 112042 7644
rect 111796 7590 111798 7642
rect 111978 7590 111980 7642
rect 111734 7588 111740 7590
rect 111796 7588 111820 7590
rect 111876 7588 111900 7590
rect 111956 7588 111980 7590
rect 112036 7588 112042 7590
rect 111734 7579 112042 7588
rect 111734 6556 112042 6565
rect 111734 6554 111740 6556
rect 111796 6554 111820 6556
rect 111876 6554 111900 6556
rect 111956 6554 111980 6556
rect 112036 6554 112042 6556
rect 111796 6502 111798 6554
rect 111978 6502 111980 6554
rect 111734 6500 111740 6502
rect 111796 6500 111820 6502
rect 111876 6500 111900 6502
rect 111956 6500 111980 6502
rect 112036 6500 112042 6502
rect 111734 6491 112042 6500
rect 111734 5468 112042 5477
rect 111734 5466 111740 5468
rect 111796 5466 111820 5468
rect 111876 5466 111900 5468
rect 111956 5466 111980 5468
rect 112036 5466 112042 5468
rect 111796 5414 111798 5466
rect 111978 5414 111980 5466
rect 111734 5412 111740 5414
rect 111796 5412 111820 5414
rect 111876 5412 111900 5414
rect 111956 5412 111980 5414
rect 112036 5412 112042 5414
rect 111734 5403 112042 5412
rect 111734 4380 112042 4389
rect 111734 4378 111740 4380
rect 111796 4378 111820 4380
rect 111876 4378 111900 4380
rect 111956 4378 111980 4380
rect 112036 4378 112042 4380
rect 111796 4326 111798 4378
rect 111978 4326 111980 4378
rect 111734 4324 111740 4326
rect 111796 4324 111820 4326
rect 111876 4324 111900 4326
rect 111956 4324 111980 4326
rect 112036 4324 112042 4326
rect 111734 4315 112042 4324
rect 111734 3292 112042 3301
rect 111734 3290 111740 3292
rect 111796 3290 111820 3292
rect 111876 3290 111900 3292
rect 111956 3290 111980 3292
rect 112036 3290 112042 3292
rect 111796 3238 111798 3290
rect 111978 3238 111980 3290
rect 111734 3236 111740 3238
rect 111796 3236 111820 3238
rect 111876 3236 111900 3238
rect 111956 3236 111980 3238
rect 112036 3236 112042 3238
rect 111734 3227 112042 3236
rect 114848 2650 114876 31726
rect 117228 3936 117280 3942
rect 117228 3878 117280 3884
rect 110512 2644 110564 2650
rect 110512 2586 110564 2592
rect 114836 2644 114888 2650
rect 114836 2586 114888 2592
rect 117240 2582 117268 3878
rect 118424 2848 118476 2854
rect 118424 2790 118476 2796
rect 117228 2576 117280 2582
rect 117228 2518 117280 2524
rect 118436 2378 118464 2790
rect 118712 2650 118740 36722
rect 119172 36582 119200 37198
rect 119908 36922 119936 37198
rect 120816 37188 120868 37194
rect 120816 37130 120868 37136
rect 119712 36916 119764 36922
rect 119712 36858 119764 36864
rect 119896 36916 119948 36922
rect 119896 36858 119948 36864
rect 119988 36916 120040 36922
rect 119988 36858 120040 36864
rect 119160 36576 119212 36582
rect 119160 36518 119212 36524
rect 119172 36310 119200 36518
rect 119724 36378 119752 36858
rect 120000 36786 120028 36858
rect 119988 36780 120040 36786
rect 119988 36722 120040 36728
rect 119712 36372 119764 36378
rect 119712 36314 119764 36320
rect 120828 36310 120856 37130
rect 121380 36786 121408 39200
rect 122300 39114 122328 39200
rect 122392 39114 122420 39222
rect 122300 39086 122420 39114
rect 122564 38480 122616 38486
rect 122564 38422 122616 38428
rect 121460 38208 121512 38214
rect 121460 38150 121512 38156
rect 121368 36780 121420 36786
rect 121368 36722 121420 36728
rect 121472 36582 121500 38150
rect 122576 37466 122604 38422
rect 122564 37460 122616 37466
rect 122564 37402 122616 37408
rect 121736 37256 121788 37262
rect 121736 37198 121788 37204
rect 121748 36802 121776 37198
rect 122668 37108 122696 39222
rect 123206 39200 123262 40000
rect 124126 39200 124182 40000
rect 125046 39200 125102 40000
rect 125966 39200 126022 40000
rect 126886 39200 126942 40000
rect 127806 39200 127862 40000
rect 127912 39222 128308 39250
rect 123116 38888 123168 38894
rect 123116 38830 123168 38836
rect 123128 37262 123156 38830
rect 122932 37256 122984 37262
rect 122932 37198 122984 37204
rect 123116 37256 123168 37262
rect 123220 37244 123248 39200
rect 123484 37324 123536 37330
rect 123484 37266 123536 37272
rect 123300 37256 123352 37262
rect 123220 37216 123300 37244
rect 123116 37198 123168 37204
rect 123300 37198 123352 37204
rect 122840 37120 122892 37126
rect 122668 37080 122840 37108
rect 122840 37062 122892 37068
rect 122944 36938 122972 37198
rect 121564 36774 121776 36802
rect 122852 36910 122972 36938
rect 122852 36786 122880 36910
rect 122840 36780 122892 36786
rect 121460 36576 121512 36582
rect 121460 36518 121512 36524
rect 119160 36304 119212 36310
rect 119160 36246 119212 36252
rect 120816 36304 120868 36310
rect 120816 36246 120868 36252
rect 120908 36236 120960 36242
rect 120908 36178 120960 36184
rect 120920 36038 120948 36178
rect 121564 36038 121592 36774
rect 122840 36722 122892 36728
rect 122852 36582 122880 36722
rect 122840 36576 122892 36582
rect 122840 36518 122892 36524
rect 120908 36032 120960 36038
rect 120908 35974 120960 35980
rect 121552 36032 121604 36038
rect 121552 35974 121604 35980
rect 121564 35562 121592 35974
rect 121552 35556 121604 35562
rect 121552 35498 121604 35504
rect 122564 2848 122616 2854
rect 122564 2790 122616 2796
rect 118700 2644 118752 2650
rect 118700 2586 118752 2592
rect 122576 2378 122604 2790
rect 122852 2650 122880 36518
rect 123128 36038 123156 37198
rect 123300 36712 123352 36718
rect 123300 36654 123352 36660
rect 123312 36378 123340 36654
rect 123208 36372 123260 36378
rect 123208 36314 123260 36320
rect 123300 36372 123352 36378
rect 123300 36314 123352 36320
rect 123220 36038 123248 36314
rect 123116 36032 123168 36038
rect 123116 35974 123168 35980
rect 123208 36032 123260 36038
rect 123208 35974 123260 35980
rect 123496 35630 123524 37266
rect 124036 37120 124088 37126
rect 124140 37108 124168 39200
rect 124956 37868 125008 37874
rect 124956 37810 125008 37816
rect 124968 37262 124996 37810
rect 124404 37256 124456 37262
rect 124404 37198 124456 37204
rect 124956 37256 125008 37262
rect 125060 37244 125088 39200
rect 125876 38072 125928 38078
rect 125876 38014 125928 38020
rect 125888 37466 125916 38014
rect 125876 37460 125928 37466
rect 125876 37402 125928 37408
rect 125140 37256 125192 37262
rect 125060 37216 125140 37244
rect 124956 37198 125008 37204
rect 125140 37198 125192 37204
rect 125600 37256 125652 37262
rect 125600 37198 125652 37204
rect 124220 37120 124272 37126
rect 124140 37080 124220 37108
rect 124036 37062 124088 37068
rect 124220 37062 124272 37068
rect 123576 36916 123628 36922
rect 123576 36858 123628 36864
rect 123588 36582 123616 36858
rect 123576 36576 123628 36582
rect 123576 36518 123628 36524
rect 123484 35624 123536 35630
rect 123484 35566 123536 35572
rect 124048 34474 124076 37062
rect 124416 36922 124444 37198
rect 124968 36922 124996 37198
rect 125612 36922 125640 37198
rect 125980 37108 126008 39200
rect 126520 38344 126572 38350
rect 126520 38286 126572 38292
rect 126428 37664 126480 37670
rect 126428 37606 126480 37612
rect 126440 37262 126468 37606
rect 126428 37256 126480 37262
rect 126428 37198 126480 37204
rect 126060 37120 126112 37126
rect 125980 37080 126060 37108
rect 126060 37062 126112 37068
rect 124404 36916 124456 36922
rect 124404 36858 124456 36864
rect 124956 36916 125008 36922
rect 124956 36858 125008 36864
rect 125600 36916 125652 36922
rect 125600 36858 125652 36864
rect 126440 36310 126468 37198
rect 126532 36922 126560 38286
rect 126900 37244 126928 39200
rect 127820 39114 127848 39200
rect 127912 39114 127940 39222
rect 127820 39086 127940 39114
rect 127094 37564 127402 37573
rect 127094 37562 127100 37564
rect 127156 37562 127180 37564
rect 127236 37562 127260 37564
rect 127316 37562 127340 37564
rect 127396 37562 127402 37564
rect 127156 37510 127158 37562
rect 127338 37510 127340 37562
rect 127094 37508 127100 37510
rect 127156 37508 127180 37510
rect 127236 37508 127260 37510
rect 127316 37508 127340 37510
rect 127396 37508 127402 37510
rect 127094 37499 127402 37508
rect 126980 37256 127032 37262
rect 126900 37216 126980 37244
rect 126980 37198 127032 37204
rect 127716 37256 127768 37262
rect 127716 37198 127768 37204
rect 127728 36922 127756 37198
rect 127808 37120 127860 37126
rect 128280 37108 128308 39222
rect 128726 39200 128782 40000
rect 129646 39200 129702 40000
rect 130566 39200 130622 40000
rect 130672 39222 131068 39250
rect 128740 37262 128768 39200
rect 128452 37256 128504 37262
rect 128452 37198 128504 37204
rect 128728 37256 128780 37262
rect 128728 37198 128780 37204
rect 129556 37256 129608 37262
rect 129556 37198 129608 37204
rect 128360 37120 128412 37126
rect 128280 37080 128360 37108
rect 127808 37062 127860 37068
rect 128360 37062 128412 37068
rect 126520 36916 126572 36922
rect 126520 36858 126572 36864
rect 127716 36916 127768 36922
rect 127716 36858 127768 36864
rect 126980 36780 127032 36786
rect 126980 36722 127032 36728
rect 126992 36582 127020 36722
rect 127820 36650 127848 37062
rect 128464 36938 128492 37198
rect 128372 36922 128492 36938
rect 128740 36922 128768 37198
rect 129280 37120 129332 37126
rect 129280 37062 129332 37068
rect 128360 36916 128492 36922
rect 128412 36910 128492 36916
rect 128728 36916 128780 36922
rect 128360 36858 128412 36864
rect 128728 36858 128780 36864
rect 128372 36825 128400 36858
rect 128358 36816 128414 36825
rect 128358 36751 128414 36760
rect 127808 36644 127860 36650
rect 127808 36586 127860 36592
rect 126520 36576 126572 36582
rect 126520 36518 126572 36524
rect 126980 36576 127032 36582
rect 126980 36518 127032 36524
rect 126532 36310 126560 36518
rect 126428 36304 126480 36310
rect 124218 36272 124274 36281
rect 126428 36246 126480 36252
rect 126520 36304 126572 36310
rect 126520 36246 126572 36252
rect 124218 36207 124220 36216
rect 124272 36207 124274 36216
rect 124220 36178 124272 36184
rect 124036 34468 124088 34474
rect 124036 34410 124088 34416
rect 125508 3188 125560 3194
rect 125508 3130 125560 3136
rect 125416 2848 125468 2854
rect 125416 2790 125468 2796
rect 122840 2644 122892 2650
rect 122840 2586 122892 2592
rect 125428 2446 125456 2790
rect 125520 2446 125548 3130
rect 126992 2650 127020 36518
rect 127094 36476 127402 36485
rect 127094 36474 127100 36476
rect 127156 36474 127180 36476
rect 127236 36474 127260 36476
rect 127316 36474 127340 36476
rect 127396 36474 127402 36476
rect 127156 36422 127158 36474
rect 127338 36422 127340 36474
rect 127094 36420 127100 36422
rect 127156 36420 127180 36422
rect 127236 36420 127260 36422
rect 127316 36420 127340 36422
rect 127396 36420 127402 36422
rect 127094 36411 127402 36420
rect 127094 35388 127402 35397
rect 127094 35386 127100 35388
rect 127156 35386 127180 35388
rect 127236 35386 127260 35388
rect 127316 35386 127340 35388
rect 127396 35386 127402 35388
rect 127156 35334 127158 35386
rect 127338 35334 127340 35386
rect 127094 35332 127100 35334
rect 127156 35332 127180 35334
rect 127236 35332 127260 35334
rect 127316 35332 127340 35334
rect 127396 35332 127402 35334
rect 127094 35323 127402 35332
rect 129292 35057 129320 37062
rect 129568 36786 129596 37198
rect 129660 37108 129688 39200
rect 130580 39114 130608 39200
rect 130672 39114 130700 39222
rect 130580 39086 130700 39114
rect 130292 38140 130344 38146
rect 130292 38082 130344 38088
rect 129740 37120 129792 37126
rect 129660 37080 129740 37108
rect 129740 37062 129792 37068
rect 129556 36780 129608 36786
rect 129556 36722 129608 36728
rect 129568 36689 129596 36722
rect 129554 36680 129610 36689
rect 129554 36615 129610 36624
rect 130304 36582 130332 38082
rect 131040 37244 131068 39222
rect 131486 39200 131542 40000
rect 132406 39200 132462 40000
rect 133326 39200 133382 40000
rect 134246 39200 134302 40000
rect 135166 39200 135222 40000
rect 136086 39200 136142 40000
rect 137006 39200 137062 40000
rect 137926 39200 137982 40000
rect 138846 39200 138902 40000
rect 139766 39200 139822 40000
rect 140686 39200 140742 40000
rect 141606 39200 141662 40000
rect 142526 39200 142582 40000
rect 143446 39200 143502 40000
rect 144366 39200 144422 40000
rect 145286 39200 145342 40000
rect 146206 39200 146262 40000
rect 147126 39200 147182 40000
rect 131120 37256 131172 37262
rect 131040 37216 131120 37244
rect 131120 37198 131172 37204
rect 130476 37120 130528 37126
rect 130476 37062 130528 37068
rect 130292 36576 130344 36582
rect 130292 36518 130344 36524
rect 130488 36038 130516 37062
rect 131132 36922 131160 37198
rect 131500 37126 131528 39200
rect 131672 37256 131724 37262
rect 132420 37244 132448 39200
rect 132500 37256 132552 37262
rect 132420 37216 132500 37244
rect 131672 37198 131724 37204
rect 133236 37256 133288 37262
rect 132500 37198 132552 37204
rect 132866 37224 132922 37233
rect 131488 37120 131540 37126
rect 131488 37062 131540 37068
rect 131120 36916 131172 36922
rect 131120 36858 131172 36864
rect 130936 36780 130988 36786
rect 130936 36722 130988 36728
rect 130948 36582 130976 36722
rect 130936 36576 130988 36582
rect 130936 36518 130988 36524
rect 130948 36038 130976 36518
rect 131684 36281 131712 37198
rect 133236 37198 133288 37204
rect 132866 37159 132922 37168
rect 132880 37126 132908 37159
rect 132868 37120 132920 37126
rect 132868 37062 132920 37068
rect 133248 36922 133276 37198
rect 133340 37126 133368 39200
rect 134260 37262 134288 39200
rect 133512 37256 133564 37262
rect 133512 37198 133564 37204
rect 134248 37256 134300 37262
rect 134248 37198 134300 37204
rect 134432 37256 134484 37262
rect 134432 37198 134484 37204
rect 133328 37120 133380 37126
rect 133328 37062 133380 37068
rect 133236 36916 133288 36922
rect 133236 36858 133288 36864
rect 133524 36854 133552 37198
rect 134260 36922 134288 37198
rect 134248 36916 134300 36922
rect 134248 36858 134300 36864
rect 132132 36848 132184 36854
rect 132132 36790 132184 36796
rect 133512 36848 133564 36854
rect 133512 36790 133564 36796
rect 132040 36780 132092 36786
rect 132040 36722 132092 36728
rect 132052 36310 132080 36722
rect 132144 36310 132172 36790
rect 134444 36718 134472 37198
rect 134524 37120 134576 37126
rect 134524 37062 134576 37068
rect 134432 36712 134484 36718
rect 134432 36654 134484 36660
rect 132040 36304 132092 36310
rect 131670 36272 131726 36281
rect 132040 36246 132092 36252
rect 132132 36304 132184 36310
rect 132132 36246 132184 36252
rect 131670 36207 131726 36216
rect 130476 36032 130528 36038
rect 130476 35974 130528 35980
rect 130936 36032 130988 36038
rect 130936 35974 130988 35980
rect 129278 35048 129334 35057
rect 129278 34983 129334 34992
rect 127094 34300 127402 34309
rect 127094 34298 127100 34300
rect 127156 34298 127180 34300
rect 127236 34298 127260 34300
rect 127316 34298 127340 34300
rect 127396 34298 127402 34300
rect 127156 34246 127158 34298
rect 127338 34246 127340 34298
rect 127094 34244 127100 34246
rect 127156 34244 127180 34246
rect 127236 34244 127260 34246
rect 127316 34244 127340 34246
rect 127396 34244 127402 34246
rect 127094 34235 127402 34244
rect 127094 33212 127402 33221
rect 127094 33210 127100 33212
rect 127156 33210 127180 33212
rect 127236 33210 127260 33212
rect 127316 33210 127340 33212
rect 127396 33210 127402 33212
rect 127156 33158 127158 33210
rect 127338 33158 127340 33210
rect 127094 33156 127100 33158
rect 127156 33156 127180 33158
rect 127236 33156 127260 33158
rect 127316 33156 127340 33158
rect 127396 33156 127402 33158
rect 127094 33147 127402 33156
rect 127094 32124 127402 32133
rect 127094 32122 127100 32124
rect 127156 32122 127180 32124
rect 127236 32122 127260 32124
rect 127316 32122 127340 32124
rect 127396 32122 127402 32124
rect 127156 32070 127158 32122
rect 127338 32070 127340 32122
rect 127094 32068 127100 32070
rect 127156 32068 127180 32070
rect 127236 32068 127260 32070
rect 127316 32068 127340 32070
rect 127396 32068 127402 32070
rect 127094 32059 127402 32068
rect 127094 31036 127402 31045
rect 127094 31034 127100 31036
rect 127156 31034 127180 31036
rect 127236 31034 127260 31036
rect 127316 31034 127340 31036
rect 127396 31034 127402 31036
rect 127156 30982 127158 31034
rect 127338 30982 127340 31034
rect 127094 30980 127100 30982
rect 127156 30980 127180 30982
rect 127236 30980 127260 30982
rect 127316 30980 127340 30982
rect 127396 30980 127402 30982
rect 127094 30971 127402 30980
rect 127094 29948 127402 29957
rect 127094 29946 127100 29948
rect 127156 29946 127180 29948
rect 127236 29946 127260 29948
rect 127316 29946 127340 29948
rect 127396 29946 127402 29948
rect 127156 29894 127158 29946
rect 127338 29894 127340 29946
rect 127094 29892 127100 29894
rect 127156 29892 127180 29894
rect 127236 29892 127260 29894
rect 127316 29892 127340 29894
rect 127396 29892 127402 29894
rect 127094 29883 127402 29892
rect 127094 28860 127402 28869
rect 127094 28858 127100 28860
rect 127156 28858 127180 28860
rect 127236 28858 127260 28860
rect 127316 28858 127340 28860
rect 127396 28858 127402 28860
rect 127156 28806 127158 28858
rect 127338 28806 127340 28858
rect 127094 28804 127100 28806
rect 127156 28804 127180 28806
rect 127236 28804 127260 28806
rect 127316 28804 127340 28806
rect 127396 28804 127402 28806
rect 127094 28795 127402 28804
rect 127094 27772 127402 27781
rect 127094 27770 127100 27772
rect 127156 27770 127180 27772
rect 127236 27770 127260 27772
rect 127316 27770 127340 27772
rect 127396 27770 127402 27772
rect 127156 27718 127158 27770
rect 127338 27718 127340 27770
rect 127094 27716 127100 27718
rect 127156 27716 127180 27718
rect 127236 27716 127260 27718
rect 127316 27716 127340 27718
rect 127396 27716 127402 27718
rect 127094 27707 127402 27716
rect 127094 26684 127402 26693
rect 127094 26682 127100 26684
rect 127156 26682 127180 26684
rect 127236 26682 127260 26684
rect 127316 26682 127340 26684
rect 127396 26682 127402 26684
rect 127156 26630 127158 26682
rect 127338 26630 127340 26682
rect 127094 26628 127100 26630
rect 127156 26628 127180 26630
rect 127236 26628 127260 26630
rect 127316 26628 127340 26630
rect 127396 26628 127402 26630
rect 127094 26619 127402 26628
rect 127094 25596 127402 25605
rect 127094 25594 127100 25596
rect 127156 25594 127180 25596
rect 127236 25594 127260 25596
rect 127316 25594 127340 25596
rect 127396 25594 127402 25596
rect 127156 25542 127158 25594
rect 127338 25542 127340 25594
rect 127094 25540 127100 25542
rect 127156 25540 127180 25542
rect 127236 25540 127260 25542
rect 127316 25540 127340 25542
rect 127396 25540 127402 25542
rect 127094 25531 127402 25540
rect 127094 24508 127402 24517
rect 127094 24506 127100 24508
rect 127156 24506 127180 24508
rect 127236 24506 127260 24508
rect 127316 24506 127340 24508
rect 127396 24506 127402 24508
rect 127156 24454 127158 24506
rect 127338 24454 127340 24506
rect 127094 24452 127100 24454
rect 127156 24452 127180 24454
rect 127236 24452 127260 24454
rect 127316 24452 127340 24454
rect 127396 24452 127402 24454
rect 127094 24443 127402 24452
rect 127094 23420 127402 23429
rect 127094 23418 127100 23420
rect 127156 23418 127180 23420
rect 127236 23418 127260 23420
rect 127316 23418 127340 23420
rect 127396 23418 127402 23420
rect 127156 23366 127158 23418
rect 127338 23366 127340 23418
rect 127094 23364 127100 23366
rect 127156 23364 127180 23366
rect 127236 23364 127260 23366
rect 127316 23364 127340 23366
rect 127396 23364 127402 23366
rect 127094 23355 127402 23364
rect 127094 22332 127402 22341
rect 127094 22330 127100 22332
rect 127156 22330 127180 22332
rect 127236 22330 127260 22332
rect 127316 22330 127340 22332
rect 127396 22330 127402 22332
rect 127156 22278 127158 22330
rect 127338 22278 127340 22330
rect 127094 22276 127100 22278
rect 127156 22276 127180 22278
rect 127236 22276 127260 22278
rect 127316 22276 127340 22278
rect 127396 22276 127402 22278
rect 127094 22267 127402 22276
rect 127094 21244 127402 21253
rect 127094 21242 127100 21244
rect 127156 21242 127180 21244
rect 127236 21242 127260 21244
rect 127316 21242 127340 21244
rect 127396 21242 127402 21244
rect 127156 21190 127158 21242
rect 127338 21190 127340 21242
rect 127094 21188 127100 21190
rect 127156 21188 127180 21190
rect 127236 21188 127260 21190
rect 127316 21188 127340 21190
rect 127396 21188 127402 21190
rect 127094 21179 127402 21188
rect 127094 20156 127402 20165
rect 127094 20154 127100 20156
rect 127156 20154 127180 20156
rect 127236 20154 127260 20156
rect 127316 20154 127340 20156
rect 127396 20154 127402 20156
rect 127156 20102 127158 20154
rect 127338 20102 127340 20154
rect 127094 20100 127100 20102
rect 127156 20100 127180 20102
rect 127236 20100 127260 20102
rect 127316 20100 127340 20102
rect 127396 20100 127402 20102
rect 127094 20091 127402 20100
rect 127094 19068 127402 19077
rect 127094 19066 127100 19068
rect 127156 19066 127180 19068
rect 127236 19066 127260 19068
rect 127316 19066 127340 19068
rect 127396 19066 127402 19068
rect 127156 19014 127158 19066
rect 127338 19014 127340 19066
rect 127094 19012 127100 19014
rect 127156 19012 127180 19014
rect 127236 19012 127260 19014
rect 127316 19012 127340 19014
rect 127396 19012 127402 19014
rect 127094 19003 127402 19012
rect 127094 17980 127402 17989
rect 127094 17978 127100 17980
rect 127156 17978 127180 17980
rect 127236 17978 127260 17980
rect 127316 17978 127340 17980
rect 127396 17978 127402 17980
rect 127156 17926 127158 17978
rect 127338 17926 127340 17978
rect 127094 17924 127100 17926
rect 127156 17924 127180 17926
rect 127236 17924 127260 17926
rect 127316 17924 127340 17926
rect 127396 17924 127402 17926
rect 127094 17915 127402 17924
rect 127094 16892 127402 16901
rect 127094 16890 127100 16892
rect 127156 16890 127180 16892
rect 127236 16890 127260 16892
rect 127316 16890 127340 16892
rect 127396 16890 127402 16892
rect 127156 16838 127158 16890
rect 127338 16838 127340 16890
rect 127094 16836 127100 16838
rect 127156 16836 127180 16838
rect 127236 16836 127260 16838
rect 127316 16836 127340 16838
rect 127396 16836 127402 16838
rect 127094 16827 127402 16836
rect 127094 15804 127402 15813
rect 127094 15802 127100 15804
rect 127156 15802 127180 15804
rect 127236 15802 127260 15804
rect 127316 15802 127340 15804
rect 127396 15802 127402 15804
rect 127156 15750 127158 15802
rect 127338 15750 127340 15802
rect 127094 15748 127100 15750
rect 127156 15748 127180 15750
rect 127236 15748 127260 15750
rect 127316 15748 127340 15750
rect 127396 15748 127402 15750
rect 127094 15739 127402 15748
rect 127094 14716 127402 14725
rect 127094 14714 127100 14716
rect 127156 14714 127180 14716
rect 127236 14714 127260 14716
rect 127316 14714 127340 14716
rect 127396 14714 127402 14716
rect 127156 14662 127158 14714
rect 127338 14662 127340 14714
rect 127094 14660 127100 14662
rect 127156 14660 127180 14662
rect 127236 14660 127260 14662
rect 127316 14660 127340 14662
rect 127396 14660 127402 14662
rect 127094 14651 127402 14660
rect 127094 13628 127402 13637
rect 127094 13626 127100 13628
rect 127156 13626 127180 13628
rect 127236 13626 127260 13628
rect 127316 13626 127340 13628
rect 127396 13626 127402 13628
rect 127156 13574 127158 13626
rect 127338 13574 127340 13626
rect 127094 13572 127100 13574
rect 127156 13572 127180 13574
rect 127236 13572 127260 13574
rect 127316 13572 127340 13574
rect 127396 13572 127402 13574
rect 127094 13563 127402 13572
rect 127094 12540 127402 12549
rect 127094 12538 127100 12540
rect 127156 12538 127180 12540
rect 127236 12538 127260 12540
rect 127316 12538 127340 12540
rect 127396 12538 127402 12540
rect 127156 12486 127158 12538
rect 127338 12486 127340 12538
rect 127094 12484 127100 12486
rect 127156 12484 127180 12486
rect 127236 12484 127260 12486
rect 127316 12484 127340 12486
rect 127396 12484 127402 12486
rect 127094 12475 127402 12484
rect 127094 11452 127402 11461
rect 127094 11450 127100 11452
rect 127156 11450 127180 11452
rect 127236 11450 127260 11452
rect 127316 11450 127340 11452
rect 127396 11450 127402 11452
rect 127156 11398 127158 11450
rect 127338 11398 127340 11450
rect 127094 11396 127100 11398
rect 127156 11396 127180 11398
rect 127236 11396 127260 11398
rect 127316 11396 127340 11398
rect 127396 11396 127402 11398
rect 127094 11387 127402 11396
rect 127094 10364 127402 10373
rect 127094 10362 127100 10364
rect 127156 10362 127180 10364
rect 127236 10362 127260 10364
rect 127316 10362 127340 10364
rect 127396 10362 127402 10364
rect 127156 10310 127158 10362
rect 127338 10310 127340 10362
rect 127094 10308 127100 10310
rect 127156 10308 127180 10310
rect 127236 10308 127260 10310
rect 127316 10308 127340 10310
rect 127396 10308 127402 10310
rect 127094 10299 127402 10308
rect 130948 9602 130976 35974
rect 134536 35193 134564 37062
rect 135180 35894 135208 39200
rect 135996 37256 136048 37262
rect 135996 37198 136048 37204
rect 135536 37120 135588 37126
rect 135536 37062 135588 37068
rect 135548 35894 135576 37062
rect 136008 36922 136036 37198
rect 136100 37194 136128 39200
rect 136088 37188 136140 37194
rect 136088 37130 136140 37136
rect 135996 36916 136048 36922
rect 135996 36858 136048 36864
rect 135904 36712 135956 36718
rect 135904 36654 135956 36660
rect 135916 36378 135944 36654
rect 136100 36378 136128 37130
rect 137020 37126 137048 39200
rect 137940 37244 137968 39200
rect 138020 37256 138072 37262
rect 137940 37216 138020 37244
rect 138020 37198 138072 37204
rect 137008 37120 137060 37126
rect 137008 37062 137060 37068
rect 137284 36848 137336 36854
rect 137284 36790 137336 36796
rect 135904 36372 135956 36378
rect 135904 36314 135956 36320
rect 136088 36372 136140 36378
rect 136088 36314 136140 36320
rect 137296 36310 137324 36790
rect 137652 36780 137704 36786
rect 137652 36722 137704 36728
rect 137284 36304 137336 36310
rect 137284 36246 137336 36252
rect 137664 36038 137692 36722
rect 138032 36378 138060 37198
rect 138860 37126 138888 39200
rect 139780 37262 139808 39200
rect 138940 37256 138992 37262
rect 138940 37198 138992 37204
rect 139768 37256 139820 37262
rect 139768 37198 139820 37204
rect 140504 37256 140556 37262
rect 140504 37198 140556 37204
rect 140700 37210 140728 39200
rect 141620 37262 141648 39200
rect 141608 37256 141660 37262
rect 138848 37120 138900 37126
rect 138848 37062 138900 37068
rect 138952 36922 138980 37198
rect 139492 37120 139544 37126
rect 139492 37062 139544 37068
rect 138940 36916 138992 36922
rect 138940 36858 138992 36864
rect 139504 36582 139532 37062
rect 140516 36922 140544 37198
rect 140700 37182 140820 37210
rect 141608 37198 141660 37204
rect 142252 37256 142304 37262
rect 142252 37198 142304 37204
rect 140792 37126 140820 37182
rect 142160 37188 142212 37194
rect 142160 37130 142212 37136
rect 140688 37120 140740 37126
rect 140688 37062 140740 37068
rect 140780 37120 140832 37126
rect 140780 37062 140832 37068
rect 140504 36916 140556 36922
rect 140504 36858 140556 36864
rect 139492 36576 139544 36582
rect 139492 36518 139544 36524
rect 138020 36372 138072 36378
rect 138020 36314 138072 36320
rect 139504 36242 139532 36518
rect 139492 36236 139544 36242
rect 139492 36178 139544 36184
rect 137652 36032 137704 36038
rect 137652 35974 137704 35980
rect 135180 35866 135576 35894
rect 134522 35184 134578 35193
rect 134522 35119 134578 35128
rect 130948 9574 131160 9602
rect 127094 9276 127402 9285
rect 127094 9274 127100 9276
rect 127156 9274 127180 9276
rect 127236 9274 127260 9276
rect 127316 9274 127340 9276
rect 127396 9274 127402 9276
rect 127156 9222 127158 9274
rect 127338 9222 127340 9274
rect 127094 9220 127100 9222
rect 127156 9220 127180 9222
rect 127236 9220 127260 9222
rect 127316 9220 127340 9222
rect 127396 9220 127402 9222
rect 127094 9211 127402 9220
rect 127094 8188 127402 8197
rect 127094 8186 127100 8188
rect 127156 8186 127180 8188
rect 127236 8186 127260 8188
rect 127316 8186 127340 8188
rect 127396 8186 127402 8188
rect 127156 8134 127158 8186
rect 127338 8134 127340 8186
rect 127094 8132 127100 8134
rect 127156 8132 127180 8134
rect 127236 8132 127260 8134
rect 127316 8132 127340 8134
rect 127396 8132 127402 8134
rect 127094 8123 127402 8132
rect 127094 7100 127402 7109
rect 127094 7098 127100 7100
rect 127156 7098 127180 7100
rect 127236 7098 127260 7100
rect 127316 7098 127340 7100
rect 127396 7098 127402 7100
rect 127156 7046 127158 7098
rect 127338 7046 127340 7098
rect 127094 7044 127100 7046
rect 127156 7044 127180 7046
rect 127236 7044 127260 7046
rect 127316 7044 127340 7046
rect 127396 7044 127402 7046
rect 127094 7035 127402 7044
rect 127094 6012 127402 6021
rect 127094 6010 127100 6012
rect 127156 6010 127180 6012
rect 127236 6010 127260 6012
rect 127316 6010 127340 6012
rect 127396 6010 127402 6012
rect 127156 5958 127158 6010
rect 127338 5958 127340 6010
rect 127094 5956 127100 5958
rect 127156 5956 127180 5958
rect 127236 5956 127260 5958
rect 127316 5956 127340 5958
rect 127396 5956 127402 5958
rect 127094 5947 127402 5956
rect 127094 4924 127402 4933
rect 127094 4922 127100 4924
rect 127156 4922 127180 4924
rect 127236 4922 127260 4924
rect 127316 4922 127340 4924
rect 127396 4922 127402 4924
rect 127156 4870 127158 4922
rect 127338 4870 127340 4922
rect 127094 4868 127100 4870
rect 127156 4868 127180 4870
rect 127236 4868 127260 4870
rect 127316 4868 127340 4870
rect 127396 4868 127402 4870
rect 127094 4859 127402 4868
rect 127094 3836 127402 3845
rect 127094 3834 127100 3836
rect 127156 3834 127180 3836
rect 127236 3834 127260 3836
rect 127316 3834 127340 3836
rect 127396 3834 127402 3836
rect 127156 3782 127158 3834
rect 127338 3782 127340 3834
rect 127094 3780 127100 3782
rect 127156 3780 127180 3782
rect 127236 3780 127260 3782
rect 127316 3780 127340 3782
rect 127396 3780 127402 3782
rect 127094 3771 127402 3780
rect 130844 2848 130896 2854
rect 130844 2790 130896 2796
rect 127094 2748 127402 2757
rect 127094 2746 127100 2748
rect 127156 2746 127180 2748
rect 127236 2746 127260 2748
rect 127316 2746 127340 2748
rect 127396 2746 127402 2748
rect 127156 2694 127158 2746
rect 127338 2694 127340 2746
rect 127094 2692 127100 2694
rect 127156 2692 127180 2694
rect 127236 2692 127260 2694
rect 127316 2692 127340 2694
rect 127396 2692 127402 2694
rect 127094 2683 127402 2692
rect 126980 2644 127032 2650
rect 126980 2586 127032 2592
rect 125416 2440 125468 2446
rect 125416 2382 125468 2388
rect 125508 2440 125560 2446
rect 125508 2382 125560 2388
rect 110420 2372 110472 2378
rect 110420 2314 110472 2320
rect 118424 2372 118476 2378
rect 118424 2314 118476 2320
rect 122564 2372 122616 2378
rect 122564 2314 122616 2320
rect 109040 2304 109092 2310
rect 109040 2246 109092 2252
rect 109052 1766 109080 2246
rect 109040 1760 109092 1766
rect 110432 1714 110460 2314
rect 112444 2304 112496 2310
rect 112444 2246 112496 2252
rect 112904 2304 112956 2310
rect 112904 2246 112956 2252
rect 114284 2304 114336 2310
rect 114284 2246 114336 2252
rect 116676 2304 116728 2310
rect 116676 2246 116728 2252
rect 117044 2304 117096 2310
rect 117044 2246 117096 2252
rect 111734 2204 112042 2213
rect 111734 2202 111740 2204
rect 111796 2202 111820 2204
rect 111876 2202 111900 2204
rect 111956 2202 111980 2204
rect 112036 2202 112042 2204
rect 111796 2150 111798 2202
rect 111978 2150 111980 2202
rect 111734 2148 111740 2150
rect 111796 2148 111820 2150
rect 111876 2148 111900 2150
rect 111956 2148 111980 2150
rect 112036 2148 112042 2150
rect 111734 2139 112042 2148
rect 109040 1702 109092 1708
rect 110156 1686 110460 1714
rect 110156 800 110184 1686
rect 112456 1494 112484 2246
rect 112444 1488 112496 1494
rect 112444 1430 112496 1436
rect 112916 800 112944 2246
rect 114296 800 114324 2246
rect 116688 1834 116716 2246
rect 116676 1828 116728 1834
rect 116676 1770 116728 1776
rect 117056 800 117084 2246
rect 118436 800 118464 2314
rect 121184 2304 121236 2310
rect 121184 2246 121236 2252
rect 121196 800 121224 2246
rect 122576 800 122604 2314
rect 125324 2304 125376 2310
rect 125324 2246 125376 2252
rect 125336 800 125364 2246
rect 125428 1562 125456 2382
rect 130856 2378 130884 2790
rect 131132 2650 131160 9574
rect 137284 3120 137336 3126
rect 137284 3062 137336 3068
rect 137296 2650 137324 3062
rect 131120 2644 131172 2650
rect 131120 2586 131172 2592
rect 137284 2644 137336 2650
rect 137284 2586 137336 2592
rect 137296 2446 137324 2586
rect 139504 2582 139532 36178
rect 140700 35290 140728 37062
rect 142172 36854 142200 37130
rect 142264 36854 142292 37198
rect 142540 37126 142568 39200
rect 143080 37256 143132 37262
rect 143080 37198 143132 37204
rect 143460 37210 143488 39200
rect 143540 37256 143592 37262
rect 143460 37204 143540 37210
rect 143460 37198 143592 37204
rect 142528 37120 142580 37126
rect 142528 37062 142580 37068
rect 142454 37020 142762 37029
rect 142454 37018 142460 37020
rect 142516 37018 142540 37020
rect 142596 37018 142620 37020
rect 142676 37018 142700 37020
rect 142756 37018 142762 37020
rect 142516 36966 142518 37018
rect 142698 36966 142700 37018
rect 142454 36964 142460 36966
rect 142516 36964 142540 36966
rect 142596 36964 142620 36966
rect 142676 36964 142700 36966
rect 142756 36964 142762 36966
rect 142454 36955 142762 36964
rect 143092 36922 143120 37198
rect 143460 37182 143580 37198
rect 143080 36916 143132 36922
rect 143080 36858 143132 36864
rect 142160 36848 142212 36854
rect 142160 36790 142212 36796
rect 142252 36848 142304 36854
rect 142252 36790 142304 36796
rect 141332 36712 141384 36718
rect 141332 36654 141384 36660
rect 140688 35284 140740 35290
rect 140688 35226 140740 35232
rect 141344 2650 141372 36654
rect 143552 36378 143580 37182
rect 144380 37126 144408 39200
rect 145300 37262 145328 39200
rect 144552 37256 144604 37262
rect 144552 37198 144604 37204
rect 145288 37256 145340 37262
rect 145288 37198 145340 37204
rect 144000 37120 144052 37126
rect 144000 37062 144052 37068
rect 144368 37120 144420 37126
rect 144368 37062 144420 37068
rect 143632 36780 143684 36786
rect 143632 36722 143684 36728
rect 143540 36372 143592 36378
rect 143540 36314 143592 36320
rect 143644 36174 143672 36722
rect 143632 36168 143684 36174
rect 143632 36110 143684 36116
rect 142454 35932 142762 35941
rect 142454 35930 142460 35932
rect 142516 35930 142540 35932
rect 142596 35930 142620 35932
rect 142676 35930 142700 35932
rect 142756 35930 142762 35932
rect 142516 35878 142518 35930
rect 142698 35878 142700 35930
rect 142454 35876 142460 35878
rect 142516 35876 142540 35878
rect 142596 35876 142620 35878
rect 142676 35876 142700 35878
rect 142756 35876 142762 35878
rect 142454 35867 142762 35876
rect 142454 34844 142762 34853
rect 142454 34842 142460 34844
rect 142516 34842 142540 34844
rect 142596 34842 142620 34844
rect 142676 34842 142700 34844
rect 142756 34842 142762 34844
rect 142516 34790 142518 34842
rect 142698 34790 142700 34842
rect 142454 34788 142460 34790
rect 142516 34788 142540 34790
rect 142596 34788 142620 34790
rect 142676 34788 142700 34790
rect 142756 34788 142762 34790
rect 142454 34779 142762 34788
rect 142454 33756 142762 33765
rect 142454 33754 142460 33756
rect 142516 33754 142540 33756
rect 142596 33754 142620 33756
rect 142676 33754 142700 33756
rect 142756 33754 142762 33756
rect 142516 33702 142518 33754
rect 142698 33702 142700 33754
rect 142454 33700 142460 33702
rect 142516 33700 142540 33702
rect 142596 33700 142620 33702
rect 142676 33700 142700 33702
rect 142756 33700 142762 33702
rect 142454 33691 142762 33700
rect 142454 32668 142762 32677
rect 142454 32666 142460 32668
rect 142516 32666 142540 32668
rect 142596 32666 142620 32668
rect 142676 32666 142700 32668
rect 142756 32666 142762 32668
rect 142516 32614 142518 32666
rect 142698 32614 142700 32666
rect 142454 32612 142460 32614
rect 142516 32612 142540 32614
rect 142596 32612 142620 32614
rect 142676 32612 142700 32614
rect 142756 32612 142762 32614
rect 142454 32603 142762 32612
rect 142454 31580 142762 31589
rect 142454 31578 142460 31580
rect 142516 31578 142540 31580
rect 142596 31578 142620 31580
rect 142676 31578 142700 31580
rect 142756 31578 142762 31580
rect 142516 31526 142518 31578
rect 142698 31526 142700 31578
rect 142454 31524 142460 31526
rect 142516 31524 142540 31526
rect 142596 31524 142620 31526
rect 142676 31524 142700 31526
rect 142756 31524 142762 31526
rect 142454 31515 142762 31524
rect 142454 30492 142762 30501
rect 142454 30490 142460 30492
rect 142516 30490 142540 30492
rect 142596 30490 142620 30492
rect 142676 30490 142700 30492
rect 142756 30490 142762 30492
rect 142516 30438 142518 30490
rect 142698 30438 142700 30490
rect 142454 30436 142460 30438
rect 142516 30436 142540 30438
rect 142596 30436 142620 30438
rect 142676 30436 142700 30438
rect 142756 30436 142762 30438
rect 142454 30427 142762 30436
rect 142454 29404 142762 29413
rect 142454 29402 142460 29404
rect 142516 29402 142540 29404
rect 142596 29402 142620 29404
rect 142676 29402 142700 29404
rect 142756 29402 142762 29404
rect 142516 29350 142518 29402
rect 142698 29350 142700 29402
rect 142454 29348 142460 29350
rect 142516 29348 142540 29350
rect 142596 29348 142620 29350
rect 142676 29348 142700 29350
rect 142756 29348 142762 29350
rect 142454 29339 142762 29348
rect 142454 28316 142762 28325
rect 142454 28314 142460 28316
rect 142516 28314 142540 28316
rect 142596 28314 142620 28316
rect 142676 28314 142700 28316
rect 142756 28314 142762 28316
rect 142516 28262 142518 28314
rect 142698 28262 142700 28314
rect 142454 28260 142460 28262
rect 142516 28260 142540 28262
rect 142596 28260 142620 28262
rect 142676 28260 142700 28262
rect 142756 28260 142762 28262
rect 142454 28251 142762 28260
rect 142454 27228 142762 27237
rect 142454 27226 142460 27228
rect 142516 27226 142540 27228
rect 142596 27226 142620 27228
rect 142676 27226 142700 27228
rect 142756 27226 142762 27228
rect 142516 27174 142518 27226
rect 142698 27174 142700 27226
rect 142454 27172 142460 27174
rect 142516 27172 142540 27174
rect 142596 27172 142620 27174
rect 142676 27172 142700 27174
rect 142756 27172 142762 27174
rect 142454 27163 142762 27172
rect 143644 26234 143672 36110
rect 144012 34406 144040 37062
rect 144564 36922 144592 37198
rect 145300 36922 145328 37198
rect 146220 37126 146248 39200
rect 147140 37262 147168 39200
rect 146300 37256 146352 37262
rect 146300 37198 146352 37204
rect 147128 37256 147180 37262
rect 147128 37198 147180 37204
rect 146208 37120 146260 37126
rect 146208 37062 146260 37068
rect 146312 36922 146340 37198
rect 147140 36922 147168 37198
rect 147404 37120 147456 37126
rect 147404 37062 147456 37068
rect 144552 36916 144604 36922
rect 144552 36858 144604 36864
rect 145288 36916 145340 36922
rect 145288 36858 145340 36864
rect 146300 36916 146352 36922
rect 146300 36858 146352 36864
rect 147128 36916 147180 36922
rect 147128 36858 147180 36864
rect 146300 36780 146352 36786
rect 146300 36722 146352 36728
rect 146312 36106 146340 36722
rect 146300 36100 146352 36106
rect 146300 36042 146352 36048
rect 147312 36100 147364 36106
rect 147312 36042 147364 36048
rect 144000 34400 144052 34406
rect 144000 34342 144052 34348
rect 143552 26206 143672 26234
rect 142454 26140 142762 26149
rect 142454 26138 142460 26140
rect 142516 26138 142540 26140
rect 142596 26138 142620 26140
rect 142676 26138 142700 26140
rect 142756 26138 142762 26140
rect 142516 26086 142518 26138
rect 142698 26086 142700 26138
rect 142454 26084 142460 26086
rect 142516 26084 142540 26086
rect 142596 26084 142620 26086
rect 142676 26084 142700 26086
rect 142756 26084 142762 26086
rect 142454 26075 142762 26084
rect 142454 25052 142762 25061
rect 142454 25050 142460 25052
rect 142516 25050 142540 25052
rect 142596 25050 142620 25052
rect 142676 25050 142700 25052
rect 142756 25050 142762 25052
rect 142516 24998 142518 25050
rect 142698 24998 142700 25050
rect 142454 24996 142460 24998
rect 142516 24996 142540 24998
rect 142596 24996 142620 24998
rect 142676 24996 142700 24998
rect 142756 24996 142762 24998
rect 142454 24987 142762 24996
rect 142454 23964 142762 23973
rect 142454 23962 142460 23964
rect 142516 23962 142540 23964
rect 142596 23962 142620 23964
rect 142676 23962 142700 23964
rect 142756 23962 142762 23964
rect 142516 23910 142518 23962
rect 142698 23910 142700 23962
rect 142454 23908 142460 23910
rect 142516 23908 142540 23910
rect 142596 23908 142620 23910
rect 142676 23908 142700 23910
rect 142756 23908 142762 23910
rect 142454 23899 142762 23908
rect 142454 22876 142762 22885
rect 142454 22874 142460 22876
rect 142516 22874 142540 22876
rect 142596 22874 142620 22876
rect 142676 22874 142700 22876
rect 142756 22874 142762 22876
rect 142516 22822 142518 22874
rect 142698 22822 142700 22874
rect 142454 22820 142460 22822
rect 142516 22820 142540 22822
rect 142596 22820 142620 22822
rect 142676 22820 142700 22822
rect 142756 22820 142762 22822
rect 142454 22811 142762 22820
rect 142454 21788 142762 21797
rect 142454 21786 142460 21788
rect 142516 21786 142540 21788
rect 142596 21786 142620 21788
rect 142676 21786 142700 21788
rect 142756 21786 142762 21788
rect 142516 21734 142518 21786
rect 142698 21734 142700 21786
rect 142454 21732 142460 21734
rect 142516 21732 142540 21734
rect 142596 21732 142620 21734
rect 142676 21732 142700 21734
rect 142756 21732 142762 21734
rect 142454 21723 142762 21732
rect 142454 20700 142762 20709
rect 142454 20698 142460 20700
rect 142516 20698 142540 20700
rect 142596 20698 142620 20700
rect 142676 20698 142700 20700
rect 142756 20698 142762 20700
rect 142516 20646 142518 20698
rect 142698 20646 142700 20698
rect 142454 20644 142460 20646
rect 142516 20644 142540 20646
rect 142596 20644 142620 20646
rect 142676 20644 142700 20646
rect 142756 20644 142762 20646
rect 142454 20635 142762 20644
rect 142454 19612 142762 19621
rect 142454 19610 142460 19612
rect 142516 19610 142540 19612
rect 142596 19610 142620 19612
rect 142676 19610 142700 19612
rect 142756 19610 142762 19612
rect 142516 19558 142518 19610
rect 142698 19558 142700 19610
rect 142454 19556 142460 19558
rect 142516 19556 142540 19558
rect 142596 19556 142620 19558
rect 142676 19556 142700 19558
rect 142756 19556 142762 19558
rect 142454 19547 142762 19556
rect 142454 18524 142762 18533
rect 142454 18522 142460 18524
rect 142516 18522 142540 18524
rect 142596 18522 142620 18524
rect 142676 18522 142700 18524
rect 142756 18522 142762 18524
rect 142516 18470 142518 18522
rect 142698 18470 142700 18522
rect 142454 18468 142460 18470
rect 142516 18468 142540 18470
rect 142596 18468 142620 18470
rect 142676 18468 142700 18470
rect 142756 18468 142762 18470
rect 142454 18459 142762 18468
rect 142454 17436 142762 17445
rect 142454 17434 142460 17436
rect 142516 17434 142540 17436
rect 142596 17434 142620 17436
rect 142676 17434 142700 17436
rect 142756 17434 142762 17436
rect 142516 17382 142518 17434
rect 142698 17382 142700 17434
rect 142454 17380 142460 17382
rect 142516 17380 142540 17382
rect 142596 17380 142620 17382
rect 142676 17380 142700 17382
rect 142756 17380 142762 17382
rect 142454 17371 142762 17380
rect 142454 16348 142762 16357
rect 142454 16346 142460 16348
rect 142516 16346 142540 16348
rect 142596 16346 142620 16348
rect 142676 16346 142700 16348
rect 142756 16346 142762 16348
rect 142516 16294 142518 16346
rect 142698 16294 142700 16346
rect 142454 16292 142460 16294
rect 142516 16292 142540 16294
rect 142596 16292 142620 16294
rect 142676 16292 142700 16294
rect 142756 16292 142762 16294
rect 142454 16283 142762 16292
rect 142454 15260 142762 15269
rect 142454 15258 142460 15260
rect 142516 15258 142540 15260
rect 142596 15258 142620 15260
rect 142676 15258 142700 15260
rect 142756 15258 142762 15260
rect 142516 15206 142518 15258
rect 142698 15206 142700 15258
rect 142454 15204 142460 15206
rect 142516 15204 142540 15206
rect 142596 15204 142620 15206
rect 142676 15204 142700 15206
rect 142756 15204 142762 15206
rect 142454 15195 142762 15204
rect 142454 14172 142762 14181
rect 142454 14170 142460 14172
rect 142516 14170 142540 14172
rect 142596 14170 142620 14172
rect 142676 14170 142700 14172
rect 142756 14170 142762 14172
rect 142516 14118 142518 14170
rect 142698 14118 142700 14170
rect 142454 14116 142460 14118
rect 142516 14116 142540 14118
rect 142596 14116 142620 14118
rect 142676 14116 142700 14118
rect 142756 14116 142762 14118
rect 142454 14107 142762 14116
rect 142454 13084 142762 13093
rect 142454 13082 142460 13084
rect 142516 13082 142540 13084
rect 142596 13082 142620 13084
rect 142676 13082 142700 13084
rect 142756 13082 142762 13084
rect 142516 13030 142518 13082
rect 142698 13030 142700 13082
rect 142454 13028 142460 13030
rect 142516 13028 142540 13030
rect 142596 13028 142620 13030
rect 142676 13028 142700 13030
rect 142756 13028 142762 13030
rect 142454 13019 142762 13028
rect 142454 11996 142762 12005
rect 142454 11994 142460 11996
rect 142516 11994 142540 11996
rect 142596 11994 142620 11996
rect 142676 11994 142700 11996
rect 142756 11994 142762 11996
rect 142516 11942 142518 11994
rect 142698 11942 142700 11994
rect 142454 11940 142460 11942
rect 142516 11940 142540 11942
rect 142596 11940 142620 11942
rect 142676 11940 142700 11942
rect 142756 11940 142762 11942
rect 142454 11931 142762 11940
rect 142454 10908 142762 10917
rect 142454 10906 142460 10908
rect 142516 10906 142540 10908
rect 142596 10906 142620 10908
rect 142676 10906 142700 10908
rect 142756 10906 142762 10908
rect 142516 10854 142518 10906
rect 142698 10854 142700 10906
rect 142454 10852 142460 10854
rect 142516 10852 142540 10854
rect 142596 10852 142620 10854
rect 142676 10852 142700 10854
rect 142756 10852 142762 10854
rect 142454 10843 142762 10852
rect 142454 9820 142762 9829
rect 142454 9818 142460 9820
rect 142516 9818 142540 9820
rect 142596 9818 142620 9820
rect 142676 9818 142700 9820
rect 142756 9818 142762 9820
rect 142516 9766 142518 9818
rect 142698 9766 142700 9818
rect 142454 9764 142460 9766
rect 142516 9764 142540 9766
rect 142596 9764 142620 9766
rect 142676 9764 142700 9766
rect 142756 9764 142762 9766
rect 142454 9755 142762 9764
rect 142454 8732 142762 8741
rect 142454 8730 142460 8732
rect 142516 8730 142540 8732
rect 142596 8730 142620 8732
rect 142676 8730 142700 8732
rect 142756 8730 142762 8732
rect 142516 8678 142518 8730
rect 142698 8678 142700 8730
rect 142454 8676 142460 8678
rect 142516 8676 142540 8678
rect 142596 8676 142620 8678
rect 142676 8676 142700 8678
rect 142756 8676 142762 8678
rect 142454 8667 142762 8676
rect 142454 7644 142762 7653
rect 142454 7642 142460 7644
rect 142516 7642 142540 7644
rect 142596 7642 142620 7644
rect 142676 7642 142700 7644
rect 142756 7642 142762 7644
rect 142516 7590 142518 7642
rect 142698 7590 142700 7642
rect 142454 7588 142460 7590
rect 142516 7588 142540 7590
rect 142596 7588 142620 7590
rect 142676 7588 142700 7590
rect 142756 7588 142762 7590
rect 142454 7579 142762 7588
rect 142454 6556 142762 6565
rect 142454 6554 142460 6556
rect 142516 6554 142540 6556
rect 142596 6554 142620 6556
rect 142676 6554 142700 6556
rect 142756 6554 142762 6556
rect 142516 6502 142518 6554
rect 142698 6502 142700 6554
rect 142454 6500 142460 6502
rect 142516 6500 142540 6502
rect 142596 6500 142620 6502
rect 142676 6500 142700 6502
rect 142756 6500 142762 6502
rect 142454 6491 142762 6500
rect 142454 5468 142762 5477
rect 142454 5466 142460 5468
rect 142516 5466 142540 5468
rect 142596 5466 142620 5468
rect 142676 5466 142700 5468
rect 142756 5466 142762 5468
rect 142516 5414 142518 5466
rect 142698 5414 142700 5466
rect 142454 5412 142460 5414
rect 142516 5412 142540 5414
rect 142596 5412 142620 5414
rect 142676 5412 142700 5414
rect 142756 5412 142762 5414
rect 142454 5403 142762 5412
rect 142454 4380 142762 4389
rect 142454 4378 142460 4380
rect 142516 4378 142540 4380
rect 142596 4378 142620 4380
rect 142676 4378 142700 4380
rect 142756 4378 142762 4380
rect 142516 4326 142518 4378
rect 142698 4326 142700 4378
rect 142454 4324 142460 4326
rect 142516 4324 142540 4326
rect 142596 4324 142620 4326
rect 142676 4324 142700 4326
rect 142756 4324 142762 4326
rect 142454 4315 142762 4324
rect 142454 3292 142762 3301
rect 142454 3290 142460 3292
rect 142516 3290 142540 3292
rect 142596 3290 142620 3292
rect 142676 3290 142700 3292
rect 142756 3290 142762 3292
rect 142516 3238 142518 3290
rect 142698 3238 142700 3290
rect 142454 3236 142460 3238
rect 142516 3236 142540 3238
rect 142596 3236 142620 3238
rect 142676 3236 142700 3238
rect 142756 3236 142762 3238
rect 142454 3227 142762 3236
rect 143264 2848 143316 2854
rect 143264 2790 143316 2796
rect 141332 2644 141384 2650
rect 141332 2586 141384 2592
rect 139492 2576 139544 2582
rect 139492 2518 139544 2524
rect 137284 2440 137336 2446
rect 137284 2382 137336 2388
rect 139124 2440 139176 2446
rect 139124 2382 139176 2388
rect 126704 2372 126756 2378
rect 126704 2314 126756 2320
rect 130844 2372 130896 2378
rect 130844 2314 130896 2320
rect 125416 1556 125468 1562
rect 125416 1498 125468 1504
rect 126716 800 126744 2314
rect 129648 2304 129700 2310
rect 129648 2246 129700 2252
rect 129660 1170 129688 2246
rect 129476 1142 129688 1170
rect 129476 800 129504 1142
rect 130856 800 130884 2314
rect 133604 2304 133656 2310
rect 133604 2246 133656 2252
rect 134984 2304 135036 2310
rect 134984 2246 135036 2252
rect 137744 2304 137796 2310
rect 137744 2246 137796 2252
rect 133616 800 133644 2246
rect 134996 800 135024 2246
rect 137756 800 137784 2246
rect 139136 800 139164 2382
rect 143276 2378 143304 2790
rect 143552 2650 143580 26206
rect 145932 3732 145984 3738
rect 145932 3674 145984 3680
rect 145944 3194 145972 3674
rect 145932 3188 145984 3194
rect 145932 3130 145984 3136
rect 143540 2644 143592 2650
rect 143540 2586 143592 2592
rect 145944 2446 145972 3130
rect 147324 2650 147352 36042
rect 147416 33114 147444 37062
rect 147404 33108 147456 33114
rect 147404 33050 147456 33056
rect 147312 2644 147364 2650
rect 147312 2586 147364 2592
rect 145932 2440 145984 2446
rect 145932 2382 145984 2388
rect 143264 2372 143316 2378
rect 143264 2314 143316 2320
rect 147404 2372 147456 2378
rect 147404 2314 147456 2320
rect 141424 2304 141476 2310
rect 141424 2246 141476 2252
rect 141884 2304 141936 2310
rect 141884 2246 141936 2252
rect 141436 1698 141464 2246
rect 141424 1692 141476 1698
rect 141424 1634 141476 1640
rect 141896 800 141924 2246
rect 142454 2204 142762 2213
rect 142454 2202 142460 2204
rect 142516 2202 142540 2204
rect 142596 2202 142620 2204
rect 142676 2202 142700 2204
rect 142756 2202 142762 2204
rect 142516 2150 142518 2202
rect 142698 2150 142700 2202
rect 142454 2148 142460 2150
rect 142516 2148 142540 2150
rect 142596 2148 142620 2150
rect 142676 2148 142700 2150
rect 142756 2148 142762 2150
rect 142454 2139 142762 2148
rect 143276 800 143304 2314
rect 146024 2304 146076 2310
rect 146024 2246 146076 2252
rect 146036 800 146064 2246
rect 147416 800 147444 2314
rect 2502 0 2558 800
rect 3882 0 3938 800
rect 5262 0 5318 800
rect 6642 0 6698 800
rect 8022 0 8078 800
rect 9402 0 9458 800
rect 10782 0 10838 800
rect 12162 0 12218 800
rect 13542 0 13598 800
rect 14922 0 14978 800
rect 16302 0 16358 800
rect 17682 0 17738 800
rect 19062 0 19118 800
rect 20442 0 20498 800
rect 21822 0 21878 800
rect 23202 0 23258 800
rect 24582 0 24638 800
rect 25962 0 26018 800
rect 27342 0 27398 800
rect 28722 0 28778 800
rect 30102 0 30158 800
rect 31482 0 31538 800
rect 32862 0 32918 800
rect 34242 0 34298 800
rect 35622 0 35678 800
rect 37002 0 37058 800
rect 38382 0 38438 800
rect 39762 0 39818 800
rect 41142 0 41198 800
rect 42522 0 42578 800
rect 43902 0 43958 800
rect 45282 0 45338 800
rect 46662 0 46718 800
rect 48042 0 48098 800
rect 49422 0 49478 800
rect 50802 0 50858 800
rect 52182 0 52238 800
rect 53562 0 53618 800
rect 54942 0 54998 800
rect 56322 0 56378 800
rect 57702 0 57758 800
rect 59082 0 59138 800
rect 60462 0 60518 800
rect 61842 0 61898 800
rect 63222 0 63278 800
rect 64602 0 64658 800
rect 65982 0 66038 800
rect 67362 0 67418 800
rect 68742 0 68798 800
rect 70122 0 70178 800
rect 71502 0 71558 800
rect 72882 0 72938 800
rect 74262 0 74318 800
rect 75642 0 75698 800
rect 77022 0 77078 800
rect 78402 0 78458 800
rect 79782 0 79838 800
rect 81162 0 81218 800
rect 82542 0 82598 800
rect 83922 0 83978 800
rect 85302 0 85358 800
rect 86682 0 86738 800
rect 88062 0 88118 800
rect 89442 0 89498 800
rect 90822 0 90878 800
rect 92202 0 92258 800
rect 93582 0 93638 800
rect 94962 0 95018 800
rect 96342 0 96398 800
rect 97722 0 97778 800
rect 99102 0 99158 800
rect 100482 0 100538 800
rect 101862 0 101918 800
rect 103242 0 103298 800
rect 104622 0 104678 800
rect 106002 0 106058 800
rect 107382 0 107438 800
rect 108762 0 108818 800
rect 110142 0 110198 800
rect 111522 0 111578 800
rect 112902 0 112958 800
rect 114282 0 114338 800
rect 115662 0 115718 800
rect 117042 0 117098 800
rect 118422 0 118478 800
rect 119802 0 119858 800
rect 121182 0 121238 800
rect 122562 0 122618 800
rect 123942 0 123998 800
rect 125322 0 125378 800
rect 126702 0 126758 800
rect 128082 0 128138 800
rect 129462 0 129518 800
rect 130842 0 130898 800
rect 132222 0 132278 800
rect 133602 0 133658 800
rect 134982 0 135038 800
rect 136362 0 136418 800
rect 137742 0 137798 800
rect 139122 0 139178 800
rect 140502 0 140558 800
rect 141882 0 141938 800
rect 143262 0 143318 800
rect 144642 0 144698 800
rect 146022 0 146078 800
rect 147402 0 147458 800
<< via2 >>
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 12898 36644 12954 36680
rect 12898 36624 12900 36644
rect 12900 36624 12952 36644
rect 12952 36624 12954 36644
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 16578 36760 16634 36816
rect 15106 36100 15162 36136
rect 15106 36080 15108 36100
rect 15108 36080 15160 36100
rect 15160 36080 15162 36100
rect 19706 37204 19708 37224
rect 19708 37204 19760 37224
rect 19760 37204 19762 37224
rect 19706 37168 19762 37204
rect 19982 37168 20038 37224
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 20442 37440 20498 37496
rect 20258 36524 20260 36544
rect 20260 36524 20312 36544
rect 20312 36524 20314 36544
rect 20258 36488 20314 36524
rect 20810 36524 20812 36544
rect 20812 36524 20864 36544
rect 20864 36524 20866 36544
rect 20810 36488 20866 36524
rect 21270 36216 21326 36272
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 22282 37204 22284 37224
rect 22284 37204 22336 37224
rect 22336 37204 22338 37224
rect 22282 37168 22338 37204
rect 23294 37032 23350 37088
rect 22742 36624 22798 36680
rect 23386 36624 23442 36680
rect 24490 36896 24546 36952
rect 22006 3596 22062 3632
rect 22006 3576 22008 3596
rect 22008 3576 22060 3596
rect 22060 3576 22062 3596
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 24858 37168 24914 37224
rect 28170 37440 28226 37496
rect 28998 37304 29054 37360
rect 28078 3596 28134 3632
rect 28078 3576 28080 3596
rect 28080 3576 28132 3596
rect 28132 3576 28134 3596
rect 30562 36760 30618 36816
rect 30010 35672 30066 35728
rect 31758 33904 31814 33960
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34426 36236 34482 36272
rect 34426 36216 34428 36236
rect 34428 36216 34480 36236
rect 34480 36216 34482 36236
rect 34702 35128 34758 35184
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 35714 37032 35770 37088
rect 36634 37068 36636 37088
rect 36636 37068 36688 37088
rect 36688 37068 36690 37088
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 36450 36760 36506 36816
rect 36634 37032 36690 37068
rect 36818 37304 36874 37360
rect 37094 36780 37150 36816
rect 37094 36760 37096 36780
rect 37096 36760 37148 36780
rect 37148 36760 37150 36780
rect 37186 34448 37242 34504
rect 38566 36488 38622 36544
rect 39946 36352 40002 36408
rect 40314 37168 40370 37224
rect 41050 36644 41106 36680
rect 41050 36624 41052 36644
rect 41052 36624 41104 36644
rect 41104 36624 41106 36644
rect 41050 36100 41106 36136
rect 41050 36080 41052 36100
rect 41052 36080 41104 36100
rect 41104 36080 41106 36100
rect 41234 36080 41290 36136
rect 41142 35572 41144 35592
rect 41144 35572 41196 35592
rect 41196 35572 41198 35592
rect 41142 35536 41198 35572
rect 41418 35572 41420 35592
rect 41420 35572 41472 35592
rect 41472 35572 41474 35592
rect 41418 35536 41474 35572
rect 41326 33496 41382 33552
rect 41694 36080 41750 36136
rect 43074 36760 43130 36816
rect 42890 36216 42946 36272
rect 43350 35028 43352 35048
rect 43352 35028 43404 35048
rect 43404 35028 43406 35048
rect 43350 34992 43406 35028
rect 41970 34040 42026 34096
rect 41694 2916 41750 2952
rect 41694 2896 41696 2916
rect 41696 2896 41748 2916
rect 41748 2896 41750 2916
rect 42614 2896 42670 2952
rect 43718 36352 43774 36408
rect 43810 36216 43866 36272
rect 44178 36624 44234 36680
rect 44178 36352 44234 36408
rect 44546 35028 44548 35048
rect 44548 35028 44600 35048
rect 44600 35028 44602 35048
rect 44546 34992 44602 35028
rect 45282 35980 45284 36000
rect 45284 35980 45336 36000
rect 45336 35980 45338 36000
rect 45282 35944 45338 35980
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50710 35980 50712 36000
rect 50712 35980 50764 36000
rect 50764 35980 50766 36000
rect 50710 35944 50766 35980
rect 50894 35536 50950 35592
rect 51262 36624 51318 36680
rect 51446 35128 51502 35184
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 53010 37168 53066 37224
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 53010 36352 53066 36408
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 53746 35808 53802 35864
rect 55678 37188 55734 37224
rect 55678 37168 55680 37188
rect 55680 37168 55732 37188
rect 55732 37168 55734 37188
rect 56138 35944 56194 36000
rect 57150 36624 57206 36680
rect 58346 37440 58402 37496
rect 58254 37324 58310 37360
rect 58254 37304 58256 37324
rect 58256 37304 58308 37324
rect 58308 37304 58310 37324
rect 58346 37204 58348 37224
rect 58348 37204 58400 37224
rect 58400 37204 58402 37224
rect 58346 37168 58402 37204
rect 58622 37324 58678 37360
rect 58622 37304 58624 37324
rect 58624 37304 58676 37324
rect 58676 37304 58678 37324
rect 59818 37440 59874 37496
rect 61382 37324 61438 37360
rect 61382 37304 61384 37324
rect 61384 37304 61436 37324
rect 61436 37304 61438 37324
rect 61750 35944 61806 36000
rect 64786 37204 64788 37224
rect 64788 37204 64840 37224
rect 64840 37204 64842 37224
rect 64786 37168 64842 37204
rect 64970 37168 65026 37224
rect 65660 37562 65716 37564
rect 65740 37562 65796 37564
rect 65820 37562 65876 37564
rect 65900 37562 65956 37564
rect 65660 37510 65706 37562
rect 65706 37510 65716 37562
rect 65740 37510 65770 37562
rect 65770 37510 65782 37562
rect 65782 37510 65796 37562
rect 65820 37510 65834 37562
rect 65834 37510 65846 37562
rect 65846 37510 65876 37562
rect 65900 37510 65910 37562
rect 65910 37510 65956 37562
rect 65660 37508 65716 37510
rect 65740 37508 65796 37510
rect 65820 37508 65876 37510
rect 65900 37508 65956 37510
rect 65798 37168 65854 37224
rect 65246 35028 65248 35048
rect 65248 35028 65300 35048
rect 65300 35028 65302 35048
rect 65246 34992 65302 35028
rect 65660 36474 65716 36476
rect 65740 36474 65796 36476
rect 65820 36474 65876 36476
rect 65900 36474 65956 36476
rect 65660 36422 65706 36474
rect 65706 36422 65716 36474
rect 65740 36422 65770 36474
rect 65770 36422 65782 36474
rect 65782 36422 65796 36474
rect 65820 36422 65834 36474
rect 65834 36422 65846 36474
rect 65846 36422 65876 36474
rect 65900 36422 65910 36474
rect 65910 36422 65956 36474
rect 65660 36420 65716 36422
rect 65740 36420 65796 36422
rect 65820 36420 65876 36422
rect 65900 36420 65956 36422
rect 65660 35386 65716 35388
rect 65740 35386 65796 35388
rect 65820 35386 65876 35388
rect 65900 35386 65956 35388
rect 65660 35334 65706 35386
rect 65706 35334 65716 35386
rect 65740 35334 65770 35386
rect 65770 35334 65782 35386
rect 65782 35334 65796 35386
rect 65820 35334 65834 35386
rect 65834 35334 65846 35386
rect 65846 35334 65876 35386
rect 65900 35334 65910 35386
rect 65910 35334 65956 35386
rect 65660 35332 65716 35334
rect 65740 35332 65796 35334
rect 65820 35332 65876 35334
rect 65900 35332 65956 35334
rect 65660 34298 65716 34300
rect 65740 34298 65796 34300
rect 65820 34298 65876 34300
rect 65900 34298 65956 34300
rect 65660 34246 65706 34298
rect 65706 34246 65716 34298
rect 65740 34246 65770 34298
rect 65770 34246 65782 34298
rect 65782 34246 65796 34298
rect 65820 34246 65834 34298
rect 65834 34246 65846 34298
rect 65846 34246 65876 34298
rect 65900 34246 65910 34298
rect 65910 34246 65956 34298
rect 65660 34244 65716 34246
rect 65740 34244 65796 34246
rect 65820 34244 65876 34246
rect 65900 34244 65956 34246
rect 65660 33210 65716 33212
rect 65740 33210 65796 33212
rect 65820 33210 65876 33212
rect 65900 33210 65956 33212
rect 65660 33158 65706 33210
rect 65706 33158 65716 33210
rect 65740 33158 65770 33210
rect 65770 33158 65782 33210
rect 65782 33158 65796 33210
rect 65820 33158 65834 33210
rect 65834 33158 65846 33210
rect 65846 33158 65876 33210
rect 65900 33158 65910 33210
rect 65910 33158 65956 33210
rect 65660 33156 65716 33158
rect 65740 33156 65796 33158
rect 65820 33156 65876 33158
rect 65900 33156 65956 33158
rect 65660 32122 65716 32124
rect 65740 32122 65796 32124
rect 65820 32122 65876 32124
rect 65900 32122 65956 32124
rect 65660 32070 65706 32122
rect 65706 32070 65716 32122
rect 65740 32070 65770 32122
rect 65770 32070 65782 32122
rect 65782 32070 65796 32122
rect 65820 32070 65834 32122
rect 65834 32070 65846 32122
rect 65846 32070 65876 32122
rect 65900 32070 65910 32122
rect 65910 32070 65956 32122
rect 65660 32068 65716 32070
rect 65740 32068 65796 32070
rect 65820 32068 65876 32070
rect 65900 32068 65956 32070
rect 66442 35980 66444 36000
rect 66444 35980 66496 36000
rect 66496 35980 66498 36000
rect 66442 35944 66498 35980
rect 65660 31034 65716 31036
rect 65740 31034 65796 31036
rect 65820 31034 65876 31036
rect 65900 31034 65956 31036
rect 65660 30982 65706 31034
rect 65706 30982 65716 31034
rect 65740 30982 65770 31034
rect 65770 30982 65782 31034
rect 65782 30982 65796 31034
rect 65820 30982 65834 31034
rect 65834 30982 65846 31034
rect 65846 30982 65876 31034
rect 65900 30982 65910 31034
rect 65910 30982 65956 31034
rect 65660 30980 65716 30982
rect 65740 30980 65796 30982
rect 65820 30980 65876 30982
rect 65900 30980 65956 30982
rect 65660 29946 65716 29948
rect 65740 29946 65796 29948
rect 65820 29946 65876 29948
rect 65900 29946 65956 29948
rect 65660 29894 65706 29946
rect 65706 29894 65716 29946
rect 65740 29894 65770 29946
rect 65770 29894 65782 29946
rect 65782 29894 65796 29946
rect 65820 29894 65834 29946
rect 65834 29894 65846 29946
rect 65846 29894 65876 29946
rect 65900 29894 65910 29946
rect 65910 29894 65956 29946
rect 65660 29892 65716 29894
rect 65740 29892 65796 29894
rect 65820 29892 65876 29894
rect 65900 29892 65956 29894
rect 65660 28858 65716 28860
rect 65740 28858 65796 28860
rect 65820 28858 65876 28860
rect 65900 28858 65956 28860
rect 65660 28806 65706 28858
rect 65706 28806 65716 28858
rect 65740 28806 65770 28858
rect 65770 28806 65782 28858
rect 65782 28806 65796 28858
rect 65820 28806 65834 28858
rect 65834 28806 65846 28858
rect 65846 28806 65876 28858
rect 65900 28806 65910 28858
rect 65910 28806 65956 28858
rect 65660 28804 65716 28806
rect 65740 28804 65796 28806
rect 65820 28804 65876 28806
rect 65900 28804 65956 28806
rect 65660 27770 65716 27772
rect 65740 27770 65796 27772
rect 65820 27770 65876 27772
rect 65900 27770 65956 27772
rect 65660 27718 65706 27770
rect 65706 27718 65716 27770
rect 65740 27718 65770 27770
rect 65770 27718 65782 27770
rect 65782 27718 65796 27770
rect 65820 27718 65834 27770
rect 65834 27718 65846 27770
rect 65846 27718 65876 27770
rect 65900 27718 65910 27770
rect 65910 27718 65956 27770
rect 65660 27716 65716 27718
rect 65740 27716 65796 27718
rect 65820 27716 65876 27718
rect 65900 27716 65956 27718
rect 65660 26682 65716 26684
rect 65740 26682 65796 26684
rect 65820 26682 65876 26684
rect 65900 26682 65956 26684
rect 65660 26630 65706 26682
rect 65706 26630 65716 26682
rect 65740 26630 65770 26682
rect 65770 26630 65782 26682
rect 65782 26630 65796 26682
rect 65820 26630 65834 26682
rect 65834 26630 65846 26682
rect 65846 26630 65876 26682
rect 65900 26630 65910 26682
rect 65910 26630 65956 26682
rect 65660 26628 65716 26630
rect 65740 26628 65796 26630
rect 65820 26628 65876 26630
rect 65900 26628 65956 26630
rect 65660 25594 65716 25596
rect 65740 25594 65796 25596
rect 65820 25594 65876 25596
rect 65900 25594 65956 25596
rect 65660 25542 65706 25594
rect 65706 25542 65716 25594
rect 65740 25542 65770 25594
rect 65770 25542 65782 25594
rect 65782 25542 65796 25594
rect 65820 25542 65834 25594
rect 65834 25542 65846 25594
rect 65846 25542 65876 25594
rect 65900 25542 65910 25594
rect 65910 25542 65956 25594
rect 65660 25540 65716 25542
rect 65740 25540 65796 25542
rect 65820 25540 65876 25542
rect 65900 25540 65956 25542
rect 65660 24506 65716 24508
rect 65740 24506 65796 24508
rect 65820 24506 65876 24508
rect 65900 24506 65956 24508
rect 65660 24454 65706 24506
rect 65706 24454 65716 24506
rect 65740 24454 65770 24506
rect 65770 24454 65782 24506
rect 65782 24454 65796 24506
rect 65820 24454 65834 24506
rect 65834 24454 65846 24506
rect 65846 24454 65876 24506
rect 65900 24454 65910 24506
rect 65910 24454 65956 24506
rect 65660 24452 65716 24454
rect 65740 24452 65796 24454
rect 65820 24452 65876 24454
rect 65900 24452 65956 24454
rect 65660 23418 65716 23420
rect 65740 23418 65796 23420
rect 65820 23418 65876 23420
rect 65900 23418 65956 23420
rect 65660 23366 65706 23418
rect 65706 23366 65716 23418
rect 65740 23366 65770 23418
rect 65770 23366 65782 23418
rect 65782 23366 65796 23418
rect 65820 23366 65834 23418
rect 65834 23366 65846 23418
rect 65846 23366 65876 23418
rect 65900 23366 65910 23418
rect 65910 23366 65956 23418
rect 65660 23364 65716 23366
rect 65740 23364 65796 23366
rect 65820 23364 65876 23366
rect 65900 23364 65956 23366
rect 65660 22330 65716 22332
rect 65740 22330 65796 22332
rect 65820 22330 65876 22332
rect 65900 22330 65956 22332
rect 65660 22278 65706 22330
rect 65706 22278 65716 22330
rect 65740 22278 65770 22330
rect 65770 22278 65782 22330
rect 65782 22278 65796 22330
rect 65820 22278 65834 22330
rect 65834 22278 65846 22330
rect 65846 22278 65876 22330
rect 65900 22278 65910 22330
rect 65910 22278 65956 22330
rect 65660 22276 65716 22278
rect 65740 22276 65796 22278
rect 65820 22276 65876 22278
rect 65900 22276 65956 22278
rect 65660 21242 65716 21244
rect 65740 21242 65796 21244
rect 65820 21242 65876 21244
rect 65900 21242 65956 21244
rect 65660 21190 65706 21242
rect 65706 21190 65716 21242
rect 65740 21190 65770 21242
rect 65770 21190 65782 21242
rect 65782 21190 65796 21242
rect 65820 21190 65834 21242
rect 65834 21190 65846 21242
rect 65846 21190 65876 21242
rect 65900 21190 65910 21242
rect 65910 21190 65956 21242
rect 65660 21188 65716 21190
rect 65740 21188 65796 21190
rect 65820 21188 65876 21190
rect 65900 21188 65956 21190
rect 65660 20154 65716 20156
rect 65740 20154 65796 20156
rect 65820 20154 65876 20156
rect 65900 20154 65956 20156
rect 65660 20102 65706 20154
rect 65706 20102 65716 20154
rect 65740 20102 65770 20154
rect 65770 20102 65782 20154
rect 65782 20102 65796 20154
rect 65820 20102 65834 20154
rect 65834 20102 65846 20154
rect 65846 20102 65876 20154
rect 65900 20102 65910 20154
rect 65910 20102 65956 20154
rect 65660 20100 65716 20102
rect 65740 20100 65796 20102
rect 65820 20100 65876 20102
rect 65900 20100 65956 20102
rect 65660 19066 65716 19068
rect 65740 19066 65796 19068
rect 65820 19066 65876 19068
rect 65900 19066 65956 19068
rect 65660 19014 65706 19066
rect 65706 19014 65716 19066
rect 65740 19014 65770 19066
rect 65770 19014 65782 19066
rect 65782 19014 65796 19066
rect 65820 19014 65834 19066
rect 65834 19014 65846 19066
rect 65846 19014 65876 19066
rect 65900 19014 65910 19066
rect 65910 19014 65956 19066
rect 65660 19012 65716 19014
rect 65740 19012 65796 19014
rect 65820 19012 65876 19014
rect 65900 19012 65956 19014
rect 65660 17978 65716 17980
rect 65740 17978 65796 17980
rect 65820 17978 65876 17980
rect 65900 17978 65956 17980
rect 65660 17926 65706 17978
rect 65706 17926 65716 17978
rect 65740 17926 65770 17978
rect 65770 17926 65782 17978
rect 65782 17926 65796 17978
rect 65820 17926 65834 17978
rect 65834 17926 65846 17978
rect 65846 17926 65876 17978
rect 65900 17926 65910 17978
rect 65910 17926 65956 17978
rect 65660 17924 65716 17926
rect 65740 17924 65796 17926
rect 65820 17924 65876 17926
rect 65900 17924 65956 17926
rect 65660 16890 65716 16892
rect 65740 16890 65796 16892
rect 65820 16890 65876 16892
rect 65900 16890 65956 16892
rect 65660 16838 65706 16890
rect 65706 16838 65716 16890
rect 65740 16838 65770 16890
rect 65770 16838 65782 16890
rect 65782 16838 65796 16890
rect 65820 16838 65834 16890
rect 65834 16838 65846 16890
rect 65846 16838 65876 16890
rect 65900 16838 65910 16890
rect 65910 16838 65956 16890
rect 65660 16836 65716 16838
rect 65740 16836 65796 16838
rect 65820 16836 65876 16838
rect 65900 16836 65956 16838
rect 65660 15802 65716 15804
rect 65740 15802 65796 15804
rect 65820 15802 65876 15804
rect 65900 15802 65956 15804
rect 65660 15750 65706 15802
rect 65706 15750 65716 15802
rect 65740 15750 65770 15802
rect 65770 15750 65782 15802
rect 65782 15750 65796 15802
rect 65820 15750 65834 15802
rect 65834 15750 65846 15802
rect 65846 15750 65876 15802
rect 65900 15750 65910 15802
rect 65910 15750 65956 15802
rect 65660 15748 65716 15750
rect 65740 15748 65796 15750
rect 65820 15748 65876 15750
rect 65900 15748 65956 15750
rect 65660 14714 65716 14716
rect 65740 14714 65796 14716
rect 65820 14714 65876 14716
rect 65900 14714 65956 14716
rect 65660 14662 65706 14714
rect 65706 14662 65716 14714
rect 65740 14662 65770 14714
rect 65770 14662 65782 14714
rect 65782 14662 65796 14714
rect 65820 14662 65834 14714
rect 65834 14662 65846 14714
rect 65846 14662 65876 14714
rect 65900 14662 65910 14714
rect 65910 14662 65956 14714
rect 65660 14660 65716 14662
rect 65740 14660 65796 14662
rect 65820 14660 65876 14662
rect 65900 14660 65956 14662
rect 65660 13626 65716 13628
rect 65740 13626 65796 13628
rect 65820 13626 65876 13628
rect 65900 13626 65956 13628
rect 65660 13574 65706 13626
rect 65706 13574 65716 13626
rect 65740 13574 65770 13626
rect 65770 13574 65782 13626
rect 65782 13574 65796 13626
rect 65820 13574 65834 13626
rect 65834 13574 65846 13626
rect 65846 13574 65876 13626
rect 65900 13574 65910 13626
rect 65910 13574 65956 13626
rect 65660 13572 65716 13574
rect 65740 13572 65796 13574
rect 65820 13572 65876 13574
rect 65900 13572 65956 13574
rect 65660 12538 65716 12540
rect 65740 12538 65796 12540
rect 65820 12538 65876 12540
rect 65900 12538 65956 12540
rect 65660 12486 65706 12538
rect 65706 12486 65716 12538
rect 65740 12486 65770 12538
rect 65770 12486 65782 12538
rect 65782 12486 65796 12538
rect 65820 12486 65834 12538
rect 65834 12486 65846 12538
rect 65846 12486 65876 12538
rect 65900 12486 65910 12538
rect 65910 12486 65956 12538
rect 65660 12484 65716 12486
rect 65740 12484 65796 12486
rect 65820 12484 65876 12486
rect 65900 12484 65956 12486
rect 65660 11450 65716 11452
rect 65740 11450 65796 11452
rect 65820 11450 65876 11452
rect 65900 11450 65956 11452
rect 65660 11398 65706 11450
rect 65706 11398 65716 11450
rect 65740 11398 65770 11450
rect 65770 11398 65782 11450
rect 65782 11398 65796 11450
rect 65820 11398 65834 11450
rect 65834 11398 65846 11450
rect 65846 11398 65876 11450
rect 65900 11398 65910 11450
rect 65910 11398 65956 11450
rect 65660 11396 65716 11398
rect 65740 11396 65796 11398
rect 65820 11396 65876 11398
rect 65900 11396 65956 11398
rect 65660 10362 65716 10364
rect 65740 10362 65796 10364
rect 65820 10362 65876 10364
rect 65900 10362 65956 10364
rect 65660 10310 65706 10362
rect 65706 10310 65716 10362
rect 65740 10310 65770 10362
rect 65770 10310 65782 10362
rect 65782 10310 65796 10362
rect 65820 10310 65834 10362
rect 65834 10310 65846 10362
rect 65846 10310 65876 10362
rect 65900 10310 65910 10362
rect 65910 10310 65956 10362
rect 65660 10308 65716 10310
rect 65740 10308 65796 10310
rect 65820 10308 65876 10310
rect 65900 10308 65956 10310
rect 65660 9274 65716 9276
rect 65740 9274 65796 9276
rect 65820 9274 65876 9276
rect 65900 9274 65956 9276
rect 65660 9222 65706 9274
rect 65706 9222 65716 9274
rect 65740 9222 65770 9274
rect 65770 9222 65782 9274
rect 65782 9222 65796 9274
rect 65820 9222 65834 9274
rect 65834 9222 65846 9274
rect 65846 9222 65876 9274
rect 65900 9222 65910 9274
rect 65910 9222 65956 9274
rect 65660 9220 65716 9222
rect 65740 9220 65796 9222
rect 65820 9220 65876 9222
rect 65900 9220 65956 9222
rect 65660 8186 65716 8188
rect 65740 8186 65796 8188
rect 65820 8186 65876 8188
rect 65900 8186 65956 8188
rect 65660 8134 65706 8186
rect 65706 8134 65716 8186
rect 65740 8134 65770 8186
rect 65770 8134 65782 8186
rect 65782 8134 65796 8186
rect 65820 8134 65834 8186
rect 65834 8134 65846 8186
rect 65846 8134 65876 8186
rect 65900 8134 65910 8186
rect 65910 8134 65956 8186
rect 65660 8132 65716 8134
rect 65740 8132 65796 8134
rect 65820 8132 65876 8134
rect 65900 8132 65956 8134
rect 65660 7098 65716 7100
rect 65740 7098 65796 7100
rect 65820 7098 65876 7100
rect 65900 7098 65956 7100
rect 65660 7046 65706 7098
rect 65706 7046 65716 7098
rect 65740 7046 65770 7098
rect 65770 7046 65782 7098
rect 65782 7046 65796 7098
rect 65820 7046 65834 7098
rect 65834 7046 65846 7098
rect 65846 7046 65876 7098
rect 65900 7046 65910 7098
rect 65910 7046 65956 7098
rect 65660 7044 65716 7046
rect 65740 7044 65796 7046
rect 65820 7044 65876 7046
rect 65900 7044 65956 7046
rect 65660 6010 65716 6012
rect 65740 6010 65796 6012
rect 65820 6010 65876 6012
rect 65900 6010 65956 6012
rect 65660 5958 65706 6010
rect 65706 5958 65716 6010
rect 65740 5958 65770 6010
rect 65770 5958 65782 6010
rect 65782 5958 65796 6010
rect 65820 5958 65834 6010
rect 65834 5958 65846 6010
rect 65846 5958 65876 6010
rect 65900 5958 65910 6010
rect 65910 5958 65956 6010
rect 65660 5956 65716 5958
rect 65740 5956 65796 5958
rect 65820 5956 65876 5958
rect 65900 5956 65956 5958
rect 68558 37188 68614 37224
rect 68558 37168 68560 37188
rect 68560 37168 68612 37188
rect 68612 37168 68614 37188
rect 68190 35944 68246 36000
rect 65660 4922 65716 4924
rect 65740 4922 65796 4924
rect 65820 4922 65876 4924
rect 65900 4922 65956 4924
rect 65660 4870 65706 4922
rect 65706 4870 65716 4922
rect 65740 4870 65770 4922
rect 65770 4870 65782 4922
rect 65782 4870 65796 4922
rect 65820 4870 65834 4922
rect 65834 4870 65846 4922
rect 65846 4870 65876 4922
rect 65900 4870 65910 4922
rect 65910 4870 65956 4922
rect 65660 4868 65716 4870
rect 65740 4868 65796 4870
rect 65820 4868 65876 4870
rect 65900 4868 65956 4870
rect 65660 3834 65716 3836
rect 65740 3834 65796 3836
rect 65820 3834 65876 3836
rect 65900 3834 65956 3836
rect 65660 3782 65706 3834
rect 65706 3782 65716 3834
rect 65740 3782 65770 3834
rect 65770 3782 65782 3834
rect 65782 3782 65796 3834
rect 65820 3782 65834 3834
rect 65834 3782 65846 3834
rect 65846 3782 65876 3834
rect 65900 3782 65910 3834
rect 65910 3782 65956 3834
rect 65660 3780 65716 3782
rect 65740 3780 65796 3782
rect 65820 3780 65876 3782
rect 65900 3780 65956 3782
rect 65660 2746 65716 2748
rect 65740 2746 65796 2748
rect 65820 2746 65876 2748
rect 65900 2746 65956 2748
rect 65660 2694 65706 2746
rect 65706 2694 65716 2746
rect 65740 2694 65770 2746
rect 65770 2694 65782 2746
rect 65782 2694 65796 2746
rect 65820 2694 65834 2746
rect 65834 2694 65846 2746
rect 65846 2694 65876 2746
rect 65900 2694 65910 2746
rect 65910 2694 65956 2746
rect 65660 2692 65716 2694
rect 65740 2692 65796 2694
rect 65820 2692 65876 2694
rect 65900 2692 65956 2694
rect 68466 3476 68468 3496
rect 68468 3476 68520 3496
rect 68520 3476 68522 3496
rect 68466 3440 68522 3476
rect 73158 37304 73214 37360
rect 71686 35128 71742 35184
rect 74906 36896 74962 36952
rect 74998 36760 75054 36816
rect 74998 36488 75054 36544
rect 74906 36352 74962 36408
rect 75458 36896 75514 36952
rect 69938 2932 69940 2952
rect 69940 2932 69992 2952
rect 69992 2932 69994 2952
rect 69938 2896 69994 2932
rect 71226 3440 71282 3496
rect 76654 36896 76710 36952
rect 79046 37440 79102 37496
rect 79506 37576 79562 37632
rect 76562 35944 76618 36000
rect 77298 35808 77354 35864
rect 75734 2896 75790 2952
rect 79966 36896 80022 36952
rect 80426 37440 80482 37496
rect 80334 36916 80390 36952
rect 80334 36896 80336 36916
rect 80336 36896 80388 36916
rect 80388 36896 80390 36916
rect 81020 37018 81076 37020
rect 81100 37018 81156 37020
rect 81180 37018 81236 37020
rect 81260 37018 81316 37020
rect 81020 36966 81066 37018
rect 81066 36966 81076 37018
rect 81100 36966 81130 37018
rect 81130 36966 81142 37018
rect 81142 36966 81156 37018
rect 81180 36966 81194 37018
rect 81194 36966 81206 37018
rect 81206 36966 81236 37018
rect 81260 36966 81270 37018
rect 81270 36966 81316 37018
rect 81020 36964 81076 36966
rect 81100 36964 81156 36966
rect 81180 36964 81236 36966
rect 81260 36964 81316 36966
rect 81020 35930 81076 35932
rect 81100 35930 81156 35932
rect 81180 35930 81236 35932
rect 81260 35930 81316 35932
rect 81020 35878 81066 35930
rect 81066 35878 81076 35930
rect 81100 35878 81130 35930
rect 81130 35878 81142 35930
rect 81142 35878 81156 35930
rect 81180 35878 81194 35930
rect 81194 35878 81206 35930
rect 81206 35878 81236 35930
rect 81260 35878 81270 35930
rect 81270 35878 81316 35930
rect 81020 35876 81076 35878
rect 81100 35876 81156 35878
rect 81180 35876 81236 35878
rect 81260 35876 81316 35878
rect 80426 35692 80482 35728
rect 80426 35672 80428 35692
rect 80428 35672 80480 35692
rect 80480 35672 80482 35692
rect 81020 34842 81076 34844
rect 81100 34842 81156 34844
rect 81180 34842 81236 34844
rect 81260 34842 81316 34844
rect 81020 34790 81066 34842
rect 81066 34790 81076 34842
rect 81100 34790 81130 34842
rect 81130 34790 81142 34842
rect 81142 34790 81156 34842
rect 81180 34790 81194 34842
rect 81194 34790 81206 34842
rect 81206 34790 81236 34842
rect 81260 34790 81270 34842
rect 81270 34790 81316 34842
rect 81020 34788 81076 34790
rect 81100 34788 81156 34790
rect 81180 34788 81236 34790
rect 81260 34788 81316 34790
rect 81020 33754 81076 33756
rect 81100 33754 81156 33756
rect 81180 33754 81236 33756
rect 81260 33754 81316 33756
rect 81020 33702 81066 33754
rect 81066 33702 81076 33754
rect 81100 33702 81130 33754
rect 81130 33702 81142 33754
rect 81142 33702 81156 33754
rect 81180 33702 81194 33754
rect 81194 33702 81206 33754
rect 81206 33702 81236 33754
rect 81260 33702 81270 33754
rect 81270 33702 81316 33754
rect 81020 33700 81076 33702
rect 81100 33700 81156 33702
rect 81180 33700 81236 33702
rect 81260 33700 81316 33702
rect 81020 32666 81076 32668
rect 81100 32666 81156 32668
rect 81180 32666 81236 32668
rect 81260 32666 81316 32668
rect 81020 32614 81066 32666
rect 81066 32614 81076 32666
rect 81100 32614 81130 32666
rect 81130 32614 81142 32666
rect 81142 32614 81156 32666
rect 81180 32614 81194 32666
rect 81194 32614 81206 32666
rect 81206 32614 81236 32666
rect 81260 32614 81270 32666
rect 81270 32614 81316 32666
rect 81020 32612 81076 32614
rect 81100 32612 81156 32614
rect 81180 32612 81236 32614
rect 81260 32612 81316 32614
rect 81020 31578 81076 31580
rect 81100 31578 81156 31580
rect 81180 31578 81236 31580
rect 81260 31578 81316 31580
rect 81020 31526 81066 31578
rect 81066 31526 81076 31578
rect 81100 31526 81130 31578
rect 81130 31526 81142 31578
rect 81142 31526 81156 31578
rect 81180 31526 81194 31578
rect 81194 31526 81206 31578
rect 81206 31526 81236 31578
rect 81260 31526 81270 31578
rect 81270 31526 81316 31578
rect 81020 31524 81076 31526
rect 81100 31524 81156 31526
rect 81180 31524 81236 31526
rect 81260 31524 81316 31526
rect 81020 30490 81076 30492
rect 81100 30490 81156 30492
rect 81180 30490 81236 30492
rect 81260 30490 81316 30492
rect 81020 30438 81066 30490
rect 81066 30438 81076 30490
rect 81100 30438 81130 30490
rect 81130 30438 81142 30490
rect 81142 30438 81156 30490
rect 81180 30438 81194 30490
rect 81194 30438 81206 30490
rect 81206 30438 81236 30490
rect 81260 30438 81270 30490
rect 81270 30438 81316 30490
rect 81020 30436 81076 30438
rect 81100 30436 81156 30438
rect 81180 30436 81236 30438
rect 81260 30436 81316 30438
rect 81020 29402 81076 29404
rect 81100 29402 81156 29404
rect 81180 29402 81236 29404
rect 81260 29402 81316 29404
rect 81020 29350 81066 29402
rect 81066 29350 81076 29402
rect 81100 29350 81130 29402
rect 81130 29350 81142 29402
rect 81142 29350 81156 29402
rect 81180 29350 81194 29402
rect 81194 29350 81206 29402
rect 81206 29350 81236 29402
rect 81260 29350 81270 29402
rect 81270 29350 81316 29402
rect 81020 29348 81076 29350
rect 81100 29348 81156 29350
rect 81180 29348 81236 29350
rect 81260 29348 81316 29350
rect 81020 28314 81076 28316
rect 81100 28314 81156 28316
rect 81180 28314 81236 28316
rect 81260 28314 81316 28316
rect 81020 28262 81066 28314
rect 81066 28262 81076 28314
rect 81100 28262 81130 28314
rect 81130 28262 81142 28314
rect 81142 28262 81156 28314
rect 81180 28262 81194 28314
rect 81194 28262 81206 28314
rect 81206 28262 81236 28314
rect 81260 28262 81270 28314
rect 81270 28262 81316 28314
rect 81020 28260 81076 28262
rect 81100 28260 81156 28262
rect 81180 28260 81236 28262
rect 81260 28260 81316 28262
rect 81020 27226 81076 27228
rect 81100 27226 81156 27228
rect 81180 27226 81236 27228
rect 81260 27226 81316 27228
rect 81020 27174 81066 27226
rect 81066 27174 81076 27226
rect 81100 27174 81130 27226
rect 81130 27174 81142 27226
rect 81142 27174 81156 27226
rect 81180 27174 81194 27226
rect 81194 27174 81206 27226
rect 81206 27174 81236 27226
rect 81260 27174 81270 27226
rect 81270 27174 81316 27226
rect 81020 27172 81076 27174
rect 81100 27172 81156 27174
rect 81180 27172 81236 27174
rect 81260 27172 81316 27174
rect 82818 37304 82874 37360
rect 81020 26138 81076 26140
rect 81100 26138 81156 26140
rect 81180 26138 81236 26140
rect 81260 26138 81316 26140
rect 81020 26086 81066 26138
rect 81066 26086 81076 26138
rect 81100 26086 81130 26138
rect 81130 26086 81142 26138
rect 81142 26086 81156 26138
rect 81180 26086 81194 26138
rect 81194 26086 81206 26138
rect 81206 26086 81236 26138
rect 81260 26086 81270 26138
rect 81270 26086 81316 26138
rect 81020 26084 81076 26086
rect 81100 26084 81156 26086
rect 81180 26084 81236 26086
rect 81260 26084 81316 26086
rect 81020 25050 81076 25052
rect 81100 25050 81156 25052
rect 81180 25050 81236 25052
rect 81260 25050 81316 25052
rect 81020 24998 81066 25050
rect 81066 24998 81076 25050
rect 81100 24998 81130 25050
rect 81130 24998 81142 25050
rect 81142 24998 81156 25050
rect 81180 24998 81194 25050
rect 81194 24998 81206 25050
rect 81206 24998 81236 25050
rect 81260 24998 81270 25050
rect 81270 24998 81316 25050
rect 81020 24996 81076 24998
rect 81100 24996 81156 24998
rect 81180 24996 81236 24998
rect 81260 24996 81316 24998
rect 81020 23962 81076 23964
rect 81100 23962 81156 23964
rect 81180 23962 81236 23964
rect 81260 23962 81316 23964
rect 81020 23910 81066 23962
rect 81066 23910 81076 23962
rect 81100 23910 81130 23962
rect 81130 23910 81142 23962
rect 81142 23910 81156 23962
rect 81180 23910 81194 23962
rect 81194 23910 81206 23962
rect 81206 23910 81236 23962
rect 81260 23910 81270 23962
rect 81270 23910 81316 23962
rect 81020 23908 81076 23910
rect 81100 23908 81156 23910
rect 81180 23908 81236 23910
rect 81260 23908 81316 23910
rect 81020 22874 81076 22876
rect 81100 22874 81156 22876
rect 81180 22874 81236 22876
rect 81260 22874 81316 22876
rect 81020 22822 81066 22874
rect 81066 22822 81076 22874
rect 81100 22822 81130 22874
rect 81130 22822 81142 22874
rect 81142 22822 81156 22874
rect 81180 22822 81194 22874
rect 81194 22822 81206 22874
rect 81206 22822 81236 22874
rect 81260 22822 81270 22874
rect 81270 22822 81316 22874
rect 81020 22820 81076 22822
rect 81100 22820 81156 22822
rect 81180 22820 81236 22822
rect 81260 22820 81316 22822
rect 81020 21786 81076 21788
rect 81100 21786 81156 21788
rect 81180 21786 81236 21788
rect 81260 21786 81316 21788
rect 81020 21734 81066 21786
rect 81066 21734 81076 21786
rect 81100 21734 81130 21786
rect 81130 21734 81142 21786
rect 81142 21734 81156 21786
rect 81180 21734 81194 21786
rect 81194 21734 81206 21786
rect 81206 21734 81236 21786
rect 81260 21734 81270 21786
rect 81270 21734 81316 21786
rect 81020 21732 81076 21734
rect 81100 21732 81156 21734
rect 81180 21732 81236 21734
rect 81260 21732 81316 21734
rect 81020 20698 81076 20700
rect 81100 20698 81156 20700
rect 81180 20698 81236 20700
rect 81260 20698 81316 20700
rect 81020 20646 81066 20698
rect 81066 20646 81076 20698
rect 81100 20646 81130 20698
rect 81130 20646 81142 20698
rect 81142 20646 81156 20698
rect 81180 20646 81194 20698
rect 81194 20646 81206 20698
rect 81206 20646 81236 20698
rect 81260 20646 81270 20698
rect 81270 20646 81316 20698
rect 81020 20644 81076 20646
rect 81100 20644 81156 20646
rect 81180 20644 81236 20646
rect 81260 20644 81316 20646
rect 81020 19610 81076 19612
rect 81100 19610 81156 19612
rect 81180 19610 81236 19612
rect 81260 19610 81316 19612
rect 81020 19558 81066 19610
rect 81066 19558 81076 19610
rect 81100 19558 81130 19610
rect 81130 19558 81142 19610
rect 81142 19558 81156 19610
rect 81180 19558 81194 19610
rect 81194 19558 81206 19610
rect 81206 19558 81236 19610
rect 81260 19558 81270 19610
rect 81270 19558 81316 19610
rect 81020 19556 81076 19558
rect 81100 19556 81156 19558
rect 81180 19556 81236 19558
rect 81260 19556 81316 19558
rect 81020 18522 81076 18524
rect 81100 18522 81156 18524
rect 81180 18522 81236 18524
rect 81260 18522 81316 18524
rect 81020 18470 81066 18522
rect 81066 18470 81076 18522
rect 81100 18470 81130 18522
rect 81130 18470 81142 18522
rect 81142 18470 81156 18522
rect 81180 18470 81194 18522
rect 81194 18470 81206 18522
rect 81206 18470 81236 18522
rect 81260 18470 81270 18522
rect 81270 18470 81316 18522
rect 81020 18468 81076 18470
rect 81100 18468 81156 18470
rect 81180 18468 81236 18470
rect 81260 18468 81316 18470
rect 81020 17434 81076 17436
rect 81100 17434 81156 17436
rect 81180 17434 81236 17436
rect 81260 17434 81316 17436
rect 81020 17382 81066 17434
rect 81066 17382 81076 17434
rect 81100 17382 81130 17434
rect 81130 17382 81142 17434
rect 81142 17382 81156 17434
rect 81180 17382 81194 17434
rect 81194 17382 81206 17434
rect 81206 17382 81236 17434
rect 81260 17382 81270 17434
rect 81270 17382 81316 17434
rect 81020 17380 81076 17382
rect 81100 17380 81156 17382
rect 81180 17380 81236 17382
rect 81260 17380 81316 17382
rect 81020 16346 81076 16348
rect 81100 16346 81156 16348
rect 81180 16346 81236 16348
rect 81260 16346 81316 16348
rect 81020 16294 81066 16346
rect 81066 16294 81076 16346
rect 81100 16294 81130 16346
rect 81130 16294 81142 16346
rect 81142 16294 81156 16346
rect 81180 16294 81194 16346
rect 81194 16294 81206 16346
rect 81206 16294 81236 16346
rect 81260 16294 81270 16346
rect 81270 16294 81316 16346
rect 81020 16292 81076 16294
rect 81100 16292 81156 16294
rect 81180 16292 81236 16294
rect 81260 16292 81316 16294
rect 81020 15258 81076 15260
rect 81100 15258 81156 15260
rect 81180 15258 81236 15260
rect 81260 15258 81316 15260
rect 81020 15206 81066 15258
rect 81066 15206 81076 15258
rect 81100 15206 81130 15258
rect 81130 15206 81142 15258
rect 81142 15206 81156 15258
rect 81180 15206 81194 15258
rect 81194 15206 81206 15258
rect 81206 15206 81236 15258
rect 81260 15206 81270 15258
rect 81270 15206 81316 15258
rect 81020 15204 81076 15206
rect 81100 15204 81156 15206
rect 81180 15204 81236 15206
rect 81260 15204 81316 15206
rect 81020 14170 81076 14172
rect 81100 14170 81156 14172
rect 81180 14170 81236 14172
rect 81260 14170 81316 14172
rect 81020 14118 81066 14170
rect 81066 14118 81076 14170
rect 81100 14118 81130 14170
rect 81130 14118 81142 14170
rect 81142 14118 81156 14170
rect 81180 14118 81194 14170
rect 81194 14118 81206 14170
rect 81206 14118 81236 14170
rect 81260 14118 81270 14170
rect 81270 14118 81316 14170
rect 81020 14116 81076 14118
rect 81100 14116 81156 14118
rect 81180 14116 81236 14118
rect 81260 14116 81316 14118
rect 81020 13082 81076 13084
rect 81100 13082 81156 13084
rect 81180 13082 81236 13084
rect 81260 13082 81316 13084
rect 81020 13030 81066 13082
rect 81066 13030 81076 13082
rect 81100 13030 81130 13082
rect 81130 13030 81142 13082
rect 81142 13030 81156 13082
rect 81180 13030 81194 13082
rect 81194 13030 81206 13082
rect 81206 13030 81236 13082
rect 81260 13030 81270 13082
rect 81270 13030 81316 13082
rect 81020 13028 81076 13030
rect 81100 13028 81156 13030
rect 81180 13028 81236 13030
rect 81260 13028 81316 13030
rect 81020 11994 81076 11996
rect 81100 11994 81156 11996
rect 81180 11994 81236 11996
rect 81260 11994 81316 11996
rect 81020 11942 81066 11994
rect 81066 11942 81076 11994
rect 81100 11942 81130 11994
rect 81130 11942 81142 11994
rect 81142 11942 81156 11994
rect 81180 11942 81194 11994
rect 81194 11942 81206 11994
rect 81206 11942 81236 11994
rect 81260 11942 81270 11994
rect 81270 11942 81316 11994
rect 81020 11940 81076 11942
rect 81100 11940 81156 11942
rect 81180 11940 81236 11942
rect 81260 11940 81316 11942
rect 81020 10906 81076 10908
rect 81100 10906 81156 10908
rect 81180 10906 81236 10908
rect 81260 10906 81316 10908
rect 81020 10854 81066 10906
rect 81066 10854 81076 10906
rect 81100 10854 81130 10906
rect 81130 10854 81142 10906
rect 81142 10854 81156 10906
rect 81180 10854 81194 10906
rect 81194 10854 81206 10906
rect 81206 10854 81236 10906
rect 81260 10854 81270 10906
rect 81270 10854 81316 10906
rect 81020 10852 81076 10854
rect 81100 10852 81156 10854
rect 81180 10852 81236 10854
rect 81260 10852 81316 10854
rect 81020 9818 81076 9820
rect 81100 9818 81156 9820
rect 81180 9818 81236 9820
rect 81260 9818 81316 9820
rect 81020 9766 81066 9818
rect 81066 9766 81076 9818
rect 81100 9766 81130 9818
rect 81130 9766 81142 9818
rect 81142 9766 81156 9818
rect 81180 9766 81194 9818
rect 81194 9766 81206 9818
rect 81206 9766 81236 9818
rect 81260 9766 81270 9818
rect 81270 9766 81316 9818
rect 81020 9764 81076 9766
rect 81100 9764 81156 9766
rect 81180 9764 81236 9766
rect 81260 9764 81316 9766
rect 81020 8730 81076 8732
rect 81100 8730 81156 8732
rect 81180 8730 81236 8732
rect 81260 8730 81316 8732
rect 81020 8678 81066 8730
rect 81066 8678 81076 8730
rect 81100 8678 81130 8730
rect 81130 8678 81142 8730
rect 81142 8678 81156 8730
rect 81180 8678 81194 8730
rect 81194 8678 81206 8730
rect 81206 8678 81236 8730
rect 81260 8678 81270 8730
rect 81270 8678 81316 8730
rect 81020 8676 81076 8678
rect 81100 8676 81156 8678
rect 81180 8676 81236 8678
rect 81260 8676 81316 8678
rect 81020 7642 81076 7644
rect 81100 7642 81156 7644
rect 81180 7642 81236 7644
rect 81260 7642 81316 7644
rect 81020 7590 81066 7642
rect 81066 7590 81076 7642
rect 81100 7590 81130 7642
rect 81130 7590 81142 7642
rect 81142 7590 81156 7642
rect 81180 7590 81194 7642
rect 81194 7590 81206 7642
rect 81206 7590 81236 7642
rect 81260 7590 81270 7642
rect 81270 7590 81316 7642
rect 81020 7588 81076 7590
rect 81100 7588 81156 7590
rect 81180 7588 81236 7590
rect 81260 7588 81316 7590
rect 81020 6554 81076 6556
rect 81100 6554 81156 6556
rect 81180 6554 81236 6556
rect 81260 6554 81316 6556
rect 81020 6502 81066 6554
rect 81066 6502 81076 6554
rect 81100 6502 81130 6554
rect 81130 6502 81142 6554
rect 81142 6502 81156 6554
rect 81180 6502 81194 6554
rect 81194 6502 81206 6554
rect 81206 6502 81236 6554
rect 81260 6502 81270 6554
rect 81270 6502 81316 6554
rect 81020 6500 81076 6502
rect 81100 6500 81156 6502
rect 81180 6500 81236 6502
rect 81260 6500 81316 6502
rect 81020 5466 81076 5468
rect 81100 5466 81156 5468
rect 81180 5466 81236 5468
rect 81260 5466 81316 5468
rect 81020 5414 81066 5466
rect 81066 5414 81076 5466
rect 81100 5414 81130 5466
rect 81130 5414 81142 5466
rect 81142 5414 81156 5466
rect 81180 5414 81194 5466
rect 81194 5414 81206 5466
rect 81206 5414 81236 5466
rect 81260 5414 81270 5466
rect 81270 5414 81316 5466
rect 81020 5412 81076 5414
rect 81100 5412 81156 5414
rect 81180 5412 81236 5414
rect 81260 5412 81316 5414
rect 81020 4378 81076 4380
rect 81100 4378 81156 4380
rect 81180 4378 81236 4380
rect 81260 4378 81316 4380
rect 81020 4326 81066 4378
rect 81066 4326 81076 4378
rect 81100 4326 81130 4378
rect 81130 4326 81142 4378
rect 81142 4326 81156 4378
rect 81180 4326 81194 4378
rect 81194 4326 81206 4378
rect 81206 4326 81236 4378
rect 81260 4326 81270 4378
rect 81270 4326 81316 4378
rect 81020 4324 81076 4326
rect 81100 4324 81156 4326
rect 81180 4324 81236 4326
rect 81260 4324 81316 4326
rect 81346 3596 81402 3632
rect 81346 3576 81348 3596
rect 81348 3576 81400 3596
rect 81400 3576 81402 3596
rect 81020 3290 81076 3292
rect 81100 3290 81156 3292
rect 81180 3290 81236 3292
rect 81260 3290 81316 3292
rect 81020 3238 81066 3290
rect 81066 3238 81076 3290
rect 81100 3238 81130 3290
rect 81130 3238 81142 3290
rect 81142 3238 81156 3290
rect 81180 3238 81194 3290
rect 81194 3238 81206 3290
rect 81206 3238 81236 3290
rect 81260 3238 81270 3290
rect 81270 3238 81316 3290
rect 81020 3236 81076 3238
rect 81100 3236 81156 3238
rect 81180 3236 81236 3238
rect 81260 3236 81316 3238
rect 81020 2202 81076 2204
rect 81100 2202 81156 2204
rect 81180 2202 81236 2204
rect 81260 2202 81316 2204
rect 81020 2150 81066 2202
rect 81066 2150 81076 2202
rect 81100 2150 81130 2202
rect 81130 2150 81142 2202
rect 81142 2150 81156 2202
rect 81180 2150 81194 2202
rect 81194 2150 81206 2202
rect 81206 2150 81236 2202
rect 81260 2150 81270 2202
rect 81270 2150 81316 2202
rect 81020 2148 81076 2150
rect 81100 2148 81156 2150
rect 81180 2148 81236 2150
rect 81260 2148 81316 2150
rect 84750 36760 84806 36816
rect 84750 36488 84806 36544
rect 84658 36352 84714 36408
rect 85762 37576 85818 37632
rect 83278 3596 83334 3632
rect 83278 3576 83280 3596
rect 83280 3576 83332 3596
rect 83332 3576 83334 3596
rect 89074 33904 89130 33960
rect 96380 37562 96436 37564
rect 96460 37562 96516 37564
rect 96540 37562 96596 37564
rect 96620 37562 96676 37564
rect 96380 37510 96426 37562
rect 96426 37510 96436 37562
rect 96460 37510 96490 37562
rect 96490 37510 96502 37562
rect 96502 37510 96516 37562
rect 96540 37510 96554 37562
rect 96554 37510 96566 37562
rect 96566 37510 96596 37562
rect 96620 37510 96630 37562
rect 96630 37510 96676 37562
rect 96380 37508 96436 37510
rect 96460 37508 96516 37510
rect 96540 37508 96596 37510
rect 96620 37508 96676 37510
rect 96802 37068 96804 37088
rect 96804 37068 96856 37088
rect 96856 37068 96858 37088
rect 96802 37032 96858 37068
rect 92846 34448 92902 34504
rect 92110 34040 92166 34096
rect 95882 33496 95938 33552
rect 96380 36474 96436 36476
rect 96460 36474 96516 36476
rect 96540 36474 96596 36476
rect 96620 36474 96676 36476
rect 96380 36422 96426 36474
rect 96426 36422 96436 36474
rect 96460 36422 96490 36474
rect 96490 36422 96502 36474
rect 96502 36422 96516 36474
rect 96540 36422 96554 36474
rect 96554 36422 96566 36474
rect 96566 36422 96596 36474
rect 96620 36422 96630 36474
rect 96630 36422 96676 36474
rect 96380 36420 96436 36422
rect 96460 36420 96516 36422
rect 96540 36420 96596 36422
rect 96620 36420 96676 36422
rect 96380 35386 96436 35388
rect 96460 35386 96516 35388
rect 96540 35386 96596 35388
rect 96620 35386 96676 35388
rect 96380 35334 96426 35386
rect 96426 35334 96436 35386
rect 96460 35334 96490 35386
rect 96490 35334 96502 35386
rect 96502 35334 96516 35386
rect 96540 35334 96554 35386
rect 96554 35334 96566 35386
rect 96566 35334 96596 35386
rect 96620 35334 96630 35386
rect 96630 35334 96676 35386
rect 96380 35332 96436 35334
rect 96460 35332 96516 35334
rect 96540 35332 96596 35334
rect 96620 35332 96676 35334
rect 96380 34298 96436 34300
rect 96460 34298 96516 34300
rect 96540 34298 96596 34300
rect 96620 34298 96676 34300
rect 96380 34246 96426 34298
rect 96426 34246 96436 34298
rect 96460 34246 96490 34298
rect 96490 34246 96502 34298
rect 96502 34246 96516 34298
rect 96540 34246 96554 34298
rect 96554 34246 96566 34298
rect 96566 34246 96596 34298
rect 96620 34246 96630 34298
rect 96630 34246 96676 34298
rect 96380 34244 96436 34246
rect 96460 34244 96516 34246
rect 96540 34244 96596 34246
rect 96620 34244 96676 34246
rect 96380 33210 96436 33212
rect 96460 33210 96516 33212
rect 96540 33210 96596 33212
rect 96620 33210 96676 33212
rect 96380 33158 96426 33210
rect 96426 33158 96436 33210
rect 96460 33158 96490 33210
rect 96490 33158 96502 33210
rect 96502 33158 96516 33210
rect 96540 33158 96554 33210
rect 96554 33158 96566 33210
rect 96566 33158 96596 33210
rect 96620 33158 96630 33210
rect 96630 33158 96676 33210
rect 96380 33156 96436 33158
rect 96460 33156 96516 33158
rect 96540 33156 96596 33158
rect 96620 33156 96676 33158
rect 96380 32122 96436 32124
rect 96460 32122 96516 32124
rect 96540 32122 96596 32124
rect 96620 32122 96676 32124
rect 96380 32070 96426 32122
rect 96426 32070 96436 32122
rect 96460 32070 96490 32122
rect 96490 32070 96502 32122
rect 96502 32070 96516 32122
rect 96540 32070 96554 32122
rect 96554 32070 96566 32122
rect 96566 32070 96596 32122
rect 96620 32070 96630 32122
rect 96630 32070 96676 32122
rect 96380 32068 96436 32070
rect 96460 32068 96516 32070
rect 96540 32068 96596 32070
rect 96620 32068 96676 32070
rect 96380 31034 96436 31036
rect 96460 31034 96516 31036
rect 96540 31034 96596 31036
rect 96620 31034 96676 31036
rect 96380 30982 96426 31034
rect 96426 30982 96436 31034
rect 96460 30982 96490 31034
rect 96490 30982 96502 31034
rect 96502 30982 96516 31034
rect 96540 30982 96554 31034
rect 96554 30982 96566 31034
rect 96566 30982 96596 31034
rect 96620 30982 96630 31034
rect 96630 30982 96676 31034
rect 96380 30980 96436 30982
rect 96460 30980 96516 30982
rect 96540 30980 96596 30982
rect 96620 30980 96676 30982
rect 96380 29946 96436 29948
rect 96460 29946 96516 29948
rect 96540 29946 96596 29948
rect 96620 29946 96676 29948
rect 96380 29894 96426 29946
rect 96426 29894 96436 29946
rect 96460 29894 96490 29946
rect 96490 29894 96502 29946
rect 96502 29894 96516 29946
rect 96540 29894 96554 29946
rect 96554 29894 96566 29946
rect 96566 29894 96596 29946
rect 96620 29894 96630 29946
rect 96630 29894 96676 29946
rect 96380 29892 96436 29894
rect 96460 29892 96516 29894
rect 96540 29892 96596 29894
rect 96620 29892 96676 29894
rect 96380 28858 96436 28860
rect 96460 28858 96516 28860
rect 96540 28858 96596 28860
rect 96620 28858 96676 28860
rect 96380 28806 96426 28858
rect 96426 28806 96436 28858
rect 96460 28806 96490 28858
rect 96490 28806 96502 28858
rect 96502 28806 96516 28858
rect 96540 28806 96554 28858
rect 96554 28806 96566 28858
rect 96566 28806 96596 28858
rect 96620 28806 96630 28858
rect 96630 28806 96676 28858
rect 96380 28804 96436 28806
rect 96460 28804 96516 28806
rect 96540 28804 96596 28806
rect 96620 28804 96676 28806
rect 96380 27770 96436 27772
rect 96460 27770 96516 27772
rect 96540 27770 96596 27772
rect 96620 27770 96676 27772
rect 96380 27718 96426 27770
rect 96426 27718 96436 27770
rect 96460 27718 96490 27770
rect 96490 27718 96502 27770
rect 96502 27718 96516 27770
rect 96540 27718 96554 27770
rect 96554 27718 96566 27770
rect 96566 27718 96596 27770
rect 96620 27718 96630 27770
rect 96630 27718 96676 27770
rect 96380 27716 96436 27718
rect 96460 27716 96516 27718
rect 96540 27716 96596 27718
rect 96620 27716 96676 27718
rect 96380 26682 96436 26684
rect 96460 26682 96516 26684
rect 96540 26682 96596 26684
rect 96620 26682 96676 26684
rect 96380 26630 96426 26682
rect 96426 26630 96436 26682
rect 96460 26630 96490 26682
rect 96490 26630 96502 26682
rect 96502 26630 96516 26682
rect 96540 26630 96554 26682
rect 96554 26630 96566 26682
rect 96566 26630 96596 26682
rect 96620 26630 96630 26682
rect 96630 26630 96676 26682
rect 96380 26628 96436 26630
rect 96460 26628 96516 26630
rect 96540 26628 96596 26630
rect 96620 26628 96676 26630
rect 96380 25594 96436 25596
rect 96460 25594 96516 25596
rect 96540 25594 96596 25596
rect 96620 25594 96676 25596
rect 96380 25542 96426 25594
rect 96426 25542 96436 25594
rect 96460 25542 96490 25594
rect 96490 25542 96502 25594
rect 96502 25542 96516 25594
rect 96540 25542 96554 25594
rect 96554 25542 96566 25594
rect 96566 25542 96596 25594
rect 96620 25542 96630 25594
rect 96630 25542 96676 25594
rect 96380 25540 96436 25542
rect 96460 25540 96516 25542
rect 96540 25540 96596 25542
rect 96620 25540 96676 25542
rect 96380 24506 96436 24508
rect 96460 24506 96516 24508
rect 96540 24506 96596 24508
rect 96620 24506 96676 24508
rect 96380 24454 96426 24506
rect 96426 24454 96436 24506
rect 96460 24454 96490 24506
rect 96490 24454 96502 24506
rect 96502 24454 96516 24506
rect 96540 24454 96554 24506
rect 96554 24454 96566 24506
rect 96566 24454 96596 24506
rect 96620 24454 96630 24506
rect 96630 24454 96676 24506
rect 96380 24452 96436 24454
rect 96460 24452 96516 24454
rect 96540 24452 96596 24454
rect 96620 24452 96676 24454
rect 96380 23418 96436 23420
rect 96460 23418 96516 23420
rect 96540 23418 96596 23420
rect 96620 23418 96676 23420
rect 96380 23366 96426 23418
rect 96426 23366 96436 23418
rect 96460 23366 96490 23418
rect 96490 23366 96502 23418
rect 96502 23366 96516 23418
rect 96540 23366 96554 23418
rect 96554 23366 96566 23418
rect 96566 23366 96596 23418
rect 96620 23366 96630 23418
rect 96630 23366 96676 23418
rect 96380 23364 96436 23366
rect 96460 23364 96516 23366
rect 96540 23364 96596 23366
rect 96620 23364 96676 23366
rect 96380 22330 96436 22332
rect 96460 22330 96516 22332
rect 96540 22330 96596 22332
rect 96620 22330 96676 22332
rect 96380 22278 96426 22330
rect 96426 22278 96436 22330
rect 96460 22278 96490 22330
rect 96490 22278 96502 22330
rect 96502 22278 96516 22330
rect 96540 22278 96554 22330
rect 96554 22278 96566 22330
rect 96566 22278 96596 22330
rect 96620 22278 96630 22330
rect 96630 22278 96676 22330
rect 96380 22276 96436 22278
rect 96460 22276 96516 22278
rect 96540 22276 96596 22278
rect 96620 22276 96676 22278
rect 96380 21242 96436 21244
rect 96460 21242 96516 21244
rect 96540 21242 96596 21244
rect 96620 21242 96676 21244
rect 96380 21190 96426 21242
rect 96426 21190 96436 21242
rect 96460 21190 96490 21242
rect 96490 21190 96502 21242
rect 96502 21190 96516 21242
rect 96540 21190 96554 21242
rect 96554 21190 96566 21242
rect 96566 21190 96596 21242
rect 96620 21190 96630 21242
rect 96630 21190 96676 21242
rect 96380 21188 96436 21190
rect 96460 21188 96516 21190
rect 96540 21188 96596 21190
rect 96620 21188 96676 21190
rect 96380 20154 96436 20156
rect 96460 20154 96516 20156
rect 96540 20154 96596 20156
rect 96620 20154 96676 20156
rect 96380 20102 96426 20154
rect 96426 20102 96436 20154
rect 96460 20102 96490 20154
rect 96490 20102 96502 20154
rect 96502 20102 96516 20154
rect 96540 20102 96554 20154
rect 96554 20102 96566 20154
rect 96566 20102 96596 20154
rect 96620 20102 96630 20154
rect 96630 20102 96676 20154
rect 96380 20100 96436 20102
rect 96460 20100 96516 20102
rect 96540 20100 96596 20102
rect 96620 20100 96676 20102
rect 96380 19066 96436 19068
rect 96460 19066 96516 19068
rect 96540 19066 96596 19068
rect 96620 19066 96676 19068
rect 96380 19014 96426 19066
rect 96426 19014 96436 19066
rect 96460 19014 96490 19066
rect 96490 19014 96502 19066
rect 96502 19014 96516 19066
rect 96540 19014 96554 19066
rect 96554 19014 96566 19066
rect 96566 19014 96596 19066
rect 96620 19014 96630 19066
rect 96630 19014 96676 19066
rect 96380 19012 96436 19014
rect 96460 19012 96516 19014
rect 96540 19012 96596 19014
rect 96620 19012 96676 19014
rect 96380 17978 96436 17980
rect 96460 17978 96516 17980
rect 96540 17978 96596 17980
rect 96620 17978 96676 17980
rect 96380 17926 96426 17978
rect 96426 17926 96436 17978
rect 96460 17926 96490 17978
rect 96490 17926 96502 17978
rect 96502 17926 96516 17978
rect 96540 17926 96554 17978
rect 96554 17926 96566 17978
rect 96566 17926 96596 17978
rect 96620 17926 96630 17978
rect 96630 17926 96676 17978
rect 96380 17924 96436 17926
rect 96460 17924 96516 17926
rect 96540 17924 96596 17926
rect 96620 17924 96676 17926
rect 96380 16890 96436 16892
rect 96460 16890 96516 16892
rect 96540 16890 96596 16892
rect 96620 16890 96676 16892
rect 96380 16838 96426 16890
rect 96426 16838 96436 16890
rect 96460 16838 96490 16890
rect 96490 16838 96502 16890
rect 96502 16838 96516 16890
rect 96540 16838 96554 16890
rect 96554 16838 96566 16890
rect 96566 16838 96596 16890
rect 96620 16838 96630 16890
rect 96630 16838 96676 16890
rect 96380 16836 96436 16838
rect 96460 16836 96516 16838
rect 96540 16836 96596 16838
rect 96620 16836 96676 16838
rect 96380 15802 96436 15804
rect 96460 15802 96516 15804
rect 96540 15802 96596 15804
rect 96620 15802 96676 15804
rect 96380 15750 96426 15802
rect 96426 15750 96436 15802
rect 96460 15750 96490 15802
rect 96490 15750 96502 15802
rect 96502 15750 96516 15802
rect 96540 15750 96554 15802
rect 96554 15750 96566 15802
rect 96566 15750 96596 15802
rect 96620 15750 96630 15802
rect 96630 15750 96676 15802
rect 96380 15748 96436 15750
rect 96460 15748 96516 15750
rect 96540 15748 96596 15750
rect 96620 15748 96676 15750
rect 96380 14714 96436 14716
rect 96460 14714 96516 14716
rect 96540 14714 96596 14716
rect 96620 14714 96676 14716
rect 96380 14662 96426 14714
rect 96426 14662 96436 14714
rect 96460 14662 96490 14714
rect 96490 14662 96502 14714
rect 96502 14662 96516 14714
rect 96540 14662 96554 14714
rect 96554 14662 96566 14714
rect 96566 14662 96596 14714
rect 96620 14662 96630 14714
rect 96630 14662 96676 14714
rect 96380 14660 96436 14662
rect 96460 14660 96516 14662
rect 96540 14660 96596 14662
rect 96620 14660 96676 14662
rect 96380 13626 96436 13628
rect 96460 13626 96516 13628
rect 96540 13626 96596 13628
rect 96620 13626 96676 13628
rect 96380 13574 96426 13626
rect 96426 13574 96436 13626
rect 96460 13574 96490 13626
rect 96490 13574 96502 13626
rect 96502 13574 96516 13626
rect 96540 13574 96554 13626
rect 96554 13574 96566 13626
rect 96566 13574 96596 13626
rect 96620 13574 96630 13626
rect 96630 13574 96676 13626
rect 96380 13572 96436 13574
rect 96460 13572 96516 13574
rect 96540 13572 96596 13574
rect 96620 13572 96676 13574
rect 96380 12538 96436 12540
rect 96460 12538 96516 12540
rect 96540 12538 96596 12540
rect 96620 12538 96676 12540
rect 96380 12486 96426 12538
rect 96426 12486 96436 12538
rect 96460 12486 96490 12538
rect 96490 12486 96502 12538
rect 96502 12486 96516 12538
rect 96540 12486 96554 12538
rect 96554 12486 96566 12538
rect 96566 12486 96596 12538
rect 96620 12486 96630 12538
rect 96630 12486 96676 12538
rect 96380 12484 96436 12486
rect 96460 12484 96516 12486
rect 96540 12484 96596 12486
rect 96620 12484 96676 12486
rect 96380 11450 96436 11452
rect 96460 11450 96516 11452
rect 96540 11450 96596 11452
rect 96620 11450 96676 11452
rect 96380 11398 96426 11450
rect 96426 11398 96436 11450
rect 96460 11398 96490 11450
rect 96490 11398 96502 11450
rect 96502 11398 96516 11450
rect 96540 11398 96554 11450
rect 96554 11398 96566 11450
rect 96566 11398 96596 11450
rect 96620 11398 96630 11450
rect 96630 11398 96676 11450
rect 96380 11396 96436 11398
rect 96460 11396 96516 11398
rect 96540 11396 96596 11398
rect 96620 11396 96676 11398
rect 96380 10362 96436 10364
rect 96460 10362 96516 10364
rect 96540 10362 96596 10364
rect 96620 10362 96676 10364
rect 96380 10310 96426 10362
rect 96426 10310 96436 10362
rect 96460 10310 96490 10362
rect 96490 10310 96502 10362
rect 96502 10310 96516 10362
rect 96540 10310 96554 10362
rect 96554 10310 96566 10362
rect 96566 10310 96596 10362
rect 96620 10310 96630 10362
rect 96630 10310 96676 10362
rect 96380 10308 96436 10310
rect 96460 10308 96516 10310
rect 96540 10308 96596 10310
rect 96620 10308 96676 10310
rect 96380 9274 96436 9276
rect 96460 9274 96516 9276
rect 96540 9274 96596 9276
rect 96620 9274 96676 9276
rect 96380 9222 96426 9274
rect 96426 9222 96436 9274
rect 96460 9222 96490 9274
rect 96490 9222 96502 9274
rect 96502 9222 96516 9274
rect 96540 9222 96554 9274
rect 96554 9222 96566 9274
rect 96566 9222 96596 9274
rect 96620 9222 96630 9274
rect 96630 9222 96676 9274
rect 96380 9220 96436 9222
rect 96460 9220 96516 9222
rect 96540 9220 96596 9222
rect 96620 9220 96676 9222
rect 96380 8186 96436 8188
rect 96460 8186 96516 8188
rect 96540 8186 96596 8188
rect 96620 8186 96676 8188
rect 96380 8134 96426 8186
rect 96426 8134 96436 8186
rect 96460 8134 96490 8186
rect 96490 8134 96502 8186
rect 96502 8134 96516 8186
rect 96540 8134 96554 8186
rect 96554 8134 96566 8186
rect 96566 8134 96596 8186
rect 96620 8134 96630 8186
rect 96630 8134 96676 8186
rect 96380 8132 96436 8134
rect 96460 8132 96516 8134
rect 96540 8132 96596 8134
rect 96620 8132 96676 8134
rect 96380 7098 96436 7100
rect 96460 7098 96516 7100
rect 96540 7098 96596 7100
rect 96620 7098 96676 7100
rect 96380 7046 96426 7098
rect 96426 7046 96436 7098
rect 96460 7046 96490 7098
rect 96490 7046 96502 7098
rect 96502 7046 96516 7098
rect 96540 7046 96554 7098
rect 96554 7046 96566 7098
rect 96566 7046 96596 7098
rect 96620 7046 96630 7098
rect 96630 7046 96676 7098
rect 96380 7044 96436 7046
rect 96460 7044 96516 7046
rect 96540 7044 96596 7046
rect 96620 7044 96676 7046
rect 96380 6010 96436 6012
rect 96460 6010 96516 6012
rect 96540 6010 96596 6012
rect 96620 6010 96676 6012
rect 96380 5958 96426 6010
rect 96426 5958 96436 6010
rect 96460 5958 96490 6010
rect 96490 5958 96502 6010
rect 96502 5958 96516 6010
rect 96540 5958 96554 6010
rect 96554 5958 96566 6010
rect 96566 5958 96596 6010
rect 96620 5958 96630 6010
rect 96630 5958 96676 6010
rect 96380 5956 96436 5958
rect 96460 5956 96516 5958
rect 96540 5956 96596 5958
rect 96620 5956 96676 5958
rect 96380 4922 96436 4924
rect 96460 4922 96516 4924
rect 96540 4922 96596 4924
rect 96620 4922 96676 4924
rect 96380 4870 96426 4922
rect 96426 4870 96436 4922
rect 96460 4870 96490 4922
rect 96490 4870 96502 4922
rect 96502 4870 96516 4922
rect 96540 4870 96554 4922
rect 96554 4870 96566 4922
rect 96566 4870 96596 4922
rect 96620 4870 96630 4922
rect 96630 4870 96676 4922
rect 96380 4868 96436 4870
rect 96460 4868 96516 4870
rect 96540 4868 96596 4870
rect 96620 4868 96676 4870
rect 96380 3834 96436 3836
rect 96460 3834 96516 3836
rect 96540 3834 96596 3836
rect 96620 3834 96676 3836
rect 96380 3782 96426 3834
rect 96426 3782 96436 3834
rect 96460 3782 96490 3834
rect 96490 3782 96502 3834
rect 96502 3782 96516 3834
rect 96540 3782 96554 3834
rect 96554 3782 96566 3834
rect 96566 3782 96596 3834
rect 96620 3782 96630 3834
rect 96630 3782 96676 3834
rect 96380 3780 96436 3782
rect 96460 3780 96516 3782
rect 96540 3780 96596 3782
rect 96620 3780 96676 3782
rect 96380 2746 96436 2748
rect 96460 2746 96516 2748
rect 96540 2746 96596 2748
rect 96620 2746 96676 2748
rect 96380 2694 96426 2746
rect 96426 2694 96436 2746
rect 96460 2694 96490 2746
rect 96490 2694 96502 2746
rect 96502 2694 96516 2746
rect 96540 2694 96554 2746
rect 96554 2694 96566 2746
rect 96566 2694 96596 2746
rect 96620 2694 96630 2746
rect 96630 2694 96676 2746
rect 96380 2692 96436 2694
rect 96460 2692 96516 2694
rect 96540 2692 96596 2694
rect 96620 2692 96676 2694
rect 100206 36624 100262 36680
rect 98366 35536 98422 35592
rect 102690 36080 102746 36136
rect 105358 36216 105414 36272
rect 107106 36760 107162 36816
rect 109406 36760 109462 36816
rect 110234 36352 110290 36408
rect 111740 37018 111796 37020
rect 111820 37018 111876 37020
rect 111900 37018 111956 37020
rect 111980 37018 112036 37020
rect 111740 36966 111786 37018
rect 111786 36966 111796 37018
rect 111820 36966 111850 37018
rect 111850 36966 111862 37018
rect 111862 36966 111876 37018
rect 111900 36966 111914 37018
rect 111914 36966 111926 37018
rect 111926 36966 111956 37018
rect 111980 36966 111990 37018
rect 111990 36966 112036 37018
rect 111740 36964 111796 36966
rect 111820 36964 111876 36966
rect 111900 36964 111956 36966
rect 111980 36964 112036 36966
rect 111890 36624 111946 36680
rect 111740 35930 111796 35932
rect 111820 35930 111876 35932
rect 111900 35930 111956 35932
rect 111980 35930 112036 35932
rect 111740 35878 111786 35930
rect 111786 35878 111796 35930
rect 111820 35878 111850 35930
rect 111850 35878 111862 35930
rect 111862 35878 111876 35930
rect 111900 35878 111914 35930
rect 111914 35878 111926 35930
rect 111926 35878 111956 35930
rect 111980 35878 111990 35930
rect 111990 35878 112036 35930
rect 111740 35876 111796 35878
rect 111820 35876 111876 35878
rect 111900 35876 111956 35878
rect 111980 35876 112036 35878
rect 111740 34842 111796 34844
rect 111820 34842 111876 34844
rect 111900 34842 111956 34844
rect 111980 34842 112036 34844
rect 111740 34790 111786 34842
rect 111786 34790 111796 34842
rect 111820 34790 111850 34842
rect 111850 34790 111862 34842
rect 111862 34790 111876 34842
rect 111900 34790 111914 34842
rect 111914 34790 111926 34842
rect 111926 34790 111956 34842
rect 111980 34790 111990 34842
rect 111990 34790 112036 34842
rect 111740 34788 111796 34790
rect 111820 34788 111876 34790
rect 111900 34788 111956 34790
rect 111980 34788 112036 34790
rect 111740 33754 111796 33756
rect 111820 33754 111876 33756
rect 111900 33754 111956 33756
rect 111980 33754 112036 33756
rect 111740 33702 111786 33754
rect 111786 33702 111796 33754
rect 111820 33702 111850 33754
rect 111850 33702 111862 33754
rect 111862 33702 111876 33754
rect 111900 33702 111914 33754
rect 111914 33702 111926 33754
rect 111926 33702 111956 33754
rect 111980 33702 111990 33754
rect 111990 33702 112036 33754
rect 111740 33700 111796 33702
rect 111820 33700 111876 33702
rect 111900 33700 111956 33702
rect 111980 33700 112036 33702
rect 115846 36352 115902 36408
rect 111740 32666 111796 32668
rect 111820 32666 111876 32668
rect 111900 32666 111956 32668
rect 111980 32666 112036 32668
rect 111740 32614 111786 32666
rect 111786 32614 111796 32666
rect 111820 32614 111850 32666
rect 111850 32614 111862 32666
rect 111862 32614 111876 32666
rect 111900 32614 111914 32666
rect 111914 32614 111926 32666
rect 111926 32614 111956 32666
rect 111980 32614 111990 32666
rect 111990 32614 112036 32666
rect 111740 32612 111796 32614
rect 111820 32612 111876 32614
rect 111900 32612 111956 32614
rect 111980 32612 112036 32614
rect 111740 31578 111796 31580
rect 111820 31578 111876 31580
rect 111900 31578 111956 31580
rect 111980 31578 112036 31580
rect 111740 31526 111786 31578
rect 111786 31526 111796 31578
rect 111820 31526 111850 31578
rect 111850 31526 111862 31578
rect 111862 31526 111876 31578
rect 111900 31526 111914 31578
rect 111914 31526 111926 31578
rect 111926 31526 111956 31578
rect 111980 31526 111990 31578
rect 111990 31526 112036 31578
rect 111740 31524 111796 31526
rect 111820 31524 111876 31526
rect 111900 31524 111956 31526
rect 111980 31524 112036 31526
rect 111740 30490 111796 30492
rect 111820 30490 111876 30492
rect 111900 30490 111956 30492
rect 111980 30490 112036 30492
rect 111740 30438 111786 30490
rect 111786 30438 111796 30490
rect 111820 30438 111850 30490
rect 111850 30438 111862 30490
rect 111862 30438 111876 30490
rect 111900 30438 111914 30490
rect 111914 30438 111926 30490
rect 111926 30438 111956 30490
rect 111980 30438 111990 30490
rect 111990 30438 112036 30490
rect 111740 30436 111796 30438
rect 111820 30436 111876 30438
rect 111900 30436 111956 30438
rect 111980 30436 112036 30438
rect 111740 29402 111796 29404
rect 111820 29402 111876 29404
rect 111900 29402 111956 29404
rect 111980 29402 112036 29404
rect 111740 29350 111786 29402
rect 111786 29350 111796 29402
rect 111820 29350 111850 29402
rect 111850 29350 111862 29402
rect 111862 29350 111876 29402
rect 111900 29350 111914 29402
rect 111914 29350 111926 29402
rect 111926 29350 111956 29402
rect 111980 29350 111990 29402
rect 111990 29350 112036 29402
rect 111740 29348 111796 29350
rect 111820 29348 111876 29350
rect 111900 29348 111956 29350
rect 111980 29348 112036 29350
rect 111740 28314 111796 28316
rect 111820 28314 111876 28316
rect 111900 28314 111956 28316
rect 111980 28314 112036 28316
rect 111740 28262 111786 28314
rect 111786 28262 111796 28314
rect 111820 28262 111850 28314
rect 111850 28262 111862 28314
rect 111862 28262 111876 28314
rect 111900 28262 111914 28314
rect 111914 28262 111926 28314
rect 111926 28262 111956 28314
rect 111980 28262 111990 28314
rect 111990 28262 112036 28314
rect 111740 28260 111796 28262
rect 111820 28260 111876 28262
rect 111900 28260 111956 28262
rect 111980 28260 112036 28262
rect 111740 27226 111796 27228
rect 111820 27226 111876 27228
rect 111900 27226 111956 27228
rect 111980 27226 112036 27228
rect 111740 27174 111786 27226
rect 111786 27174 111796 27226
rect 111820 27174 111850 27226
rect 111850 27174 111862 27226
rect 111862 27174 111876 27226
rect 111900 27174 111914 27226
rect 111914 27174 111926 27226
rect 111926 27174 111956 27226
rect 111980 27174 111990 27226
rect 111990 27174 112036 27226
rect 111740 27172 111796 27174
rect 111820 27172 111876 27174
rect 111900 27172 111956 27174
rect 111980 27172 112036 27174
rect 111740 26138 111796 26140
rect 111820 26138 111876 26140
rect 111900 26138 111956 26140
rect 111980 26138 112036 26140
rect 111740 26086 111786 26138
rect 111786 26086 111796 26138
rect 111820 26086 111850 26138
rect 111850 26086 111862 26138
rect 111862 26086 111876 26138
rect 111900 26086 111914 26138
rect 111914 26086 111926 26138
rect 111926 26086 111956 26138
rect 111980 26086 111990 26138
rect 111990 26086 112036 26138
rect 111740 26084 111796 26086
rect 111820 26084 111876 26086
rect 111900 26084 111956 26086
rect 111980 26084 112036 26086
rect 111740 25050 111796 25052
rect 111820 25050 111876 25052
rect 111900 25050 111956 25052
rect 111980 25050 112036 25052
rect 111740 24998 111786 25050
rect 111786 24998 111796 25050
rect 111820 24998 111850 25050
rect 111850 24998 111862 25050
rect 111862 24998 111876 25050
rect 111900 24998 111914 25050
rect 111914 24998 111926 25050
rect 111926 24998 111956 25050
rect 111980 24998 111990 25050
rect 111990 24998 112036 25050
rect 111740 24996 111796 24998
rect 111820 24996 111876 24998
rect 111900 24996 111956 24998
rect 111980 24996 112036 24998
rect 111740 23962 111796 23964
rect 111820 23962 111876 23964
rect 111900 23962 111956 23964
rect 111980 23962 112036 23964
rect 111740 23910 111786 23962
rect 111786 23910 111796 23962
rect 111820 23910 111850 23962
rect 111850 23910 111862 23962
rect 111862 23910 111876 23962
rect 111900 23910 111914 23962
rect 111914 23910 111926 23962
rect 111926 23910 111956 23962
rect 111980 23910 111990 23962
rect 111990 23910 112036 23962
rect 111740 23908 111796 23910
rect 111820 23908 111876 23910
rect 111900 23908 111956 23910
rect 111980 23908 112036 23910
rect 111740 22874 111796 22876
rect 111820 22874 111876 22876
rect 111900 22874 111956 22876
rect 111980 22874 112036 22876
rect 111740 22822 111786 22874
rect 111786 22822 111796 22874
rect 111820 22822 111850 22874
rect 111850 22822 111862 22874
rect 111862 22822 111876 22874
rect 111900 22822 111914 22874
rect 111914 22822 111926 22874
rect 111926 22822 111956 22874
rect 111980 22822 111990 22874
rect 111990 22822 112036 22874
rect 111740 22820 111796 22822
rect 111820 22820 111876 22822
rect 111900 22820 111956 22822
rect 111980 22820 112036 22822
rect 111740 21786 111796 21788
rect 111820 21786 111876 21788
rect 111900 21786 111956 21788
rect 111980 21786 112036 21788
rect 111740 21734 111786 21786
rect 111786 21734 111796 21786
rect 111820 21734 111850 21786
rect 111850 21734 111862 21786
rect 111862 21734 111876 21786
rect 111900 21734 111914 21786
rect 111914 21734 111926 21786
rect 111926 21734 111956 21786
rect 111980 21734 111990 21786
rect 111990 21734 112036 21786
rect 111740 21732 111796 21734
rect 111820 21732 111876 21734
rect 111900 21732 111956 21734
rect 111980 21732 112036 21734
rect 111740 20698 111796 20700
rect 111820 20698 111876 20700
rect 111900 20698 111956 20700
rect 111980 20698 112036 20700
rect 111740 20646 111786 20698
rect 111786 20646 111796 20698
rect 111820 20646 111850 20698
rect 111850 20646 111862 20698
rect 111862 20646 111876 20698
rect 111900 20646 111914 20698
rect 111914 20646 111926 20698
rect 111926 20646 111956 20698
rect 111980 20646 111990 20698
rect 111990 20646 112036 20698
rect 111740 20644 111796 20646
rect 111820 20644 111876 20646
rect 111900 20644 111956 20646
rect 111980 20644 112036 20646
rect 111740 19610 111796 19612
rect 111820 19610 111876 19612
rect 111900 19610 111956 19612
rect 111980 19610 112036 19612
rect 111740 19558 111786 19610
rect 111786 19558 111796 19610
rect 111820 19558 111850 19610
rect 111850 19558 111862 19610
rect 111862 19558 111876 19610
rect 111900 19558 111914 19610
rect 111914 19558 111926 19610
rect 111926 19558 111956 19610
rect 111980 19558 111990 19610
rect 111990 19558 112036 19610
rect 111740 19556 111796 19558
rect 111820 19556 111876 19558
rect 111900 19556 111956 19558
rect 111980 19556 112036 19558
rect 111740 18522 111796 18524
rect 111820 18522 111876 18524
rect 111900 18522 111956 18524
rect 111980 18522 112036 18524
rect 111740 18470 111786 18522
rect 111786 18470 111796 18522
rect 111820 18470 111850 18522
rect 111850 18470 111862 18522
rect 111862 18470 111876 18522
rect 111900 18470 111914 18522
rect 111914 18470 111926 18522
rect 111926 18470 111956 18522
rect 111980 18470 111990 18522
rect 111990 18470 112036 18522
rect 111740 18468 111796 18470
rect 111820 18468 111876 18470
rect 111900 18468 111956 18470
rect 111980 18468 112036 18470
rect 111740 17434 111796 17436
rect 111820 17434 111876 17436
rect 111900 17434 111956 17436
rect 111980 17434 112036 17436
rect 111740 17382 111786 17434
rect 111786 17382 111796 17434
rect 111820 17382 111850 17434
rect 111850 17382 111862 17434
rect 111862 17382 111876 17434
rect 111900 17382 111914 17434
rect 111914 17382 111926 17434
rect 111926 17382 111956 17434
rect 111980 17382 111990 17434
rect 111990 17382 112036 17434
rect 111740 17380 111796 17382
rect 111820 17380 111876 17382
rect 111900 17380 111956 17382
rect 111980 17380 112036 17382
rect 111740 16346 111796 16348
rect 111820 16346 111876 16348
rect 111900 16346 111956 16348
rect 111980 16346 112036 16348
rect 111740 16294 111786 16346
rect 111786 16294 111796 16346
rect 111820 16294 111850 16346
rect 111850 16294 111862 16346
rect 111862 16294 111876 16346
rect 111900 16294 111914 16346
rect 111914 16294 111926 16346
rect 111926 16294 111956 16346
rect 111980 16294 111990 16346
rect 111990 16294 112036 16346
rect 111740 16292 111796 16294
rect 111820 16292 111876 16294
rect 111900 16292 111956 16294
rect 111980 16292 112036 16294
rect 111740 15258 111796 15260
rect 111820 15258 111876 15260
rect 111900 15258 111956 15260
rect 111980 15258 112036 15260
rect 111740 15206 111786 15258
rect 111786 15206 111796 15258
rect 111820 15206 111850 15258
rect 111850 15206 111862 15258
rect 111862 15206 111876 15258
rect 111900 15206 111914 15258
rect 111914 15206 111926 15258
rect 111926 15206 111956 15258
rect 111980 15206 111990 15258
rect 111990 15206 112036 15258
rect 111740 15204 111796 15206
rect 111820 15204 111876 15206
rect 111900 15204 111956 15206
rect 111980 15204 112036 15206
rect 111740 14170 111796 14172
rect 111820 14170 111876 14172
rect 111900 14170 111956 14172
rect 111980 14170 112036 14172
rect 111740 14118 111786 14170
rect 111786 14118 111796 14170
rect 111820 14118 111850 14170
rect 111850 14118 111862 14170
rect 111862 14118 111876 14170
rect 111900 14118 111914 14170
rect 111914 14118 111926 14170
rect 111926 14118 111956 14170
rect 111980 14118 111990 14170
rect 111990 14118 112036 14170
rect 111740 14116 111796 14118
rect 111820 14116 111876 14118
rect 111900 14116 111956 14118
rect 111980 14116 112036 14118
rect 111740 13082 111796 13084
rect 111820 13082 111876 13084
rect 111900 13082 111956 13084
rect 111980 13082 112036 13084
rect 111740 13030 111786 13082
rect 111786 13030 111796 13082
rect 111820 13030 111850 13082
rect 111850 13030 111862 13082
rect 111862 13030 111876 13082
rect 111900 13030 111914 13082
rect 111914 13030 111926 13082
rect 111926 13030 111956 13082
rect 111980 13030 111990 13082
rect 111990 13030 112036 13082
rect 111740 13028 111796 13030
rect 111820 13028 111876 13030
rect 111900 13028 111956 13030
rect 111980 13028 112036 13030
rect 111740 11994 111796 11996
rect 111820 11994 111876 11996
rect 111900 11994 111956 11996
rect 111980 11994 112036 11996
rect 111740 11942 111786 11994
rect 111786 11942 111796 11994
rect 111820 11942 111850 11994
rect 111850 11942 111862 11994
rect 111862 11942 111876 11994
rect 111900 11942 111914 11994
rect 111914 11942 111926 11994
rect 111926 11942 111956 11994
rect 111980 11942 111990 11994
rect 111990 11942 112036 11994
rect 111740 11940 111796 11942
rect 111820 11940 111876 11942
rect 111900 11940 111956 11942
rect 111980 11940 112036 11942
rect 111740 10906 111796 10908
rect 111820 10906 111876 10908
rect 111900 10906 111956 10908
rect 111980 10906 112036 10908
rect 111740 10854 111786 10906
rect 111786 10854 111796 10906
rect 111820 10854 111850 10906
rect 111850 10854 111862 10906
rect 111862 10854 111876 10906
rect 111900 10854 111914 10906
rect 111914 10854 111926 10906
rect 111926 10854 111956 10906
rect 111980 10854 111990 10906
rect 111990 10854 112036 10906
rect 111740 10852 111796 10854
rect 111820 10852 111876 10854
rect 111900 10852 111956 10854
rect 111980 10852 112036 10854
rect 111740 9818 111796 9820
rect 111820 9818 111876 9820
rect 111900 9818 111956 9820
rect 111980 9818 112036 9820
rect 111740 9766 111786 9818
rect 111786 9766 111796 9818
rect 111820 9766 111850 9818
rect 111850 9766 111862 9818
rect 111862 9766 111876 9818
rect 111900 9766 111914 9818
rect 111914 9766 111926 9818
rect 111926 9766 111956 9818
rect 111980 9766 111990 9818
rect 111990 9766 112036 9818
rect 111740 9764 111796 9766
rect 111820 9764 111876 9766
rect 111900 9764 111956 9766
rect 111980 9764 112036 9766
rect 111740 8730 111796 8732
rect 111820 8730 111876 8732
rect 111900 8730 111956 8732
rect 111980 8730 112036 8732
rect 111740 8678 111786 8730
rect 111786 8678 111796 8730
rect 111820 8678 111850 8730
rect 111850 8678 111862 8730
rect 111862 8678 111876 8730
rect 111900 8678 111914 8730
rect 111914 8678 111926 8730
rect 111926 8678 111956 8730
rect 111980 8678 111990 8730
rect 111990 8678 112036 8730
rect 111740 8676 111796 8678
rect 111820 8676 111876 8678
rect 111900 8676 111956 8678
rect 111980 8676 112036 8678
rect 111740 7642 111796 7644
rect 111820 7642 111876 7644
rect 111900 7642 111956 7644
rect 111980 7642 112036 7644
rect 111740 7590 111786 7642
rect 111786 7590 111796 7642
rect 111820 7590 111850 7642
rect 111850 7590 111862 7642
rect 111862 7590 111876 7642
rect 111900 7590 111914 7642
rect 111914 7590 111926 7642
rect 111926 7590 111956 7642
rect 111980 7590 111990 7642
rect 111990 7590 112036 7642
rect 111740 7588 111796 7590
rect 111820 7588 111876 7590
rect 111900 7588 111956 7590
rect 111980 7588 112036 7590
rect 111740 6554 111796 6556
rect 111820 6554 111876 6556
rect 111900 6554 111956 6556
rect 111980 6554 112036 6556
rect 111740 6502 111786 6554
rect 111786 6502 111796 6554
rect 111820 6502 111850 6554
rect 111850 6502 111862 6554
rect 111862 6502 111876 6554
rect 111900 6502 111914 6554
rect 111914 6502 111926 6554
rect 111926 6502 111956 6554
rect 111980 6502 111990 6554
rect 111990 6502 112036 6554
rect 111740 6500 111796 6502
rect 111820 6500 111876 6502
rect 111900 6500 111956 6502
rect 111980 6500 112036 6502
rect 111740 5466 111796 5468
rect 111820 5466 111876 5468
rect 111900 5466 111956 5468
rect 111980 5466 112036 5468
rect 111740 5414 111786 5466
rect 111786 5414 111796 5466
rect 111820 5414 111850 5466
rect 111850 5414 111862 5466
rect 111862 5414 111876 5466
rect 111900 5414 111914 5466
rect 111914 5414 111926 5466
rect 111926 5414 111956 5466
rect 111980 5414 111990 5466
rect 111990 5414 112036 5466
rect 111740 5412 111796 5414
rect 111820 5412 111876 5414
rect 111900 5412 111956 5414
rect 111980 5412 112036 5414
rect 111740 4378 111796 4380
rect 111820 4378 111876 4380
rect 111900 4378 111956 4380
rect 111980 4378 112036 4380
rect 111740 4326 111786 4378
rect 111786 4326 111796 4378
rect 111820 4326 111850 4378
rect 111850 4326 111862 4378
rect 111862 4326 111876 4378
rect 111900 4326 111914 4378
rect 111914 4326 111926 4378
rect 111926 4326 111956 4378
rect 111980 4326 111990 4378
rect 111990 4326 112036 4378
rect 111740 4324 111796 4326
rect 111820 4324 111876 4326
rect 111900 4324 111956 4326
rect 111980 4324 112036 4326
rect 111740 3290 111796 3292
rect 111820 3290 111876 3292
rect 111900 3290 111956 3292
rect 111980 3290 112036 3292
rect 111740 3238 111786 3290
rect 111786 3238 111796 3290
rect 111820 3238 111850 3290
rect 111850 3238 111862 3290
rect 111862 3238 111876 3290
rect 111900 3238 111914 3290
rect 111914 3238 111926 3290
rect 111926 3238 111956 3290
rect 111980 3238 111990 3290
rect 111990 3238 112036 3290
rect 111740 3236 111796 3238
rect 111820 3236 111876 3238
rect 111900 3236 111956 3238
rect 111980 3236 112036 3238
rect 127100 37562 127156 37564
rect 127180 37562 127236 37564
rect 127260 37562 127316 37564
rect 127340 37562 127396 37564
rect 127100 37510 127146 37562
rect 127146 37510 127156 37562
rect 127180 37510 127210 37562
rect 127210 37510 127222 37562
rect 127222 37510 127236 37562
rect 127260 37510 127274 37562
rect 127274 37510 127286 37562
rect 127286 37510 127316 37562
rect 127340 37510 127350 37562
rect 127350 37510 127396 37562
rect 127100 37508 127156 37510
rect 127180 37508 127236 37510
rect 127260 37508 127316 37510
rect 127340 37508 127396 37510
rect 128358 36760 128414 36816
rect 124218 36236 124274 36272
rect 124218 36216 124220 36236
rect 124220 36216 124272 36236
rect 124272 36216 124274 36236
rect 127100 36474 127156 36476
rect 127180 36474 127236 36476
rect 127260 36474 127316 36476
rect 127340 36474 127396 36476
rect 127100 36422 127146 36474
rect 127146 36422 127156 36474
rect 127180 36422 127210 36474
rect 127210 36422 127222 36474
rect 127222 36422 127236 36474
rect 127260 36422 127274 36474
rect 127274 36422 127286 36474
rect 127286 36422 127316 36474
rect 127340 36422 127350 36474
rect 127350 36422 127396 36474
rect 127100 36420 127156 36422
rect 127180 36420 127236 36422
rect 127260 36420 127316 36422
rect 127340 36420 127396 36422
rect 127100 35386 127156 35388
rect 127180 35386 127236 35388
rect 127260 35386 127316 35388
rect 127340 35386 127396 35388
rect 127100 35334 127146 35386
rect 127146 35334 127156 35386
rect 127180 35334 127210 35386
rect 127210 35334 127222 35386
rect 127222 35334 127236 35386
rect 127260 35334 127274 35386
rect 127274 35334 127286 35386
rect 127286 35334 127316 35386
rect 127340 35334 127350 35386
rect 127350 35334 127396 35386
rect 127100 35332 127156 35334
rect 127180 35332 127236 35334
rect 127260 35332 127316 35334
rect 127340 35332 127396 35334
rect 129554 36624 129610 36680
rect 132866 37168 132922 37224
rect 131670 36216 131726 36272
rect 129278 34992 129334 35048
rect 127100 34298 127156 34300
rect 127180 34298 127236 34300
rect 127260 34298 127316 34300
rect 127340 34298 127396 34300
rect 127100 34246 127146 34298
rect 127146 34246 127156 34298
rect 127180 34246 127210 34298
rect 127210 34246 127222 34298
rect 127222 34246 127236 34298
rect 127260 34246 127274 34298
rect 127274 34246 127286 34298
rect 127286 34246 127316 34298
rect 127340 34246 127350 34298
rect 127350 34246 127396 34298
rect 127100 34244 127156 34246
rect 127180 34244 127236 34246
rect 127260 34244 127316 34246
rect 127340 34244 127396 34246
rect 127100 33210 127156 33212
rect 127180 33210 127236 33212
rect 127260 33210 127316 33212
rect 127340 33210 127396 33212
rect 127100 33158 127146 33210
rect 127146 33158 127156 33210
rect 127180 33158 127210 33210
rect 127210 33158 127222 33210
rect 127222 33158 127236 33210
rect 127260 33158 127274 33210
rect 127274 33158 127286 33210
rect 127286 33158 127316 33210
rect 127340 33158 127350 33210
rect 127350 33158 127396 33210
rect 127100 33156 127156 33158
rect 127180 33156 127236 33158
rect 127260 33156 127316 33158
rect 127340 33156 127396 33158
rect 127100 32122 127156 32124
rect 127180 32122 127236 32124
rect 127260 32122 127316 32124
rect 127340 32122 127396 32124
rect 127100 32070 127146 32122
rect 127146 32070 127156 32122
rect 127180 32070 127210 32122
rect 127210 32070 127222 32122
rect 127222 32070 127236 32122
rect 127260 32070 127274 32122
rect 127274 32070 127286 32122
rect 127286 32070 127316 32122
rect 127340 32070 127350 32122
rect 127350 32070 127396 32122
rect 127100 32068 127156 32070
rect 127180 32068 127236 32070
rect 127260 32068 127316 32070
rect 127340 32068 127396 32070
rect 127100 31034 127156 31036
rect 127180 31034 127236 31036
rect 127260 31034 127316 31036
rect 127340 31034 127396 31036
rect 127100 30982 127146 31034
rect 127146 30982 127156 31034
rect 127180 30982 127210 31034
rect 127210 30982 127222 31034
rect 127222 30982 127236 31034
rect 127260 30982 127274 31034
rect 127274 30982 127286 31034
rect 127286 30982 127316 31034
rect 127340 30982 127350 31034
rect 127350 30982 127396 31034
rect 127100 30980 127156 30982
rect 127180 30980 127236 30982
rect 127260 30980 127316 30982
rect 127340 30980 127396 30982
rect 127100 29946 127156 29948
rect 127180 29946 127236 29948
rect 127260 29946 127316 29948
rect 127340 29946 127396 29948
rect 127100 29894 127146 29946
rect 127146 29894 127156 29946
rect 127180 29894 127210 29946
rect 127210 29894 127222 29946
rect 127222 29894 127236 29946
rect 127260 29894 127274 29946
rect 127274 29894 127286 29946
rect 127286 29894 127316 29946
rect 127340 29894 127350 29946
rect 127350 29894 127396 29946
rect 127100 29892 127156 29894
rect 127180 29892 127236 29894
rect 127260 29892 127316 29894
rect 127340 29892 127396 29894
rect 127100 28858 127156 28860
rect 127180 28858 127236 28860
rect 127260 28858 127316 28860
rect 127340 28858 127396 28860
rect 127100 28806 127146 28858
rect 127146 28806 127156 28858
rect 127180 28806 127210 28858
rect 127210 28806 127222 28858
rect 127222 28806 127236 28858
rect 127260 28806 127274 28858
rect 127274 28806 127286 28858
rect 127286 28806 127316 28858
rect 127340 28806 127350 28858
rect 127350 28806 127396 28858
rect 127100 28804 127156 28806
rect 127180 28804 127236 28806
rect 127260 28804 127316 28806
rect 127340 28804 127396 28806
rect 127100 27770 127156 27772
rect 127180 27770 127236 27772
rect 127260 27770 127316 27772
rect 127340 27770 127396 27772
rect 127100 27718 127146 27770
rect 127146 27718 127156 27770
rect 127180 27718 127210 27770
rect 127210 27718 127222 27770
rect 127222 27718 127236 27770
rect 127260 27718 127274 27770
rect 127274 27718 127286 27770
rect 127286 27718 127316 27770
rect 127340 27718 127350 27770
rect 127350 27718 127396 27770
rect 127100 27716 127156 27718
rect 127180 27716 127236 27718
rect 127260 27716 127316 27718
rect 127340 27716 127396 27718
rect 127100 26682 127156 26684
rect 127180 26682 127236 26684
rect 127260 26682 127316 26684
rect 127340 26682 127396 26684
rect 127100 26630 127146 26682
rect 127146 26630 127156 26682
rect 127180 26630 127210 26682
rect 127210 26630 127222 26682
rect 127222 26630 127236 26682
rect 127260 26630 127274 26682
rect 127274 26630 127286 26682
rect 127286 26630 127316 26682
rect 127340 26630 127350 26682
rect 127350 26630 127396 26682
rect 127100 26628 127156 26630
rect 127180 26628 127236 26630
rect 127260 26628 127316 26630
rect 127340 26628 127396 26630
rect 127100 25594 127156 25596
rect 127180 25594 127236 25596
rect 127260 25594 127316 25596
rect 127340 25594 127396 25596
rect 127100 25542 127146 25594
rect 127146 25542 127156 25594
rect 127180 25542 127210 25594
rect 127210 25542 127222 25594
rect 127222 25542 127236 25594
rect 127260 25542 127274 25594
rect 127274 25542 127286 25594
rect 127286 25542 127316 25594
rect 127340 25542 127350 25594
rect 127350 25542 127396 25594
rect 127100 25540 127156 25542
rect 127180 25540 127236 25542
rect 127260 25540 127316 25542
rect 127340 25540 127396 25542
rect 127100 24506 127156 24508
rect 127180 24506 127236 24508
rect 127260 24506 127316 24508
rect 127340 24506 127396 24508
rect 127100 24454 127146 24506
rect 127146 24454 127156 24506
rect 127180 24454 127210 24506
rect 127210 24454 127222 24506
rect 127222 24454 127236 24506
rect 127260 24454 127274 24506
rect 127274 24454 127286 24506
rect 127286 24454 127316 24506
rect 127340 24454 127350 24506
rect 127350 24454 127396 24506
rect 127100 24452 127156 24454
rect 127180 24452 127236 24454
rect 127260 24452 127316 24454
rect 127340 24452 127396 24454
rect 127100 23418 127156 23420
rect 127180 23418 127236 23420
rect 127260 23418 127316 23420
rect 127340 23418 127396 23420
rect 127100 23366 127146 23418
rect 127146 23366 127156 23418
rect 127180 23366 127210 23418
rect 127210 23366 127222 23418
rect 127222 23366 127236 23418
rect 127260 23366 127274 23418
rect 127274 23366 127286 23418
rect 127286 23366 127316 23418
rect 127340 23366 127350 23418
rect 127350 23366 127396 23418
rect 127100 23364 127156 23366
rect 127180 23364 127236 23366
rect 127260 23364 127316 23366
rect 127340 23364 127396 23366
rect 127100 22330 127156 22332
rect 127180 22330 127236 22332
rect 127260 22330 127316 22332
rect 127340 22330 127396 22332
rect 127100 22278 127146 22330
rect 127146 22278 127156 22330
rect 127180 22278 127210 22330
rect 127210 22278 127222 22330
rect 127222 22278 127236 22330
rect 127260 22278 127274 22330
rect 127274 22278 127286 22330
rect 127286 22278 127316 22330
rect 127340 22278 127350 22330
rect 127350 22278 127396 22330
rect 127100 22276 127156 22278
rect 127180 22276 127236 22278
rect 127260 22276 127316 22278
rect 127340 22276 127396 22278
rect 127100 21242 127156 21244
rect 127180 21242 127236 21244
rect 127260 21242 127316 21244
rect 127340 21242 127396 21244
rect 127100 21190 127146 21242
rect 127146 21190 127156 21242
rect 127180 21190 127210 21242
rect 127210 21190 127222 21242
rect 127222 21190 127236 21242
rect 127260 21190 127274 21242
rect 127274 21190 127286 21242
rect 127286 21190 127316 21242
rect 127340 21190 127350 21242
rect 127350 21190 127396 21242
rect 127100 21188 127156 21190
rect 127180 21188 127236 21190
rect 127260 21188 127316 21190
rect 127340 21188 127396 21190
rect 127100 20154 127156 20156
rect 127180 20154 127236 20156
rect 127260 20154 127316 20156
rect 127340 20154 127396 20156
rect 127100 20102 127146 20154
rect 127146 20102 127156 20154
rect 127180 20102 127210 20154
rect 127210 20102 127222 20154
rect 127222 20102 127236 20154
rect 127260 20102 127274 20154
rect 127274 20102 127286 20154
rect 127286 20102 127316 20154
rect 127340 20102 127350 20154
rect 127350 20102 127396 20154
rect 127100 20100 127156 20102
rect 127180 20100 127236 20102
rect 127260 20100 127316 20102
rect 127340 20100 127396 20102
rect 127100 19066 127156 19068
rect 127180 19066 127236 19068
rect 127260 19066 127316 19068
rect 127340 19066 127396 19068
rect 127100 19014 127146 19066
rect 127146 19014 127156 19066
rect 127180 19014 127210 19066
rect 127210 19014 127222 19066
rect 127222 19014 127236 19066
rect 127260 19014 127274 19066
rect 127274 19014 127286 19066
rect 127286 19014 127316 19066
rect 127340 19014 127350 19066
rect 127350 19014 127396 19066
rect 127100 19012 127156 19014
rect 127180 19012 127236 19014
rect 127260 19012 127316 19014
rect 127340 19012 127396 19014
rect 127100 17978 127156 17980
rect 127180 17978 127236 17980
rect 127260 17978 127316 17980
rect 127340 17978 127396 17980
rect 127100 17926 127146 17978
rect 127146 17926 127156 17978
rect 127180 17926 127210 17978
rect 127210 17926 127222 17978
rect 127222 17926 127236 17978
rect 127260 17926 127274 17978
rect 127274 17926 127286 17978
rect 127286 17926 127316 17978
rect 127340 17926 127350 17978
rect 127350 17926 127396 17978
rect 127100 17924 127156 17926
rect 127180 17924 127236 17926
rect 127260 17924 127316 17926
rect 127340 17924 127396 17926
rect 127100 16890 127156 16892
rect 127180 16890 127236 16892
rect 127260 16890 127316 16892
rect 127340 16890 127396 16892
rect 127100 16838 127146 16890
rect 127146 16838 127156 16890
rect 127180 16838 127210 16890
rect 127210 16838 127222 16890
rect 127222 16838 127236 16890
rect 127260 16838 127274 16890
rect 127274 16838 127286 16890
rect 127286 16838 127316 16890
rect 127340 16838 127350 16890
rect 127350 16838 127396 16890
rect 127100 16836 127156 16838
rect 127180 16836 127236 16838
rect 127260 16836 127316 16838
rect 127340 16836 127396 16838
rect 127100 15802 127156 15804
rect 127180 15802 127236 15804
rect 127260 15802 127316 15804
rect 127340 15802 127396 15804
rect 127100 15750 127146 15802
rect 127146 15750 127156 15802
rect 127180 15750 127210 15802
rect 127210 15750 127222 15802
rect 127222 15750 127236 15802
rect 127260 15750 127274 15802
rect 127274 15750 127286 15802
rect 127286 15750 127316 15802
rect 127340 15750 127350 15802
rect 127350 15750 127396 15802
rect 127100 15748 127156 15750
rect 127180 15748 127236 15750
rect 127260 15748 127316 15750
rect 127340 15748 127396 15750
rect 127100 14714 127156 14716
rect 127180 14714 127236 14716
rect 127260 14714 127316 14716
rect 127340 14714 127396 14716
rect 127100 14662 127146 14714
rect 127146 14662 127156 14714
rect 127180 14662 127210 14714
rect 127210 14662 127222 14714
rect 127222 14662 127236 14714
rect 127260 14662 127274 14714
rect 127274 14662 127286 14714
rect 127286 14662 127316 14714
rect 127340 14662 127350 14714
rect 127350 14662 127396 14714
rect 127100 14660 127156 14662
rect 127180 14660 127236 14662
rect 127260 14660 127316 14662
rect 127340 14660 127396 14662
rect 127100 13626 127156 13628
rect 127180 13626 127236 13628
rect 127260 13626 127316 13628
rect 127340 13626 127396 13628
rect 127100 13574 127146 13626
rect 127146 13574 127156 13626
rect 127180 13574 127210 13626
rect 127210 13574 127222 13626
rect 127222 13574 127236 13626
rect 127260 13574 127274 13626
rect 127274 13574 127286 13626
rect 127286 13574 127316 13626
rect 127340 13574 127350 13626
rect 127350 13574 127396 13626
rect 127100 13572 127156 13574
rect 127180 13572 127236 13574
rect 127260 13572 127316 13574
rect 127340 13572 127396 13574
rect 127100 12538 127156 12540
rect 127180 12538 127236 12540
rect 127260 12538 127316 12540
rect 127340 12538 127396 12540
rect 127100 12486 127146 12538
rect 127146 12486 127156 12538
rect 127180 12486 127210 12538
rect 127210 12486 127222 12538
rect 127222 12486 127236 12538
rect 127260 12486 127274 12538
rect 127274 12486 127286 12538
rect 127286 12486 127316 12538
rect 127340 12486 127350 12538
rect 127350 12486 127396 12538
rect 127100 12484 127156 12486
rect 127180 12484 127236 12486
rect 127260 12484 127316 12486
rect 127340 12484 127396 12486
rect 127100 11450 127156 11452
rect 127180 11450 127236 11452
rect 127260 11450 127316 11452
rect 127340 11450 127396 11452
rect 127100 11398 127146 11450
rect 127146 11398 127156 11450
rect 127180 11398 127210 11450
rect 127210 11398 127222 11450
rect 127222 11398 127236 11450
rect 127260 11398 127274 11450
rect 127274 11398 127286 11450
rect 127286 11398 127316 11450
rect 127340 11398 127350 11450
rect 127350 11398 127396 11450
rect 127100 11396 127156 11398
rect 127180 11396 127236 11398
rect 127260 11396 127316 11398
rect 127340 11396 127396 11398
rect 127100 10362 127156 10364
rect 127180 10362 127236 10364
rect 127260 10362 127316 10364
rect 127340 10362 127396 10364
rect 127100 10310 127146 10362
rect 127146 10310 127156 10362
rect 127180 10310 127210 10362
rect 127210 10310 127222 10362
rect 127222 10310 127236 10362
rect 127260 10310 127274 10362
rect 127274 10310 127286 10362
rect 127286 10310 127316 10362
rect 127340 10310 127350 10362
rect 127350 10310 127396 10362
rect 127100 10308 127156 10310
rect 127180 10308 127236 10310
rect 127260 10308 127316 10310
rect 127340 10308 127396 10310
rect 134522 35128 134578 35184
rect 127100 9274 127156 9276
rect 127180 9274 127236 9276
rect 127260 9274 127316 9276
rect 127340 9274 127396 9276
rect 127100 9222 127146 9274
rect 127146 9222 127156 9274
rect 127180 9222 127210 9274
rect 127210 9222 127222 9274
rect 127222 9222 127236 9274
rect 127260 9222 127274 9274
rect 127274 9222 127286 9274
rect 127286 9222 127316 9274
rect 127340 9222 127350 9274
rect 127350 9222 127396 9274
rect 127100 9220 127156 9222
rect 127180 9220 127236 9222
rect 127260 9220 127316 9222
rect 127340 9220 127396 9222
rect 127100 8186 127156 8188
rect 127180 8186 127236 8188
rect 127260 8186 127316 8188
rect 127340 8186 127396 8188
rect 127100 8134 127146 8186
rect 127146 8134 127156 8186
rect 127180 8134 127210 8186
rect 127210 8134 127222 8186
rect 127222 8134 127236 8186
rect 127260 8134 127274 8186
rect 127274 8134 127286 8186
rect 127286 8134 127316 8186
rect 127340 8134 127350 8186
rect 127350 8134 127396 8186
rect 127100 8132 127156 8134
rect 127180 8132 127236 8134
rect 127260 8132 127316 8134
rect 127340 8132 127396 8134
rect 127100 7098 127156 7100
rect 127180 7098 127236 7100
rect 127260 7098 127316 7100
rect 127340 7098 127396 7100
rect 127100 7046 127146 7098
rect 127146 7046 127156 7098
rect 127180 7046 127210 7098
rect 127210 7046 127222 7098
rect 127222 7046 127236 7098
rect 127260 7046 127274 7098
rect 127274 7046 127286 7098
rect 127286 7046 127316 7098
rect 127340 7046 127350 7098
rect 127350 7046 127396 7098
rect 127100 7044 127156 7046
rect 127180 7044 127236 7046
rect 127260 7044 127316 7046
rect 127340 7044 127396 7046
rect 127100 6010 127156 6012
rect 127180 6010 127236 6012
rect 127260 6010 127316 6012
rect 127340 6010 127396 6012
rect 127100 5958 127146 6010
rect 127146 5958 127156 6010
rect 127180 5958 127210 6010
rect 127210 5958 127222 6010
rect 127222 5958 127236 6010
rect 127260 5958 127274 6010
rect 127274 5958 127286 6010
rect 127286 5958 127316 6010
rect 127340 5958 127350 6010
rect 127350 5958 127396 6010
rect 127100 5956 127156 5958
rect 127180 5956 127236 5958
rect 127260 5956 127316 5958
rect 127340 5956 127396 5958
rect 127100 4922 127156 4924
rect 127180 4922 127236 4924
rect 127260 4922 127316 4924
rect 127340 4922 127396 4924
rect 127100 4870 127146 4922
rect 127146 4870 127156 4922
rect 127180 4870 127210 4922
rect 127210 4870 127222 4922
rect 127222 4870 127236 4922
rect 127260 4870 127274 4922
rect 127274 4870 127286 4922
rect 127286 4870 127316 4922
rect 127340 4870 127350 4922
rect 127350 4870 127396 4922
rect 127100 4868 127156 4870
rect 127180 4868 127236 4870
rect 127260 4868 127316 4870
rect 127340 4868 127396 4870
rect 127100 3834 127156 3836
rect 127180 3834 127236 3836
rect 127260 3834 127316 3836
rect 127340 3834 127396 3836
rect 127100 3782 127146 3834
rect 127146 3782 127156 3834
rect 127180 3782 127210 3834
rect 127210 3782 127222 3834
rect 127222 3782 127236 3834
rect 127260 3782 127274 3834
rect 127274 3782 127286 3834
rect 127286 3782 127316 3834
rect 127340 3782 127350 3834
rect 127350 3782 127396 3834
rect 127100 3780 127156 3782
rect 127180 3780 127236 3782
rect 127260 3780 127316 3782
rect 127340 3780 127396 3782
rect 127100 2746 127156 2748
rect 127180 2746 127236 2748
rect 127260 2746 127316 2748
rect 127340 2746 127396 2748
rect 127100 2694 127146 2746
rect 127146 2694 127156 2746
rect 127180 2694 127210 2746
rect 127210 2694 127222 2746
rect 127222 2694 127236 2746
rect 127260 2694 127274 2746
rect 127274 2694 127286 2746
rect 127286 2694 127316 2746
rect 127340 2694 127350 2746
rect 127350 2694 127396 2746
rect 127100 2692 127156 2694
rect 127180 2692 127236 2694
rect 127260 2692 127316 2694
rect 127340 2692 127396 2694
rect 111740 2202 111796 2204
rect 111820 2202 111876 2204
rect 111900 2202 111956 2204
rect 111980 2202 112036 2204
rect 111740 2150 111786 2202
rect 111786 2150 111796 2202
rect 111820 2150 111850 2202
rect 111850 2150 111862 2202
rect 111862 2150 111876 2202
rect 111900 2150 111914 2202
rect 111914 2150 111926 2202
rect 111926 2150 111956 2202
rect 111980 2150 111990 2202
rect 111990 2150 112036 2202
rect 111740 2148 111796 2150
rect 111820 2148 111876 2150
rect 111900 2148 111956 2150
rect 111980 2148 112036 2150
rect 142460 37018 142516 37020
rect 142540 37018 142596 37020
rect 142620 37018 142676 37020
rect 142700 37018 142756 37020
rect 142460 36966 142506 37018
rect 142506 36966 142516 37018
rect 142540 36966 142570 37018
rect 142570 36966 142582 37018
rect 142582 36966 142596 37018
rect 142620 36966 142634 37018
rect 142634 36966 142646 37018
rect 142646 36966 142676 37018
rect 142700 36966 142710 37018
rect 142710 36966 142756 37018
rect 142460 36964 142516 36966
rect 142540 36964 142596 36966
rect 142620 36964 142676 36966
rect 142700 36964 142756 36966
rect 142460 35930 142516 35932
rect 142540 35930 142596 35932
rect 142620 35930 142676 35932
rect 142700 35930 142756 35932
rect 142460 35878 142506 35930
rect 142506 35878 142516 35930
rect 142540 35878 142570 35930
rect 142570 35878 142582 35930
rect 142582 35878 142596 35930
rect 142620 35878 142634 35930
rect 142634 35878 142646 35930
rect 142646 35878 142676 35930
rect 142700 35878 142710 35930
rect 142710 35878 142756 35930
rect 142460 35876 142516 35878
rect 142540 35876 142596 35878
rect 142620 35876 142676 35878
rect 142700 35876 142756 35878
rect 142460 34842 142516 34844
rect 142540 34842 142596 34844
rect 142620 34842 142676 34844
rect 142700 34842 142756 34844
rect 142460 34790 142506 34842
rect 142506 34790 142516 34842
rect 142540 34790 142570 34842
rect 142570 34790 142582 34842
rect 142582 34790 142596 34842
rect 142620 34790 142634 34842
rect 142634 34790 142646 34842
rect 142646 34790 142676 34842
rect 142700 34790 142710 34842
rect 142710 34790 142756 34842
rect 142460 34788 142516 34790
rect 142540 34788 142596 34790
rect 142620 34788 142676 34790
rect 142700 34788 142756 34790
rect 142460 33754 142516 33756
rect 142540 33754 142596 33756
rect 142620 33754 142676 33756
rect 142700 33754 142756 33756
rect 142460 33702 142506 33754
rect 142506 33702 142516 33754
rect 142540 33702 142570 33754
rect 142570 33702 142582 33754
rect 142582 33702 142596 33754
rect 142620 33702 142634 33754
rect 142634 33702 142646 33754
rect 142646 33702 142676 33754
rect 142700 33702 142710 33754
rect 142710 33702 142756 33754
rect 142460 33700 142516 33702
rect 142540 33700 142596 33702
rect 142620 33700 142676 33702
rect 142700 33700 142756 33702
rect 142460 32666 142516 32668
rect 142540 32666 142596 32668
rect 142620 32666 142676 32668
rect 142700 32666 142756 32668
rect 142460 32614 142506 32666
rect 142506 32614 142516 32666
rect 142540 32614 142570 32666
rect 142570 32614 142582 32666
rect 142582 32614 142596 32666
rect 142620 32614 142634 32666
rect 142634 32614 142646 32666
rect 142646 32614 142676 32666
rect 142700 32614 142710 32666
rect 142710 32614 142756 32666
rect 142460 32612 142516 32614
rect 142540 32612 142596 32614
rect 142620 32612 142676 32614
rect 142700 32612 142756 32614
rect 142460 31578 142516 31580
rect 142540 31578 142596 31580
rect 142620 31578 142676 31580
rect 142700 31578 142756 31580
rect 142460 31526 142506 31578
rect 142506 31526 142516 31578
rect 142540 31526 142570 31578
rect 142570 31526 142582 31578
rect 142582 31526 142596 31578
rect 142620 31526 142634 31578
rect 142634 31526 142646 31578
rect 142646 31526 142676 31578
rect 142700 31526 142710 31578
rect 142710 31526 142756 31578
rect 142460 31524 142516 31526
rect 142540 31524 142596 31526
rect 142620 31524 142676 31526
rect 142700 31524 142756 31526
rect 142460 30490 142516 30492
rect 142540 30490 142596 30492
rect 142620 30490 142676 30492
rect 142700 30490 142756 30492
rect 142460 30438 142506 30490
rect 142506 30438 142516 30490
rect 142540 30438 142570 30490
rect 142570 30438 142582 30490
rect 142582 30438 142596 30490
rect 142620 30438 142634 30490
rect 142634 30438 142646 30490
rect 142646 30438 142676 30490
rect 142700 30438 142710 30490
rect 142710 30438 142756 30490
rect 142460 30436 142516 30438
rect 142540 30436 142596 30438
rect 142620 30436 142676 30438
rect 142700 30436 142756 30438
rect 142460 29402 142516 29404
rect 142540 29402 142596 29404
rect 142620 29402 142676 29404
rect 142700 29402 142756 29404
rect 142460 29350 142506 29402
rect 142506 29350 142516 29402
rect 142540 29350 142570 29402
rect 142570 29350 142582 29402
rect 142582 29350 142596 29402
rect 142620 29350 142634 29402
rect 142634 29350 142646 29402
rect 142646 29350 142676 29402
rect 142700 29350 142710 29402
rect 142710 29350 142756 29402
rect 142460 29348 142516 29350
rect 142540 29348 142596 29350
rect 142620 29348 142676 29350
rect 142700 29348 142756 29350
rect 142460 28314 142516 28316
rect 142540 28314 142596 28316
rect 142620 28314 142676 28316
rect 142700 28314 142756 28316
rect 142460 28262 142506 28314
rect 142506 28262 142516 28314
rect 142540 28262 142570 28314
rect 142570 28262 142582 28314
rect 142582 28262 142596 28314
rect 142620 28262 142634 28314
rect 142634 28262 142646 28314
rect 142646 28262 142676 28314
rect 142700 28262 142710 28314
rect 142710 28262 142756 28314
rect 142460 28260 142516 28262
rect 142540 28260 142596 28262
rect 142620 28260 142676 28262
rect 142700 28260 142756 28262
rect 142460 27226 142516 27228
rect 142540 27226 142596 27228
rect 142620 27226 142676 27228
rect 142700 27226 142756 27228
rect 142460 27174 142506 27226
rect 142506 27174 142516 27226
rect 142540 27174 142570 27226
rect 142570 27174 142582 27226
rect 142582 27174 142596 27226
rect 142620 27174 142634 27226
rect 142634 27174 142646 27226
rect 142646 27174 142676 27226
rect 142700 27174 142710 27226
rect 142710 27174 142756 27226
rect 142460 27172 142516 27174
rect 142540 27172 142596 27174
rect 142620 27172 142676 27174
rect 142700 27172 142756 27174
rect 142460 26138 142516 26140
rect 142540 26138 142596 26140
rect 142620 26138 142676 26140
rect 142700 26138 142756 26140
rect 142460 26086 142506 26138
rect 142506 26086 142516 26138
rect 142540 26086 142570 26138
rect 142570 26086 142582 26138
rect 142582 26086 142596 26138
rect 142620 26086 142634 26138
rect 142634 26086 142646 26138
rect 142646 26086 142676 26138
rect 142700 26086 142710 26138
rect 142710 26086 142756 26138
rect 142460 26084 142516 26086
rect 142540 26084 142596 26086
rect 142620 26084 142676 26086
rect 142700 26084 142756 26086
rect 142460 25050 142516 25052
rect 142540 25050 142596 25052
rect 142620 25050 142676 25052
rect 142700 25050 142756 25052
rect 142460 24998 142506 25050
rect 142506 24998 142516 25050
rect 142540 24998 142570 25050
rect 142570 24998 142582 25050
rect 142582 24998 142596 25050
rect 142620 24998 142634 25050
rect 142634 24998 142646 25050
rect 142646 24998 142676 25050
rect 142700 24998 142710 25050
rect 142710 24998 142756 25050
rect 142460 24996 142516 24998
rect 142540 24996 142596 24998
rect 142620 24996 142676 24998
rect 142700 24996 142756 24998
rect 142460 23962 142516 23964
rect 142540 23962 142596 23964
rect 142620 23962 142676 23964
rect 142700 23962 142756 23964
rect 142460 23910 142506 23962
rect 142506 23910 142516 23962
rect 142540 23910 142570 23962
rect 142570 23910 142582 23962
rect 142582 23910 142596 23962
rect 142620 23910 142634 23962
rect 142634 23910 142646 23962
rect 142646 23910 142676 23962
rect 142700 23910 142710 23962
rect 142710 23910 142756 23962
rect 142460 23908 142516 23910
rect 142540 23908 142596 23910
rect 142620 23908 142676 23910
rect 142700 23908 142756 23910
rect 142460 22874 142516 22876
rect 142540 22874 142596 22876
rect 142620 22874 142676 22876
rect 142700 22874 142756 22876
rect 142460 22822 142506 22874
rect 142506 22822 142516 22874
rect 142540 22822 142570 22874
rect 142570 22822 142582 22874
rect 142582 22822 142596 22874
rect 142620 22822 142634 22874
rect 142634 22822 142646 22874
rect 142646 22822 142676 22874
rect 142700 22822 142710 22874
rect 142710 22822 142756 22874
rect 142460 22820 142516 22822
rect 142540 22820 142596 22822
rect 142620 22820 142676 22822
rect 142700 22820 142756 22822
rect 142460 21786 142516 21788
rect 142540 21786 142596 21788
rect 142620 21786 142676 21788
rect 142700 21786 142756 21788
rect 142460 21734 142506 21786
rect 142506 21734 142516 21786
rect 142540 21734 142570 21786
rect 142570 21734 142582 21786
rect 142582 21734 142596 21786
rect 142620 21734 142634 21786
rect 142634 21734 142646 21786
rect 142646 21734 142676 21786
rect 142700 21734 142710 21786
rect 142710 21734 142756 21786
rect 142460 21732 142516 21734
rect 142540 21732 142596 21734
rect 142620 21732 142676 21734
rect 142700 21732 142756 21734
rect 142460 20698 142516 20700
rect 142540 20698 142596 20700
rect 142620 20698 142676 20700
rect 142700 20698 142756 20700
rect 142460 20646 142506 20698
rect 142506 20646 142516 20698
rect 142540 20646 142570 20698
rect 142570 20646 142582 20698
rect 142582 20646 142596 20698
rect 142620 20646 142634 20698
rect 142634 20646 142646 20698
rect 142646 20646 142676 20698
rect 142700 20646 142710 20698
rect 142710 20646 142756 20698
rect 142460 20644 142516 20646
rect 142540 20644 142596 20646
rect 142620 20644 142676 20646
rect 142700 20644 142756 20646
rect 142460 19610 142516 19612
rect 142540 19610 142596 19612
rect 142620 19610 142676 19612
rect 142700 19610 142756 19612
rect 142460 19558 142506 19610
rect 142506 19558 142516 19610
rect 142540 19558 142570 19610
rect 142570 19558 142582 19610
rect 142582 19558 142596 19610
rect 142620 19558 142634 19610
rect 142634 19558 142646 19610
rect 142646 19558 142676 19610
rect 142700 19558 142710 19610
rect 142710 19558 142756 19610
rect 142460 19556 142516 19558
rect 142540 19556 142596 19558
rect 142620 19556 142676 19558
rect 142700 19556 142756 19558
rect 142460 18522 142516 18524
rect 142540 18522 142596 18524
rect 142620 18522 142676 18524
rect 142700 18522 142756 18524
rect 142460 18470 142506 18522
rect 142506 18470 142516 18522
rect 142540 18470 142570 18522
rect 142570 18470 142582 18522
rect 142582 18470 142596 18522
rect 142620 18470 142634 18522
rect 142634 18470 142646 18522
rect 142646 18470 142676 18522
rect 142700 18470 142710 18522
rect 142710 18470 142756 18522
rect 142460 18468 142516 18470
rect 142540 18468 142596 18470
rect 142620 18468 142676 18470
rect 142700 18468 142756 18470
rect 142460 17434 142516 17436
rect 142540 17434 142596 17436
rect 142620 17434 142676 17436
rect 142700 17434 142756 17436
rect 142460 17382 142506 17434
rect 142506 17382 142516 17434
rect 142540 17382 142570 17434
rect 142570 17382 142582 17434
rect 142582 17382 142596 17434
rect 142620 17382 142634 17434
rect 142634 17382 142646 17434
rect 142646 17382 142676 17434
rect 142700 17382 142710 17434
rect 142710 17382 142756 17434
rect 142460 17380 142516 17382
rect 142540 17380 142596 17382
rect 142620 17380 142676 17382
rect 142700 17380 142756 17382
rect 142460 16346 142516 16348
rect 142540 16346 142596 16348
rect 142620 16346 142676 16348
rect 142700 16346 142756 16348
rect 142460 16294 142506 16346
rect 142506 16294 142516 16346
rect 142540 16294 142570 16346
rect 142570 16294 142582 16346
rect 142582 16294 142596 16346
rect 142620 16294 142634 16346
rect 142634 16294 142646 16346
rect 142646 16294 142676 16346
rect 142700 16294 142710 16346
rect 142710 16294 142756 16346
rect 142460 16292 142516 16294
rect 142540 16292 142596 16294
rect 142620 16292 142676 16294
rect 142700 16292 142756 16294
rect 142460 15258 142516 15260
rect 142540 15258 142596 15260
rect 142620 15258 142676 15260
rect 142700 15258 142756 15260
rect 142460 15206 142506 15258
rect 142506 15206 142516 15258
rect 142540 15206 142570 15258
rect 142570 15206 142582 15258
rect 142582 15206 142596 15258
rect 142620 15206 142634 15258
rect 142634 15206 142646 15258
rect 142646 15206 142676 15258
rect 142700 15206 142710 15258
rect 142710 15206 142756 15258
rect 142460 15204 142516 15206
rect 142540 15204 142596 15206
rect 142620 15204 142676 15206
rect 142700 15204 142756 15206
rect 142460 14170 142516 14172
rect 142540 14170 142596 14172
rect 142620 14170 142676 14172
rect 142700 14170 142756 14172
rect 142460 14118 142506 14170
rect 142506 14118 142516 14170
rect 142540 14118 142570 14170
rect 142570 14118 142582 14170
rect 142582 14118 142596 14170
rect 142620 14118 142634 14170
rect 142634 14118 142646 14170
rect 142646 14118 142676 14170
rect 142700 14118 142710 14170
rect 142710 14118 142756 14170
rect 142460 14116 142516 14118
rect 142540 14116 142596 14118
rect 142620 14116 142676 14118
rect 142700 14116 142756 14118
rect 142460 13082 142516 13084
rect 142540 13082 142596 13084
rect 142620 13082 142676 13084
rect 142700 13082 142756 13084
rect 142460 13030 142506 13082
rect 142506 13030 142516 13082
rect 142540 13030 142570 13082
rect 142570 13030 142582 13082
rect 142582 13030 142596 13082
rect 142620 13030 142634 13082
rect 142634 13030 142646 13082
rect 142646 13030 142676 13082
rect 142700 13030 142710 13082
rect 142710 13030 142756 13082
rect 142460 13028 142516 13030
rect 142540 13028 142596 13030
rect 142620 13028 142676 13030
rect 142700 13028 142756 13030
rect 142460 11994 142516 11996
rect 142540 11994 142596 11996
rect 142620 11994 142676 11996
rect 142700 11994 142756 11996
rect 142460 11942 142506 11994
rect 142506 11942 142516 11994
rect 142540 11942 142570 11994
rect 142570 11942 142582 11994
rect 142582 11942 142596 11994
rect 142620 11942 142634 11994
rect 142634 11942 142646 11994
rect 142646 11942 142676 11994
rect 142700 11942 142710 11994
rect 142710 11942 142756 11994
rect 142460 11940 142516 11942
rect 142540 11940 142596 11942
rect 142620 11940 142676 11942
rect 142700 11940 142756 11942
rect 142460 10906 142516 10908
rect 142540 10906 142596 10908
rect 142620 10906 142676 10908
rect 142700 10906 142756 10908
rect 142460 10854 142506 10906
rect 142506 10854 142516 10906
rect 142540 10854 142570 10906
rect 142570 10854 142582 10906
rect 142582 10854 142596 10906
rect 142620 10854 142634 10906
rect 142634 10854 142646 10906
rect 142646 10854 142676 10906
rect 142700 10854 142710 10906
rect 142710 10854 142756 10906
rect 142460 10852 142516 10854
rect 142540 10852 142596 10854
rect 142620 10852 142676 10854
rect 142700 10852 142756 10854
rect 142460 9818 142516 9820
rect 142540 9818 142596 9820
rect 142620 9818 142676 9820
rect 142700 9818 142756 9820
rect 142460 9766 142506 9818
rect 142506 9766 142516 9818
rect 142540 9766 142570 9818
rect 142570 9766 142582 9818
rect 142582 9766 142596 9818
rect 142620 9766 142634 9818
rect 142634 9766 142646 9818
rect 142646 9766 142676 9818
rect 142700 9766 142710 9818
rect 142710 9766 142756 9818
rect 142460 9764 142516 9766
rect 142540 9764 142596 9766
rect 142620 9764 142676 9766
rect 142700 9764 142756 9766
rect 142460 8730 142516 8732
rect 142540 8730 142596 8732
rect 142620 8730 142676 8732
rect 142700 8730 142756 8732
rect 142460 8678 142506 8730
rect 142506 8678 142516 8730
rect 142540 8678 142570 8730
rect 142570 8678 142582 8730
rect 142582 8678 142596 8730
rect 142620 8678 142634 8730
rect 142634 8678 142646 8730
rect 142646 8678 142676 8730
rect 142700 8678 142710 8730
rect 142710 8678 142756 8730
rect 142460 8676 142516 8678
rect 142540 8676 142596 8678
rect 142620 8676 142676 8678
rect 142700 8676 142756 8678
rect 142460 7642 142516 7644
rect 142540 7642 142596 7644
rect 142620 7642 142676 7644
rect 142700 7642 142756 7644
rect 142460 7590 142506 7642
rect 142506 7590 142516 7642
rect 142540 7590 142570 7642
rect 142570 7590 142582 7642
rect 142582 7590 142596 7642
rect 142620 7590 142634 7642
rect 142634 7590 142646 7642
rect 142646 7590 142676 7642
rect 142700 7590 142710 7642
rect 142710 7590 142756 7642
rect 142460 7588 142516 7590
rect 142540 7588 142596 7590
rect 142620 7588 142676 7590
rect 142700 7588 142756 7590
rect 142460 6554 142516 6556
rect 142540 6554 142596 6556
rect 142620 6554 142676 6556
rect 142700 6554 142756 6556
rect 142460 6502 142506 6554
rect 142506 6502 142516 6554
rect 142540 6502 142570 6554
rect 142570 6502 142582 6554
rect 142582 6502 142596 6554
rect 142620 6502 142634 6554
rect 142634 6502 142646 6554
rect 142646 6502 142676 6554
rect 142700 6502 142710 6554
rect 142710 6502 142756 6554
rect 142460 6500 142516 6502
rect 142540 6500 142596 6502
rect 142620 6500 142676 6502
rect 142700 6500 142756 6502
rect 142460 5466 142516 5468
rect 142540 5466 142596 5468
rect 142620 5466 142676 5468
rect 142700 5466 142756 5468
rect 142460 5414 142506 5466
rect 142506 5414 142516 5466
rect 142540 5414 142570 5466
rect 142570 5414 142582 5466
rect 142582 5414 142596 5466
rect 142620 5414 142634 5466
rect 142634 5414 142646 5466
rect 142646 5414 142676 5466
rect 142700 5414 142710 5466
rect 142710 5414 142756 5466
rect 142460 5412 142516 5414
rect 142540 5412 142596 5414
rect 142620 5412 142676 5414
rect 142700 5412 142756 5414
rect 142460 4378 142516 4380
rect 142540 4378 142596 4380
rect 142620 4378 142676 4380
rect 142700 4378 142756 4380
rect 142460 4326 142506 4378
rect 142506 4326 142516 4378
rect 142540 4326 142570 4378
rect 142570 4326 142582 4378
rect 142582 4326 142596 4378
rect 142620 4326 142634 4378
rect 142634 4326 142646 4378
rect 142646 4326 142676 4378
rect 142700 4326 142710 4378
rect 142710 4326 142756 4378
rect 142460 4324 142516 4326
rect 142540 4324 142596 4326
rect 142620 4324 142676 4326
rect 142700 4324 142756 4326
rect 142460 3290 142516 3292
rect 142540 3290 142596 3292
rect 142620 3290 142676 3292
rect 142700 3290 142756 3292
rect 142460 3238 142506 3290
rect 142506 3238 142516 3290
rect 142540 3238 142570 3290
rect 142570 3238 142582 3290
rect 142582 3238 142596 3290
rect 142620 3238 142634 3290
rect 142634 3238 142646 3290
rect 142646 3238 142676 3290
rect 142700 3238 142710 3290
rect 142710 3238 142756 3290
rect 142460 3236 142516 3238
rect 142540 3236 142596 3238
rect 142620 3236 142676 3238
rect 142700 3236 142756 3238
rect 142460 2202 142516 2204
rect 142540 2202 142596 2204
rect 142620 2202 142676 2204
rect 142700 2202 142756 2204
rect 142460 2150 142506 2202
rect 142506 2150 142516 2202
rect 142540 2150 142570 2202
rect 142570 2150 142582 2202
rect 142582 2150 142596 2202
rect 142620 2150 142634 2202
rect 142634 2150 142646 2202
rect 142646 2150 142676 2202
rect 142700 2150 142710 2202
rect 142710 2150 142756 2202
rect 142460 2148 142516 2150
rect 142540 2148 142596 2150
rect 142620 2148 142676 2150
rect 142700 2148 142756 2150
<< metal3 >>
rect 79501 37634 79567 37637
rect 85757 37634 85823 37637
rect 79501 37632 85823 37634
rect 79501 37576 79506 37632
rect 79562 37576 85762 37632
rect 85818 37576 85823 37632
rect 79501 37574 85823 37576
rect 79501 37571 79567 37574
rect 85757 37571 85823 37574
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 65650 37568 65966 37569
rect 65650 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65966 37568
rect 65650 37503 65966 37504
rect 96370 37568 96686 37569
rect 96370 37504 96376 37568
rect 96440 37504 96456 37568
rect 96520 37504 96536 37568
rect 96600 37504 96616 37568
rect 96680 37504 96686 37568
rect 96370 37503 96686 37504
rect 127090 37568 127406 37569
rect 127090 37504 127096 37568
rect 127160 37504 127176 37568
rect 127240 37504 127256 37568
rect 127320 37504 127336 37568
rect 127400 37504 127406 37568
rect 127090 37503 127406 37504
rect 20437 37498 20503 37501
rect 28165 37498 28231 37501
rect 20437 37496 28231 37498
rect 20437 37440 20442 37496
rect 20498 37440 28170 37496
rect 28226 37440 28231 37496
rect 20437 37438 28231 37440
rect 20437 37435 20503 37438
rect 28165 37435 28231 37438
rect 58341 37498 58407 37501
rect 59813 37498 59879 37501
rect 58341 37496 59879 37498
rect 58341 37440 58346 37496
rect 58402 37440 59818 37496
rect 59874 37440 59879 37496
rect 58341 37438 59879 37440
rect 58341 37435 58407 37438
rect 59813 37435 59879 37438
rect 79041 37498 79107 37501
rect 80421 37498 80487 37501
rect 79041 37496 80487 37498
rect 79041 37440 79046 37496
rect 79102 37440 80426 37496
rect 80482 37440 80487 37496
rect 79041 37438 80487 37440
rect 79041 37435 79107 37438
rect 80421 37435 80487 37438
rect 28993 37362 29059 37365
rect 36813 37362 36879 37365
rect 22142 37302 25146 37362
rect 19701 37226 19767 37229
rect 19977 37226 20043 37229
rect 22142 37226 22202 37302
rect 19701 37224 22202 37226
rect 19701 37168 19706 37224
rect 19762 37168 19982 37224
rect 20038 37168 22202 37224
rect 19701 37166 22202 37168
rect 22277 37226 22343 37229
rect 24853 37226 24919 37229
rect 22277 37224 24919 37226
rect 22277 37168 22282 37224
rect 22338 37168 24858 37224
rect 24914 37168 24919 37224
rect 22277 37166 24919 37168
rect 25086 37226 25146 37302
rect 28993 37360 36879 37362
rect 28993 37304 28998 37360
rect 29054 37304 36818 37360
rect 36874 37304 36879 37360
rect 28993 37302 36879 37304
rect 28993 37299 29059 37302
rect 36813 37299 36879 37302
rect 58249 37362 58315 37365
rect 58617 37362 58683 37365
rect 61377 37362 61443 37365
rect 58249 37360 61443 37362
rect 58249 37304 58254 37360
rect 58310 37304 58622 37360
rect 58678 37304 61382 37360
rect 61438 37304 61443 37360
rect 58249 37302 61443 37304
rect 58249 37299 58315 37302
rect 58617 37299 58683 37302
rect 61377 37299 61443 37302
rect 73153 37362 73219 37365
rect 82813 37362 82879 37365
rect 73153 37360 82879 37362
rect 73153 37304 73158 37360
rect 73214 37304 82818 37360
rect 82874 37304 82879 37360
rect 73153 37302 82879 37304
rect 73153 37299 73219 37302
rect 82813 37299 82879 37302
rect 40309 37226 40375 37229
rect 53005 37226 53071 37229
rect 55673 37226 55739 37229
rect 25086 37224 40375 37226
rect 25086 37168 40314 37224
rect 40370 37168 40375 37224
rect 25086 37166 40375 37168
rect 19701 37163 19767 37166
rect 19977 37163 20043 37166
rect 22277 37163 22343 37166
rect 24853 37163 24919 37166
rect 40309 37163 40375 37166
rect 45510 37166 51090 37226
rect 23289 37090 23355 37093
rect 35709 37090 35775 37093
rect 23289 37088 35775 37090
rect 23289 37032 23294 37088
rect 23350 37032 35714 37088
rect 35770 37032 35775 37088
rect 23289 37030 35775 37032
rect 23289 37027 23355 37030
rect 35709 37027 35775 37030
rect 36629 37090 36695 37093
rect 45510 37090 45570 37166
rect 36629 37088 45570 37090
rect 36629 37032 36634 37088
rect 36690 37032 45570 37088
rect 36629 37030 45570 37032
rect 51030 37090 51090 37166
rect 53005 37224 55739 37226
rect 53005 37168 53010 37224
rect 53066 37168 55678 37224
rect 55734 37168 55739 37224
rect 53005 37166 55739 37168
rect 53005 37163 53071 37166
rect 55673 37163 55739 37166
rect 58341 37226 58407 37229
rect 64781 37226 64847 37229
rect 58341 37224 64847 37226
rect 58341 37168 58346 37224
rect 58402 37168 64786 37224
rect 64842 37168 64847 37224
rect 58341 37166 64847 37168
rect 58341 37163 58407 37166
rect 64781 37163 64847 37166
rect 64965 37226 65031 37229
rect 65793 37226 65859 37229
rect 64965 37224 65859 37226
rect 64965 37168 64970 37224
rect 65026 37168 65798 37224
rect 65854 37168 65859 37224
rect 64965 37166 65859 37168
rect 64965 37163 65031 37166
rect 65793 37163 65859 37166
rect 68553 37226 68619 37229
rect 132861 37226 132927 37229
rect 68553 37224 132927 37226
rect 68553 37168 68558 37224
rect 68614 37168 132866 37224
rect 132922 37168 132927 37224
rect 68553 37166 132927 37168
rect 68553 37163 68619 37166
rect 132861 37163 132927 37166
rect 96797 37090 96863 37093
rect 51030 37030 75194 37090
rect 36629 37027 36695 37030
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 24485 36954 24551 36957
rect 74901 36954 74967 36957
rect 24485 36952 50170 36954
rect 24485 36896 24490 36952
rect 24546 36896 50170 36952
rect 24485 36894 50170 36896
rect 24485 36891 24551 36894
rect 16573 36818 16639 36821
rect 30557 36818 30623 36821
rect 16573 36816 30623 36818
rect 16573 36760 16578 36816
rect 16634 36760 30562 36816
rect 30618 36760 30623 36816
rect 16573 36758 30623 36760
rect 16573 36755 16639 36758
rect 30557 36755 30623 36758
rect 36445 36818 36511 36821
rect 37089 36818 37155 36821
rect 36445 36816 37155 36818
rect 36445 36760 36450 36816
rect 36506 36760 37094 36816
rect 37150 36760 37155 36816
rect 36445 36758 37155 36760
rect 36445 36755 36511 36758
rect 37089 36755 37155 36758
rect 43069 36818 43135 36821
rect 50110 36818 50170 36894
rect 50846 36952 74967 36954
rect 50846 36896 74906 36952
rect 74962 36896 74967 36952
rect 50846 36894 74967 36896
rect 50846 36818 50906 36894
rect 74901 36891 74967 36894
rect 74993 36818 75059 36821
rect 43069 36816 45570 36818
rect 43069 36760 43074 36816
rect 43130 36760 45570 36816
rect 43069 36758 45570 36760
rect 50110 36758 50906 36818
rect 51030 36816 75059 36818
rect 51030 36760 74998 36816
rect 75054 36760 75059 36816
rect 51030 36758 75059 36760
rect 75134 36818 75194 37030
rect 81390 37088 96863 37090
rect 81390 37032 96802 37088
rect 96858 37032 96863 37088
rect 81390 37030 96863 37032
rect 81010 37024 81326 37025
rect 81010 36960 81016 37024
rect 81080 36960 81096 37024
rect 81160 36960 81176 37024
rect 81240 36960 81256 37024
rect 81320 36960 81326 37024
rect 81010 36959 81326 36960
rect 75453 36954 75519 36957
rect 76649 36954 76715 36957
rect 75453 36952 76715 36954
rect 75453 36896 75458 36952
rect 75514 36896 76654 36952
rect 76710 36896 76715 36952
rect 75453 36894 76715 36896
rect 75453 36891 75519 36894
rect 76649 36891 76715 36894
rect 79961 36954 80027 36957
rect 80329 36954 80395 36957
rect 79961 36952 80395 36954
rect 79961 36896 79966 36952
rect 80022 36896 80334 36952
rect 80390 36896 80395 36952
rect 79961 36894 80395 36896
rect 79961 36891 80027 36894
rect 80329 36891 80395 36894
rect 81390 36818 81450 37030
rect 96797 37027 96863 37030
rect 111730 37024 112046 37025
rect 111730 36960 111736 37024
rect 111800 36960 111816 37024
rect 111880 36960 111896 37024
rect 111960 36960 111976 37024
rect 112040 36960 112046 37024
rect 111730 36959 112046 36960
rect 142450 37024 142766 37025
rect 142450 36960 142456 37024
rect 142520 36960 142536 37024
rect 142600 36960 142616 37024
rect 142680 36960 142696 37024
rect 142760 36960 142766 37024
rect 142450 36959 142766 36960
rect 75134 36758 81450 36818
rect 84745 36818 84811 36821
rect 107101 36818 107167 36821
rect 84745 36816 107167 36818
rect 84745 36760 84750 36816
rect 84806 36760 107106 36816
rect 107162 36760 107167 36816
rect 84745 36758 107167 36760
rect 43069 36755 43135 36758
rect 12893 36682 12959 36685
rect 22737 36682 22803 36685
rect 23381 36682 23447 36685
rect 12893 36680 23447 36682
rect 12893 36624 12898 36680
rect 12954 36624 22742 36680
rect 22798 36624 23386 36680
rect 23442 36624 23447 36680
rect 12893 36622 23447 36624
rect 12893 36619 12959 36622
rect 22737 36619 22803 36622
rect 23381 36619 23447 36622
rect 41045 36682 41111 36685
rect 44173 36682 44239 36685
rect 41045 36680 44239 36682
rect 41045 36624 41050 36680
rect 41106 36624 44178 36680
rect 44234 36624 44239 36680
rect 41045 36622 44239 36624
rect 45510 36682 45570 36758
rect 51030 36682 51090 36758
rect 74993 36755 75059 36758
rect 84745 36755 84811 36758
rect 107101 36755 107167 36758
rect 109401 36818 109467 36821
rect 128353 36818 128419 36821
rect 109401 36816 128419 36818
rect 109401 36760 109406 36816
rect 109462 36760 128358 36816
rect 128414 36760 128419 36816
rect 109401 36758 128419 36760
rect 109401 36755 109467 36758
rect 128353 36755 128419 36758
rect 45510 36622 51090 36682
rect 51257 36682 51323 36685
rect 57145 36682 57211 36685
rect 100201 36682 100267 36685
rect 51257 36680 57211 36682
rect 51257 36624 51262 36680
rect 51318 36624 57150 36680
rect 57206 36624 57211 36680
rect 51257 36622 57211 36624
rect 41045 36619 41111 36622
rect 44173 36619 44239 36622
rect 51257 36619 51323 36622
rect 57145 36619 57211 36622
rect 60690 36680 100267 36682
rect 60690 36624 100206 36680
rect 100262 36624 100267 36680
rect 60690 36622 100267 36624
rect 20253 36546 20319 36549
rect 20805 36546 20871 36549
rect 20253 36544 20871 36546
rect 20253 36488 20258 36544
rect 20314 36488 20810 36544
rect 20866 36488 20871 36544
rect 20253 36486 20871 36488
rect 20253 36483 20319 36486
rect 20805 36483 20871 36486
rect 38561 36546 38627 36549
rect 60690 36546 60750 36622
rect 100201 36619 100267 36622
rect 111885 36682 111951 36685
rect 129549 36682 129615 36685
rect 111885 36680 129615 36682
rect 111885 36624 111890 36680
rect 111946 36624 129554 36680
rect 129610 36624 129615 36680
rect 111885 36622 129615 36624
rect 111885 36619 111951 36622
rect 129549 36619 129615 36622
rect 38561 36544 60750 36546
rect 38561 36488 38566 36544
rect 38622 36488 60750 36544
rect 38561 36486 60750 36488
rect 74993 36546 75059 36549
rect 84745 36546 84811 36549
rect 74993 36544 84811 36546
rect 74993 36488 74998 36544
rect 75054 36488 84750 36544
rect 84806 36488 84811 36544
rect 74993 36486 84811 36488
rect 38561 36483 38627 36486
rect 74993 36483 75059 36486
rect 84745 36483 84811 36486
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 65650 36480 65966 36481
rect 65650 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65966 36480
rect 65650 36415 65966 36416
rect 96370 36480 96686 36481
rect 96370 36416 96376 36480
rect 96440 36416 96456 36480
rect 96520 36416 96536 36480
rect 96600 36416 96616 36480
rect 96680 36416 96686 36480
rect 96370 36415 96686 36416
rect 127090 36480 127406 36481
rect 127090 36416 127096 36480
rect 127160 36416 127176 36480
rect 127240 36416 127256 36480
rect 127320 36416 127336 36480
rect 127400 36416 127406 36480
rect 127090 36415 127406 36416
rect 39941 36410 40007 36413
rect 43713 36410 43779 36413
rect 39941 36408 43779 36410
rect 39941 36352 39946 36408
rect 40002 36352 43718 36408
rect 43774 36352 43779 36408
rect 39941 36350 43779 36352
rect 39941 36347 40007 36350
rect 43713 36347 43779 36350
rect 44173 36410 44239 36413
rect 53005 36410 53071 36413
rect 44173 36408 53071 36410
rect 44173 36352 44178 36408
rect 44234 36352 53010 36408
rect 53066 36352 53071 36408
rect 44173 36350 53071 36352
rect 44173 36347 44239 36350
rect 53005 36347 53071 36350
rect 74901 36410 74967 36413
rect 84653 36410 84719 36413
rect 74901 36408 84719 36410
rect 74901 36352 74906 36408
rect 74962 36352 84658 36408
rect 84714 36352 84719 36408
rect 74901 36350 84719 36352
rect 74901 36347 74967 36350
rect 84653 36347 84719 36350
rect 110229 36410 110295 36413
rect 115841 36410 115907 36413
rect 110229 36408 115907 36410
rect 110229 36352 110234 36408
rect 110290 36352 115846 36408
rect 115902 36352 115907 36408
rect 110229 36350 115907 36352
rect 110229 36347 110295 36350
rect 115841 36347 115907 36350
rect 21265 36274 21331 36277
rect 34421 36274 34487 36277
rect 42885 36274 42951 36277
rect 21265 36272 31034 36274
rect 21265 36216 21270 36272
rect 21326 36216 31034 36272
rect 21265 36214 31034 36216
rect 21265 36211 21331 36214
rect 15101 36138 15167 36141
rect 30974 36138 31034 36214
rect 34421 36272 42951 36274
rect 34421 36216 34426 36272
rect 34482 36216 42890 36272
rect 42946 36216 42951 36272
rect 34421 36214 42951 36216
rect 34421 36211 34487 36214
rect 42885 36211 42951 36214
rect 43805 36274 43871 36277
rect 105353 36274 105419 36277
rect 43805 36272 105419 36274
rect 43805 36216 43810 36272
rect 43866 36216 105358 36272
rect 105414 36216 105419 36272
rect 43805 36214 105419 36216
rect 43805 36211 43871 36214
rect 105353 36211 105419 36214
rect 124213 36274 124279 36277
rect 131665 36274 131731 36277
rect 124213 36272 131731 36274
rect 124213 36216 124218 36272
rect 124274 36216 131670 36272
rect 131726 36216 131731 36272
rect 124213 36214 131731 36216
rect 124213 36211 124279 36214
rect 131665 36211 131731 36214
rect 41045 36138 41111 36141
rect 15101 36136 26250 36138
rect 15101 36080 15106 36136
rect 15162 36080 26250 36136
rect 15101 36078 26250 36080
rect 30974 36136 41111 36138
rect 30974 36080 41050 36136
rect 41106 36080 41111 36136
rect 30974 36078 41111 36080
rect 15101 36075 15167 36078
rect 26190 36002 26250 36078
rect 41045 36075 41111 36078
rect 41229 36138 41295 36141
rect 41689 36138 41755 36141
rect 102685 36138 102751 36141
rect 41229 36136 102751 36138
rect 41229 36080 41234 36136
rect 41290 36080 41694 36136
rect 41750 36080 102690 36136
rect 102746 36080 102751 36136
rect 41229 36078 102751 36080
rect 41229 36075 41295 36078
rect 41689 36075 41755 36078
rect 102685 36075 102751 36078
rect 45277 36002 45343 36005
rect 26190 36000 45343 36002
rect 26190 35944 45282 36000
rect 45338 35944 45343 36000
rect 26190 35942 45343 35944
rect 45277 35939 45343 35942
rect 50705 36002 50771 36005
rect 56133 36002 56199 36005
rect 50705 36000 56199 36002
rect 50705 35944 50710 36000
rect 50766 35944 56138 36000
rect 56194 35944 56199 36000
rect 50705 35942 56199 35944
rect 50705 35939 50771 35942
rect 56133 35939 56199 35942
rect 61745 36002 61811 36005
rect 66437 36002 66503 36005
rect 61745 36000 66503 36002
rect 61745 35944 61750 36000
rect 61806 35944 66442 36000
rect 66498 35944 66503 36000
rect 61745 35942 66503 35944
rect 61745 35939 61811 35942
rect 66437 35939 66503 35942
rect 68185 36002 68251 36005
rect 76557 36002 76623 36005
rect 68185 36000 76623 36002
rect 68185 35944 68190 36000
rect 68246 35944 76562 36000
rect 76618 35944 76623 36000
rect 68185 35942 76623 35944
rect 68185 35939 68251 35942
rect 76557 35939 76623 35942
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 81010 35936 81326 35937
rect 81010 35872 81016 35936
rect 81080 35872 81096 35936
rect 81160 35872 81176 35936
rect 81240 35872 81256 35936
rect 81320 35872 81326 35936
rect 81010 35871 81326 35872
rect 111730 35936 112046 35937
rect 111730 35872 111736 35936
rect 111800 35872 111816 35936
rect 111880 35872 111896 35936
rect 111960 35872 111976 35936
rect 112040 35872 112046 35936
rect 111730 35871 112046 35872
rect 142450 35936 142766 35937
rect 142450 35872 142456 35936
rect 142520 35872 142536 35936
rect 142600 35872 142616 35936
rect 142680 35872 142696 35936
rect 142760 35872 142766 35936
rect 142450 35871 142766 35872
rect 53741 35866 53807 35869
rect 77293 35866 77359 35869
rect 53741 35864 77359 35866
rect 53741 35808 53746 35864
rect 53802 35808 77298 35864
rect 77354 35808 77359 35864
rect 53741 35806 77359 35808
rect 53741 35803 53807 35806
rect 77293 35803 77359 35806
rect 30005 35730 30071 35733
rect 80421 35730 80487 35733
rect 30005 35728 80487 35730
rect 30005 35672 30010 35728
rect 30066 35672 80426 35728
rect 80482 35672 80487 35728
rect 30005 35670 80487 35672
rect 30005 35667 30071 35670
rect 80421 35667 80487 35670
rect 41137 35594 41203 35597
rect 41413 35594 41479 35597
rect 41137 35592 41479 35594
rect 41137 35536 41142 35592
rect 41198 35536 41418 35592
rect 41474 35536 41479 35592
rect 41137 35534 41479 35536
rect 41137 35531 41203 35534
rect 41413 35531 41479 35534
rect 50889 35594 50955 35597
rect 98361 35594 98427 35597
rect 50889 35592 98427 35594
rect 50889 35536 50894 35592
rect 50950 35536 98366 35592
rect 98422 35536 98427 35592
rect 50889 35534 98427 35536
rect 50889 35531 50955 35534
rect 98361 35531 98427 35534
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 65650 35392 65966 35393
rect 65650 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65966 35392
rect 65650 35327 65966 35328
rect 96370 35392 96686 35393
rect 96370 35328 96376 35392
rect 96440 35328 96456 35392
rect 96520 35328 96536 35392
rect 96600 35328 96616 35392
rect 96680 35328 96686 35392
rect 96370 35327 96686 35328
rect 127090 35392 127406 35393
rect 127090 35328 127096 35392
rect 127160 35328 127176 35392
rect 127240 35328 127256 35392
rect 127320 35328 127336 35392
rect 127400 35328 127406 35392
rect 127090 35327 127406 35328
rect 34697 35186 34763 35189
rect 51441 35186 51507 35189
rect 34697 35184 51507 35186
rect 34697 35128 34702 35184
rect 34758 35128 51446 35184
rect 51502 35128 51507 35184
rect 34697 35126 51507 35128
rect 34697 35123 34763 35126
rect 51441 35123 51507 35126
rect 71681 35186 71747 35189
rect 134517 35186 134583 35189
rect 71681 35184 134583 35186
rect 71681 35128 71686 35184
rect 71742 35128 134522 35184
rect 134578 35128 134583 35184
rect 71681 35126 134583 35128
rect 71681 35123 71747 35126
rect 134517 35123 134583 35126
rect 43345 35050 43411 35053
rect 44541 35050 44607 35053
rect 43345 35048 44607 35050
rect 43345 34992 43350 35048
rect 43406 34992 44546 35048
rect 44602 34992 44607 35048
rect 43345 34990 44607 34992
rect 43345 34987 43411 34990
rect 44541 34987 44607 34990
rect 65241 35050 65307 35053
rect 129273 35050 129339 35053
rect 65241 35048 129339 35050
rect 65241 34992 65246 35048
rect 65302 34992 129278 35048
rect 129334 34992 129339 35048
rect 65241 34990 129339 34992
rect 65241 34987 65307 34990
rect 129273 34987 129339 34990
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 81010 34848 81326 34849
rect 81010 34784 81016 34848
rect 81080 34784 81096 34848
rect 81160 34784 81176 34848
rect 81240 34784 81256 34848
rect 81320 34784 81326 34848
rect 81010 34783 81326 34784
rect 111730 34848 112046 34849
rect 111730 34784 111736 34848
rect 111800 34784 111816 34848
rect 111880 34784 111896 34848
rect 111960 34784 111976 34848
rect 112040 34784 112046 34848
rect 111730 34783 112046 34784
rect 142450 34848 142766 34849
rect 142450 34784 142456 34848
rect 142520 34784 142536 34848
rect 142600 34784 142616 34848
rect 142680 34784 142696 34848
rect 142760 34784 142766 34848
rect 142450 34783 142766 34784
rect 37181 34506 37247 34509
rect 92841 34506 92907 34509
rect 37181 34504 92907 34506
rect 37181 34448 37186 34504
rect 37242 34448 92846 34504
rect 92902 34448 92907 34504
rect 37181 34446 92907 34448
rect 37181 34443 37247 34446
rect 92841 34443 92907 34446
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 65650 34304 65966 34305
rect 65650 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65966 34304
rect 65650 34239 65966 34240
rect 96370 34304 96686 34305
rect 96370 34240 96376 34304
rect 96440 34240 96456 34304
rect 96520 34240 96536 34304
rect 96600 34240 96616 34304
rect 96680 34240 96686 34304
rect 96370 34239 96686 34240
rect 127090 34304 127406 34305
rect 127090 34240 127096 34304
rect 127160 34240 127176 34304
rect 127240 34240 127256 34304
rect 127320 34240 127336 34304
rect 127400 34240 127406 34304
rect 127090 34239 127406 34240
rect 41965 34098 42031 34101
rect 92105 34098 92171 34101
rect 41965 34096 92171 34098
rect 41965 34040 41970 34096
rect 42026 34040 92110 34096
rect 92166 34040 92171 34096
rect 41965 34038 92171 34040
rect 41965 34035 42031 34038
rect 92105 34035 92171 34038
rect 31753 33962 31819 33965
rect 89069 33962 89135 33965
rect 31753 33960 89135 33962
rect 31753 33904 31758 33960
rect 31814 33904 89074 33960
rect 89130 33904 89135 33960
rect 31753 33902 89135 33904
rect 31753 33899 31819 33902
rect 89069 33899 89135 33902
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 81010 33760 81326 33761
rect 81010 33696 81016 33760
rect 81080 33696 81096 33760
rect 81160 33696 81176 33760
rect 81240 33696 81256 33760
rect 81320 33696 81326 33760
rect 81010 33695 81326 33696
rect 111730 33760 112046 33761
rect 111730 33696 111736 33760
rect 111800 33696 111816 33760
rect 111880 33696 111896 33760
rect 111960 33696 111976 33760
rect 112040 33696 112046 33760
rect 111730 33695 112046 33696
rect 142450 33760 142766 33761
rect 142450 33696 142456 33760
rect 142520 33696 142536 33760
rect 142600 33696 142616 33760
rect 142680 33696 142696 33760
rect 142760 33696 142766 33760
rect 142450 33695 142766 33696
rect 41321 33554 41387 33557
rect 95877 33554 95943 33557
rect 41321 33552 95943 33554
rect 41321 33496 41326 33552
rect 41382 33496 95882 33552
rect 95938 33496 95943 33552
rect 41321 33494 95943 33496
rect 41321 33491 41387 33494
rect 95877 33491 95943 33494
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 65650 33216 65966 33217
rect 65650 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65966 33216
rect 65650 33151 65966 33152
rect 96370 33216 96686 33217
rect 96370 33152 96376 33216
rect 96440 33152 96456 33216
rect 96520 33152 96536 33216
rect 96600 33152 96616 33216
rect 96680 33152 96686 33216
rect 96370 33151 96686 33152
rect 127090 33216 127406 33217
rect 127090 33152 127096 33216
rect 127160 33152 127176 33216
rect 127240 33152 127256 33216
rect 127320 33152 127336 33216
rect 127400 33152 127406 33216
rect 127090 33151 127406 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 81010 32672 81326 32673
rect 81010 32608 81016 32672
rect 81080 32608 81096 32672
rect 81160 32608 81176 32672
rect 81240 32608 81256 32672
rect 81320 32608 81326 32672
rect 81010 32607 81326 32608
rect 111730 32672 112046 32673
rect 111730 32608 111736 32672
rect 111800 32608 111816 32672
rect 111880 32608 111896 32672
rect 111960 32608 111976 32672
rect 112040 32608 112046 32672
rect 111730 32607 112046 32608
rect 142450 32672 142766 32673
rect 142450 32608 142456 32672
rect 142520 32608 142536 32672
rect 142600 32608 142616 32672
rect 142680 32608 142696 32672
rect 142760 32608 142766 32672
rect 142450 32607 142766 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 65650 32128 65966 32129
rect 65650 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65966 32128
rect 65650 32063 65966 32064
rect 96370 32128 96686 32129
rect 96370 32064 96376 32128
rect 96440 32064 96456 32128
rect 96520 32064 96536 32128
rect 96600 32064 96616 32128
rect 96680 32064 96686 32128
rect 96370 32063 96686 32064
rect 127090 32128 127406 32129
rect 127090 32064 127096 32128
rect 127160 32064 127176 32128
rect 127240 32064 127256 32128
rect 127320 32064 127336 32128
rect 127400 32064 127406 32128
rect 127090 32063 127406 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 81010 31584 81326 31585
rect 81010 31520 81016 31584
rect 81080 31520 81096 31584
rect 81160 31520 81176 31584
rect 81240 31520 81256 31584
rect 81320 31520 81326 31584
rect 81010 31519 81326 31520
rect 111730 31584 112046 31585
rect 111730 31520 111736 31584
rect 111800 31520 111816 31584
rect 111880 31520 111896 31584
rect 111960 31520 111976 31584
rect 112040 31520 112046 31584
rect 111730 31519 112046 31520
rect 142450 31584 142766 31585
rect 142450 31520 142456 31584
rect 142520 31520 142536 31584
rect 142600 31520 142616 31584
rect 142680 31520 142696 31584
rect 142760 31520 142766 31584
rect 142450 31519 142766 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 65650 31040 65966 31041
rect 65650 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65966 31040
rect 65650 30975 65966 30976
rect 96370 31040 96686 31041
rect 96370 30976 96376 31040
rect 96440 30976 96456 31040
rect 96520 30976 96536 31040
rect 96600 30976 96616 31040
rect 96680 30976 96686 31040
rect 96370 30975 96686 30976
rect 127090 31040 127406 31041
rect 127090 30976 127096 31040
rect 127160 30976 127176 31040
rect 127240 30976 127256 31040
rect 127320 30976 127336 31040
rect 127400 30976 127406 31040
rect 127090 30975 127406 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 81010 30496 81326 30497
rect 81010 30432 81016 30496
rect 81080 30432 81096 30496
rect 81160 30432 81176 30496
rect 81240 30432 81256 30496
rect 81320 30432 81326 30496
rect 81010 30431 81326 30432
rect 111730 30496 112046 30497
rect 111730 30432 111736 30496
rect 111800 30432 111816 30496
rect 111880 30432 111896 30496
rect 111960 30432 111976 30496
rect 112040 30432 112046 30496
rect 111730 30431 112046 30432
rect 142450 30496 142766 30497
rect 142450 30432 142456 30496
rect 142520 30432 142536 30496
rect 142600 30432 142616 30496
rect 142680 30432 142696 30496
rect 142760 30432 142766 30496
rect 142450 30431 142766 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 65650 29952 65966 29953
rect 65650 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65966 29952
rect 65650 29887 65966 29888
rect 96370 29952 96686 29953
rect 96370 29888 96376 29952
rect 96440 29888 96456 29952
rect 96520 29888 96536 29952
rect 96600 29888 96616 29952
rect 96680 29888 96686 29952
rect 96370 29887 96686 29888
rect 127090 29952 127406 29953
rect 127090 29888 127096 29952
rect 127160 29888 127176 29952
rect 127240 29888 127256 29952
rect 127320 29888 127336 29952
rect 127400 29888 127406 29952
rect 127090 29887 127406 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 81010 29408 81326 29409
rect 81010 29344 81016 29408
rect 81080 29344 81096 29408
rect 81160 29344 81176 29408
rect 81240 29344 81256 29408
rect 81320 29344 81326 29408
rect 81010 29343 81326 29344
rect 111730 29408 112046 29409
rect 111730 29344 111736 29408
rect 111800 29344 111816 29408
rect 111880 29344 111896 29408
rect 111960 29344 111976 29408
rect 112040 29344 112046 29408
rect 111730 29343 112046 29344
rect 142450 29408 142766 29409
rect 142450 29344 142456 29408
rect 142520 29344 142536 29408
rect 142600 29344 142616 29408
rect 142680 29344 142696 29408
rect 142760 29344 142766 29408
rect 142450 29343 142766 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 65650 28864 65966 28865
rect 65650 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65966 28864
rect 65650 28799 65966 28800
rect 96370 28864 96686 28865
rect 96370 28800 96376 28864
rect 96440 28800 96456 28864
rect 96520 28800 96536 28864
rect 96600 28800 96616 28864
rect 96680 28800 96686 28864
rect 96370 28799 96686 28800
rect 127090 28864 127406 28865
rect 127090 28800 127096 28864
rect 127160 28800 127176 28864
rect 127240 28800 127256 28864
rect 127320 28800 127336 28864
rect 127400 28800 127406 28864
rect 127090 28799 127406 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 81010 28320 81326 28321
rect 81010 28256 81016 28320
rect 81080 28256 81096 28320
rect 81160 28256 81176 28320
rect 81240 28256 81256 28320
rect 81320 28256 81326 28320
rect 81010 28255 81326 28256
rect 111730 28320 112046 28321
rect 111730 28256 111736 28320
rect 111800 28256 111816 28320
rect 111880 28256 111896 28320
rect 111960 28256 111976 28320
rect 112040 28256 112046 28320
rect 111730 28255 112046 28256
rect 142450 28320 142766 28321
rect 142450 28256 142456 28320
rect 142520 28256 142536 28320
rect 142600 28256 142616 28320
rect 142680 28256 142696 28320
rect 142760 28256 142766 28320
rect 142450 28255 142766 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 65650 27776 65966 27777
rect 65650 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65966 27776
rect 65650 27711 65966 27712
rect 96370 27776 96686 27777
rect 96370 27712 96376 27776
rect 96440 27712 96456 27776
rect 96520 27712 96536 27776
rect 96600 27712 96616 27776
rect 96680 27712 96686 27776
rect 96370 27711 96686 27712
rect 127090 27776 127406 27777
rect 127090 27712 127096 27776
rect 127160 27712 127176 27776
rect 127240 27712 127256 27776
rect 127320 27712 127336 27776
rect 127400 27712 127406 27776
rect 127090 27711 127406 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 81010 27232 81326 27233
rect 81010 27168 81016 27232
rect 81080 27168 81096 27232
rect 81160 27168 81176 27232
rect 81240 27168 81256 27232
rect 81320 27168 81326 27232
rect 81010 27167 81326 27168
rect 111730 27232 112046 27233
rect 111730 27168 111736 27232
rect 111800 27168 111816 27232
rect 111880 27168 111896 27232
rect 111960 27168 111976 27232
rect 112040 27168 112046 27232
rect 111730 27167 112046 27168
rect 142450 27232 142766 27233
rect 142450 27168 142456 27232
rect 142520 27168 142536 27232
rect 142600 27168 142616 27232
rect 142680 27168 142696 27232
rect 142760 27168 142766 27232
rect 142450 27167 142766 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 65650 26688 65966 26689
rect 65650 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65966 26688
rect 65650 26623 65966 26624
rect 96370 26688 96686 26689
rect 96370 26624 96376 26688
rect 96440 26624 96456 26688
rect 96520 26624 96536 26688
rect 96600 26624 96616 26688
rect 96680 26624 96686 26688
rect 96370 26623 96686 26624
rect 127090 26688 127406 26689
rect 127090 26624 127096 26688
rect 127160 26624 127176 26688
rect 127240 26624 127256 26688
rect 127320 26624 127336 26688
rect 127400 26624 127406 26688
rect 127090 26623 127406 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 81010 26144 81326 26145
rect 81010 26080 81016 26144
rect 81080 26080 81096 26144
rect 81160 26080 81176 26144
rect 81240 26080 81256 26144
rect 81320 26080 81326 26144
rect 81010 26079 81326 26080
rect 111730 26144 112046 26145
rect 111730 26080 111736 26144
rect 111800 26080 111816 26144
rect 111880 26080 111896 26144
rect 111960 26080 111976 26144
rect 112040 26080 112046 26144
rect 111730 26079 112046 26080
rect 142450 26144 142766 26145
rect 142450 26080 142456 26144
rect 142520 26080 142536 26144
rect 142600 26080 142616 26144
rect 142680 26080 142696 26144
rect 142760 26080 142766 26144
rect 142450 26079 142766 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 65650 25600 65966 25601
rect 65650 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65966 25600
rect 65650 25535 65966 25536
rect 96370 25600 96686 25601
rect 96370 25536 96376 25600
rect 96440 25536 96456 25600
rect 96520 25536 96536 25600
rect 96600 25536 96616 25600
rect 96680 25536 96686 25600
rect 96370 25535 96686 25536
rect 127090 25600 127406 25601
rect 127090 25536 127096 25600
rect 127160 25536 127176 25600
rect 127240 25536 127256 25600
rect 127320 25536 127336 25600
rect 127400 25536 127406 25600
rect 127090 25535 127406 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 81010 25056 81326 25057
rect 81010 24992 81016 25056
rect 81080 24992 81096 25056
rect 81160 24992 81176 25056
rect 81240 24992 81256 25056
rect 81320 24992 81326 25056
rect 81010 24991 81326 24992
rect 111730 25056 112046 25057
rect 111730 24992 111736 25056
rect 111800 24992 111816 25056
rect 111880 24992 111896 25056
rect 111960 24992 111976 25056
rect 112040 24992 112046 25056
rect 111730 24991 112046 24992
rect 142450 25056 142766 25057
rect 142450 24992 142456 25056
rect 142520 24992 142536 25056
rect 142600 24992 142616 25056
rect 142680 24992 142696 25056
rect 142760 24992 142766 25056
rect 142450 24991 142766 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 65650 24512 65966 24513
rect 65650 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65966 24512
rect 65650 24447 65966 24448
rect 96370 24512 96686 24513
rect 96370 24448 96376 24512
rect 96440 24448 96456 24512
rect 96520 24448 96536 24512
rect 96600 24448 96616 24512
rect 96680 24448 96686 24512
rect 96370 24447 96686 24448
rect 127090 24512 127406 24513
rect 127090 24448 127096 24512
rect 127160 24448 127176 24512
rect 127240 24448 127256 24512
rect 127320 24448 127336 24512
rect 127400 24448 127406 24512
rect 127090 24447 127406 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 81010 23968 81326 23969
rect 81010 23904 81016 23968
rect 81080 23904 81096 23968
rect 81160 23904 81176 23968
rect 81240 23904 81256 23968
rect 81320 23904 81326 23968
rect 81010 23903 81326 23904
rect 111730 23968 112046 23969
rect 111730 23904 111736 23968
rect 111800 23904 111816 23968
rect 111880 23904 111896 23968
rect 111960 23904 111976 23968
rect 112040 23904 112046 23968
rect 111730 23903 112046 23904
rect 142450 23968 142766 23969
rect 142450 23904 142456 23968
rect 142520 23904 142536 23968
rect 142600 23904 142616 23968
rect 142680 23904 142696 23968
rect 142760 23904 142766 23968
rect 142450 23903 142766 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 65650 23424 65966 23425
rect 65650 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65966 23424
rect 65650 23359 65966 23360
rect 96370 23424 96686 23425
rect 96370 23360 96376 23424
rect 96440 23360 96456 23424
rect 96520 23360 96536 23424
rect 96600 23360 96616 23424
rect 96680 23360 96686 23424
rect 96370 23359 96686 23360
rect 127090 23424 127406 23425
rect 127090 23360 127096 23424
rect 127160 23360 127176 23424
rect 127240 23360 127256 23424
rect 127320 23360 127336 23424
rect 127400 23360 127406 23424
rect 127090 23359 127406 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 81010 22880 81326 22881
rect 81010 22816 81016 22880
rect 81080 22816 81096 22880
rect 81160 22816 81176 22880
rect 81240 22816 81256 22880
rect 81320 22816 81326 22880
rect 81010 22815 81326 22816
rect 111730 22880 112046 22881
rect 111730 22816 111736 22880
rect 111800 22816 111816 22880
rect 111880 22816 111896 22880
rect 111960 22816 111976 22880
rect 112040 22816 112046 22880
rect 111730 22815 112046 22816
rect 142450 22880 142766 22881
rect 142450 22816 142456 22880
rect 142520 22816 142536 22880
rect 142600 22816 142616 22880
rect 142680 22816 142696 22880
rect 142760 22816 142766 22880
rect 142450 22815 142766 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 65650 22336 65966 22337
rect 65650 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65966 22336
rect 65650 22271 65966 22272
rect 96370 22336 96686 22337
rect 96370 22272 96376 22336
rect 96440 22272 96456 22336
rect 96520 22272 96536 22336
rect 96600 22272 96616 22336
rect 96680 22272 96686 22336
rect 96370 22271 96686 22272
rect 127090 22336 127406 22337
rect 127090 22272 127096 22336
rect 127160 22272 127176 22336
rect 127240 22272 127256 22336
rect 127320 22272 127336 22336
rect 127400 22272 127406 22336
rect 127090 22271 127406 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 81010 21792 81326 21793
rect 81010 21728 81016 21792
rect 81080 21728 81096 21792
rect 81160 21728 81176 21792
rect 81240 21728 81256 21792
rect 81320 21728 81326 21792
rect 81010 21727 81326 21728
rect 111730 21792 112046 21793
rect 111730 21728 111736 21792
rect 111800 21728 111816 21792
rect 111880 21728 111896 21792
rect 111960 21728 111976 21792
rect 112040 21728 112046 21792
rect 111730 21727 112046 21728
rect 142450 21792 142766 21793
rect 142450 21728 142456 21792
rect 142520 21728 142536 21792
rect 142600 21728 142616 21792
rect 142680 21728 142696 21792
rect 142760 21728 142766 21792
rect 142450 21727 142766 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 65650 21248 65966 21249
rect 65650 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65966 21248
rect 65650 21183 65966 21184
rect 96370 21248 96686 21249
rect 96370 21184 96376 21248
rect 96440 21184 96456 21248
rect 96520 21184 96536 21248
rect 96600 21184 96616 21248
rect 96680 21184 96686 21248
rect 96370 21183 96686 21184
rect 127090 21248 127406 21249
rect 127090 21184 127096 21248
rect 127160 21184 127176 21248
rect 127240 21184 127256 21248
rect 127320 21184 127336 21248
rect 127400 21184 127406 21248
rect 127090 21183 127406 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 81010 20704 81326 20705
rect 81010 20640 81016 20704
rect 81080 20640 81096 20704
rect 81160 20640 81176 20704
rect 81240 20640 81256 20704
rect 81320 20640 81326 20704
rect 81010 20639 81326 20640
rect 111730 20704 112046 20705
rect 111730 20640 111736 20704
rect 111800 20640 111816 20704
rect 111880 20640 111896 20704
rect 111960 20640 111976 20704
rect 112040 20640 112046 20704
rect 111730 20639 112046 20640
rect 142450 20704 142766 20705
rect 142450 20640 142456 20704
rect 142520 20640 142536 20704
rect 142600 20640 142616 20704
rect 142680 20640 142696 20704
rect 142760 20640 142766 20704
rect 142450 20639 142766 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 65650 20160 65966 20161
rect 65650 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65966 20160
rect 65650 20095 65966 20096
rect 96370 20160 96686 20161
rect 96370 20096 96376 20160
rect 96440 20096 96456 20160
rect 96520 20096 96536 20160
rect 96600 20096 96616 20160
rect 96680 20096 96686 20160
rect 96370 20095 96686 20096
rect 127090 20160 127406 20161
rect 127090 20096 127096 20160
rect 127160 20096 127176 20160
rect 127240 20096 127256 20160
rect 127320 20096 127336 20160
rect 127400 20096 127406 20160
rect 127090 20095 127406 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 81010 19616 81326 19617
rect 81010 19552 81016 19616
rect 81080 19552 81096 19616
rect 81160 19552 81176 19616
rect 81240 19552 81256 19616
rect 81320 19552 81326 19616
rect 81010 19551 81326 19552
rect 111730 19616 112046 19617
rect 111730 19552 111736 19616
rect 111800 19552 111816 19616
rect 111880 19552 111896 19616
rect 111960 19552 111976 19616
rect 112040 19552 112046 19616
rect 111730 19551 112046 19552
rect 142450 19616 142766 19617
rect 142450 19552 142456 19616
rect 142520 19552 142536 19616
rect 142600 19552 142616 19616
rect 142680 19552 142696 19616
rect 142760 19552 142766 19616
rect 142450 19551 142766 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 65650 19072 65966 19073
rect 65650 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65966 19072
rect 65650 19007 65966 19008
rect 96370 19072 96686 19073
rect 96370 19008 96376 19072
rect 96440 19008 96456 19072
rect 96520 19008 96536 19072
rect 96600 19008 96616 19072
rect 96680 19008 96686 19072
rect 96370 19007 96686 19008
rect 127090 19072 127406 19073
rect 127090 19008 127096 19072
rect 127160 19008 127176 19072
rect 127240 19008 127256 19072
rect 127320 19008 127336 19072
rect 127400 19008 127406 19072
rect 127090 19007 127406 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 81010 18528 81326 18529
rect 81010 18464 81016 18528
rect 81080 18464 81096 18528
rect 81160 18464 81176 18528
rect 81240 18464 81256 18528
rect 81320 18464 81326 18528
rect 81010 18463 81326 18464
rect 111730 18528 112046 18529
rect 111730 18464 111736 18528
rect 111800 18464 111816 18528
rect 111880 18464 111896 18528
rect 111960 18464 111976 18528
rect 112040 18464 112046 18528
rect 111730 18463 112046 18464
rect 142450 18528 142766 18529
rect 142450 18464 142456 18528
rect 142520 18464 142536 18528
rect 142600 18464 142616 18528
rect 142680 18464 142696 18528
rect 142760 18464 142766 18528
rect 142450 18463 142766 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 65650 17984 65966 17985
rect 65650 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65966 17984
rect 65650 17919 65966 17920
rect 96370 17984 96686 17985
rect 96370 17920 96376 17984
rect 96440 17920 96456 17984
rect 96520 17920 96536 17984
rect 96600 17920 96616 17984
rect 96680 17920 96686 17984
rect 96370 17919 96686 17920
rect 127090 17984 127406 17985
rect 127090 17920 127096 17984
rect 127160 17920 127176 17984
rect 127240 17920 127256 17984
rect 127320 17920 127336 17984
rect 127400 17920 127406 17984
rect 127090 17919 127406 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 81010 17440 81326 17441
rect 81010 17376 81016 17440
rect 81080 17376 81096 17440
rect 81160 17376 81176 17440
rect 81240 17376 81256 17440
rect 81320 17376 81326 17440
rect 81010 17375 81326 17376
rect 111730 17440 112046 17441
rect 111730 17376 111736 17440
rect 111800 17376 111816 17440
rect 111880 17376 111896 17440
rect 111960 17376 111976 17440
rect 112040 17376 112046 17440
rect 111730 17375 112046 17376
rect 142450 17440 142766 17441
rect 142450 17376 142456 17440
rect 142520 17376 142536 17440
rect 142600 17376 142616 17440
rect 142680 17376 142696 17440
rect 142760 17376 142766 17440
rect 142450 17375 142766 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 65650 16896 65966 16897
rect 65650 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65966 16896
rect 65650 16831 65966 16832
rect 96370 16896 96686 16897
rect 96370 16832 96376 16896
rect 96440 16832 96456 16896
rect 96520 16832 96536 16896
rect 96600 16832 96616 16896
rect 96680 16832 96686 16896
rect 96370 16831 96686 16832
rect 127090 16896 127406 16897
rect 127090 16832 127096 16896
rect 127160 16832 127176 16896
rect 127240 16832 127256 16896
rect 127320 16832 127336 16896
rect 127400 16832 127406 16896
rect 127090 16831 127406 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 81010 16352 81326 16353
rect 81010 16288 81016 16352
rect 81080 16288 81096 16352
rect 81160 16288 81176 16352
rect 81240 16288 81256 16352
rect 81320 16288 81326 16352
rect 81010 16287 81326 16288
rect 111730 16352 112046 16353
rect 111730 16288 111736 16352
rect 111800 16288 111816 16352
rect 111880 16288 111896 16352
rect 111960 16288 111976 16352
rect 112040 16288 112046 16352
rect 111730 16287 112046 16288
rect 142450 16352 142766 16353
rect 142450 16288 142456 16352
rect 142520 16288 142536 16352
rect 142600 16288 142616 16352
rect 142680 16288 142696 16352
rect 142760 16288 142766 16352
rect 142450 16287 142766 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 65650 15808 65966 15809
rect 65650 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65966 15808
rect 65650 15743 65966 15744
rect 96370 15808 96686 15809
rect 96370 15744 96376 15808
rect 96440 15744 96456 15808
rect 96520 15744 96536 15808
rect 96600 15744 96616 15808
rect 96680 15744 96686 15808
rect 96370 15743 96686 15744
rect 127090 15808 127406 15809
rect 127090 15744 127096 15808
rect 127160 15744 127176 15808
rect 127240 15744 127256 15808
rect 127320 15744 127336 15808
rect 127400 15744 127406 15808
rect 127090 15743 127406 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 81010 15264 81326 15265
rect 81010 15200 81016 15264
rect 81080 15200 81096 15264
rect 81160 15200 81176 15264
rect 81240 15200 81256 15264
rect 81320 15200 81326 15264
rect 81010 15199 81326 15200
rect 111730 15264 112046 15265
rect 111730 15200 111736 15264
rect 111800 15200 111816 15264
rect 111880 15200 111896 15264
rect 111960 15200 111976 15264
rect 112040 15200 112046 15264
rect 111730 15199 112046 15200
rect 142450 15264 142766 15265
rect 142450 15200 142456 15264
rect 142520 15200 142536 15264
rect 142600 15200 142616 15264
rect 142680 15200 142696 15264
rect 142760 15200 142766 15264
rect 142450 15199 142766 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 65650 14720 65966 14721
rect 65650 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65966 14720
rect 65650 14655 65966 14656
rect 96370 14720 96686 14721
rect 96370 14656 96376 14720
rect 96440 14656 96456 14720
rect 96520 14656 96536 14720
rect 96600 14656 96616 14720
rect 96680 14656 96686 14720
rect 96370 14655 96686 14656
rect 127090 14720 127406 14721
rect 127090 14656 127096 14720
rect 127160 14656 127176 14720
rect 127240 14656 127256 14720
rect 127320 14656 127336 14720
rect 127400 14656 127406 14720
rect 127090 14655 127406 14656
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 81010 14176 81326 14177
rect 81010 14112 81016 14176
rect 81080 14112 81096 14176
rect 81160 14112 81176 14176
rect 81240 14112 81256 14176
rect 81320 14112 81326 14176
rect 81010 14111 81326 14112
rect 111730 14176 112046 14177
rect 111730 14112 111736 14176
rect 111800 14112 111816 14176
rect 111880 14112 111896 14176
rect 111960 14112 111976 14176
rect 112040 14112 112046 14176
rect 111730 14111 112046 14112
rect 142450 14176 142766 14177
rect 142450 14112 142456 14176
rect 142520 14112 142536 14176
rect 142600 14112 142616 14176
rect 142680 14112 142696 14176
rect 142760 14112 142766 14176
rect 142450 14111 142766 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 65650 13632 65966 13633
rect 65650 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65966 13632
rect 65650 13567 65966 13568
rect 96370 13632 96686 13633
rect 96370 13568 96376 13632
rect 96440 13568 96456 13632
rect 96520 13568 96536 13632
rect 96600 13568 96616 13632
rect 96680 13568 96686 13632
rect 96370 13567 96686 13568
rect 127090 13632 127406 13633
rect 127090 13568 127096 13632
rect 127160 13568 127176 13632
rect 127240 13568 127256 13632
rect 127320 13568 127336 13632
rect 127400 13568 127406 13632
rect 127090 13567 127406 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 81010 13088 81326 13089
rect 81010 13024 81016 13088
rect 81080 13024 81096 13088
rect 81160 13024 81176 13088
rect 81240 13024 81256 13088
rect 81320 13024 81326 13088
rect 81010 13023 81326 13024
rect 111730 13088 112046 13089
rect 111730 13024 111736 13088
rect 111800 13024 111816 13088
rect 111880 13024 111896 13088
rect 111960 13024 111976 13088
rect 112040 13024 112046 13088
rect 111730 13023 112046 13024
rect 142450 13088 142766 13089
rect 142450 13024 142456 13088
rect 142520 13024 142536 13088
rect 142600 13024 142616 13088
rect 142680 13024 142696 13088
rect 142760 13024 142766 13088
rect 142450 13023 142766 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 65650 12544 65966 12545
rect 65650 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65966 12544
rect 65650 12479 65966 12480
rect 96370 12544 96686 12545
rect 96370 12480 96376 12544
rect 96440 12480 96456 12544
rect 96520 12480 96536 12544
rect 96600 12480 96616 12544
rect 96680 12480 96686 12544
rect 96370 12479 96686 12480
rect 127090 12544 127406 12545
rect 127090 12480 127096 12544
rect 127160 12480 127176 12544
rect 127240 12480 127256 12544
rect 127320 12480 127336 12544
rect 127400 12480 127406 12544
rect 127090 12479 127406 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 81010 12000 81326 12001
rect 81010 11936 81016 12000
rect 81080 11936 81096 12000
rect 81160 11936 81176 12000
rect 81240 11936 81256 12000
rect 81320 11936 81326 12000
rect 81010 11935 81326 11936
rect 111730 12000 112046 12001
rect 111730 11936 111736 12000
rect 111800 11936 111816 12000
rect 111880 11936 111896 12000
rect 111960 11936 111976 12000
rect 112040 11936 112046 12000
rect 111730 11935 112046 11936
rect 142450 12000 142766 12001
rect 142450 11936 142456 12000
rect 142520 11936 142536 12000
rect 142600 11936 142616 12000
rect 142680 11936 142696 12000
rect 142760 11936 142766 12000
rect 142450 11935 142766 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 65650 11456 65966 11457
rect 65650 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65966 11456
rect 65650 11391 65966 11392
rect 96370 11456 96686 11457
rect 96370 11392 96376 11456
rect 96440 11392 96456 11456
rect 96520 11392 96536 11456
rect 96600 11392 96616 11456
rect 96680 11392 96686 11456
rect 96370 11391 96686 11392
rect 127090 11456 127406 11457
rect 127090 11392 127096 11456
rect 127160 11392 127176 11456
rect 127240 11392 127256 11456
rect 127320 11392 127336 11456
rect 127400 11392 127406 11456
rect 127090 11391 127406 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 81010 10912 81326 10913
rect 81010 10848 81016 10912
rect 81080 10848 81096 10912
rect 81160 10848 81176 10912
rect 81240 10848 81256 10912
rect 81320 10848 81326 10912
rect 81010 10847 81326 10848
rect 111730 10912 112046 10913
rect 111730 10848 111736 10912
rect 111800 10848 111816 10912
rect 111880 10848 111896 10912
rect 111960 10848 111976 10912
rect 112040 10848 112046 10912
rect 111730 10847 112046 10848
rect 142450 10912 142766 10913
rect 142450 10848 142456 10912
rect 142520 10848 142536 10912
rect 142600 10848 142616 10912
rect 142680 10848 142696 10912
rect 142760 10848 142766 10912
rect 142450 10847 142766 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 65650 10368 65966 10369
rect 65650 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65966 10368
rect 65650 10303 65966 10304
rect 96370 10368 96686 10369
rect 96370 10304 96376 10368
rect 96440 10304 96456 10368
rect 96520 10304 96536 10368
rect 96600 10304 96616 10368
rect 96680 10304 96686 10368
rect 96370 10303 96686 10304
rect 127090 10368 127406 10369
rect 127090 10304 127096 10368
rect 127160 10304 127176 10368
rect 127240 10304 127256 10368
rect 127320 10304 127336 10368
rect 127400 10304 127406 10368
rect 127090 10303 127406 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 81010 9824 81326 9825
rect 81010 9760 81016 9824
rect 81080 9760 81096 9824
rect 81160 9760 81176 9824
rect 81240 9760 81256 9824
rect 81320 9760 81326 9824
rect 81010 9759 81326 9760
rect 111730 9824 112046 9825
rect 111730 9760 111736 9824
rect 111800 9760 111816 9824
rect 111880 9760 111896 9824
rect 111960 9760 111976 9824
rect 112040 9760 112046 9824
rect 111730 9759 112046 9760
rect 142450 9824 142766 9825
rect 142450 9760 142456 9824
rect 142520 9760 142536 9824
rect 142600 9760 142616 9824
rect 142680 9760 142696 9824
rect 142760 9760 142766 9824
rect 142450 9759 142766 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 65650 9280 65966 9281
rect 65650 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65966 9280
rect 65650 9215 65966 9216
rect 96370 9280 96686 9281
rect 96370 9216 96376 9280
rect 96440 9216 96456 9280
rect 96520 9216 96536 9280
rect 96600 9216 96616 9280
rect 96680 9216 96686 9280
rect 96370 9215 96686 9216
rect 127090 9280 127406 9281
rect 127090 9216 127096 9280
rect 127160 9216 127176 9280
rect 127240 9216 127256 9280
rect 127320 9216 127336 9280
rect 127400 9216 127406 9280
rect 127090 9215 127406 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 81010 8736 81326 8737
rect 81010 8672 81016 8736
rect 81080 8672 81096 8736
rect 81160 8672 81176 8736
rect 81240 8672 81256 8736
rect 81320 8672 81326 8736
rect 81010 8671 81326 8672
rect 111730 8736 112046 8737
rect 111730 8672 111736 8736
rect 111800 8672 111816 8736
rect 111880 8672 111896 8736
rect 111960 8672 111976 8736
rect 112040 8672 112046 8736
rect 111730 8671 112046 8672
rect 142450 8736 142766 8737
rect 142450 8672 142456 8736
rect 142520 8672 142536 8736
rect 142600 8672 142616 8736
rect 142680 8672 142696 8736
rect 142760 8672 142766 8736
rect 142450 8671 142766 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 65650 8192 65966 8193
rect 65650 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65966 8192
rect 65650 8127 65966 8128
rect 96370 8192 96686 8193
rect 96370 8128 96376 8192
rect 96440 8128 96456 8192
rect 96520 8128 96536 8192
rect 96600 8128 96616 8192
rect 96680 8128 96686 8192
rect 96370 8127 96686 8128
rect 127090 8192 127406 8193
rect 127090 8128 127096 8192
rect 127160 8128 127176 8192
rect 127240 8128 127256 8192
rect 127320 8128 127336 8192
rect 127400 8128 127406 8192
rect 127090 8127 127406 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 81010 7648 81326 7649
rect 81010 7584 81016 7648
rect 81080 7584 81096 7648
rect 81160 7584 81176 7648
rect 81240 7584 81256 7648
rect 81320 7584 81326 7648
rect 81010 7583 81326 7584
rect 111730 7648 112046 7649
rect 111730 7584 111736 7648
rect 111800 7584 111816 7648
rect 111880 7584 111896 7648
rect 111960 7584 111976 7648
rect 112040 7584 112046 7648
rect 111730 7583 112046 7584
rect 142450 7648 142766 7649
rect 142450 7584 142456 7648
rect 142520 7584 142536 7648
rect 142600 7584 142616 7648
rect 142680 7584 142696 7648
rect 142760 7584 142766 7648
rect 142450 7583 142766 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 65650 7104 65966 7105
rect 65650 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65966 7104
rect 65650 7039 65966 7040
rect 96370 7104 96686 7105
rect 96370 7040 96376 7104
rect 96440 7040 96456 7104
rect 96520 7040 96536 7104
rect 96600 7040 96616 7104
rect 96680 7040 96686 7104
rect 96370 7039 96686 7040
rect 127090 7104 127406 7105
rect 127090 7040 127096 7104
rect 127160 7040 127176 7104
rect 127240 7040 127256 7104
rect 127320 7040 127336 7104
rect 127400 7040 127406 7104
rect 127090 7039 127406 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 81010 6560 81326 6561
rect 81010 6496 81016 6560
rect 81080 6496 81096 6560
rect 81160 6496 81176 6560
rect 81240 6496 81256 6560
rect 81320 6496 81326 6560
rect 81010 6495 81326 6496
rect 111730 6560 112046 6561
rect 111730 6496 111736 6560
rect 111800 6496 111816 6560
rect 111880 6496 111896 6560
rect 111960 6496 111976 6560
rect 112040 6496 112046 6560
rect 111730 6495 112046 6496
rect 142450 6560 142766 6561
rect 142450 6496 142456 6560
rect 142520 6496 142536 6560
rect 142600 6496 142616 6560
rect 142680 6496 142696 6560
rect 142760 6496 142766 6560
rect 142450 6495 142766 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 65650 6016 65966 6017
rect 65650 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65966 6016
rect 65650 5951 65966 5952
rect 96370 6016 96686 6017
rect 96370 5952 96376 6016
rect 96440 5952 96456 6016
rect 96520 5952 96536 6016
rect 96600 5952 96616 6016
rect 96680 5952 96686 6016
rect 96370 5951 96686 5952
rect 127090 6016 127406 6017
rect 127090 5952 127096 6016
rect 127160 5952 127176 6016
rect 127240 5952 127256 6016
rect 127320 5952 127336 6016
rect 127400 5952 127406 6016
rect 127090 5951 127406 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 81010 5472 81326 5473
rect 81010 5408 81016 5472
rect 81080 5408 81096 5472
rect 81160 5408 81176 5472
rect 81240 5408 81256 5472
rect 81320 5408 81326 5472
rect 81010 5407 81326 5408
rect 111730 5472 112046 5473
rect 111730 5408 111736 5472
rect 111800 5408 111816 5472
rect 111880 5408 111896 5472
rect 111960 5408 111976 5472
rect 112040 5408 112046 5472
rect 111730 5407 112046 5408
rect 142450 5472 142766 5473
rect 142450 5408 142456 5472
rect 142520 5408 142536 5472
rect 142600 5408 142616 5472
rect 142680 5408 142696 5472
rect 142760 5408 142766 5472
rect 142450 5407 142766 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 65650 4928 65966 4929
rect 65650 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65966 4928
rect 65650 4863 65966 4864
rect 96370 4928 96686 4929
rect 96370 4864 96376 4928
rect 96440 4864 96456 4928
rect 96520 4864 96536 4928
rect 96600 4864 96616 4928
rect 96680 4864 96686 4928
rect 96370 4863 96686 4864
rect 127090 4928 127406 4929
rect 127090 4864 127096 4928
rect 127160 4864 127176 4928
rect 127240 4864 127256 4928
rect 127320 4864 127336 4928
rect 127400 4864 127406 4928
rect 127090 4863 127406 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 81010 4384 81326 4385
rect 81010 4320 81016 4384
rect 81080 4320 81096 4384
rect 81160 4320 81176 4384
rect 81240 4320 81256 4384
rect 81320 4320 81326 4384
rect 81010 4319 81326 4320
rect 111730 4384 112046 4385
rect 111730 4320 111736 4384
rect 111800 4320 111816 4384
rect 111880 4320 111896 4384
rect 111960 4320 111976 4384
rect 112040 4320 112046 4384
rect 111730 4319 112046 4320
rect 142450 4384 142766 4385
rect 142450 4320 142456 4384
rect 142520 4320 142536 4384
rect 142600 4320 142616 4384
rect 142680 4320 142696 4384
rect 142760 4320 142766 4384
rect 142450 4319 142766 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 65650 3840 65966 3841
rect 65650 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65966 3840
rect 65650 3775 65966 3776
rect 96370 3840 96686 3841
rect 96370 3776 96376 3840
rect 96440 3776 96456 3840
rect 96520 3776 96536 3840
rect 96600 3776 96616 3840
rect 96680 3776 96686 3840
rect 96370 3775 96686 3776
rect 127090 3840 127406 3841
rect 127090 3776 127096 3840
rect 127160 3776 127176 3840
rect 127240 3776 127256 3840
rect 127320 3776 127336 3840
rect 127400 3776 127406 3840
rect 127090 3775 127406 3776
rect 22001 3634 22067 3637
rect 28073 3634 28139 3637
rect 22001 3632 28139 3634
rect 22001 3576 22006 3632
rect 22062 3576 28078 3632
rect 28134 3576 28139 3632
rect 22001 3574 28139 3576
rect 22001 3571 22067 3574
rect 28073 3571 28139 3574
rect 81341 3634 81407 3637
rect 83273 3634 83339 3637
rect 81341 3632 83339 3634
rect 81341 3576 81346 3632
rect 81402 3576 83278 3632
rect 83334 3576 83339 3632
rect 81341 3574 83339 3576
rect 81341 3571 81407 3574
rect 83273 3571 83339 3574
rect 68461 3498 68527 3501
rect 71221 3498 71287 3501
rect 68461 3496 71287 3498
rect 68461 3440 68466 3496
rect 68522 3440 71226 3496
rect 71282 3440 71287 3496
rect 68461 3438 71287 3440
rect 68461 3435 68527 3438
rect 71221 3435 71287 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 81010 3296 81326 3297
rect 81010 3232 81016 3296
rect 81080 3232 81096 3296
rect 81160 3232 81176 3296
rect 81240 3232 81256 3296
rect 81320 3232 81326 3296
rect 81010 3231 81326 3232
rect 111730 3296 112046 3297
rect 111730 3232 111736 3296
rect 111800 3232 111816 3296
rect 111880 3232 111896 3296
rect 111960 3232 111976 3296
rect 112040 3232 112046 3296
rect 111730 3231 112046 3232
rect 142450 3296 142766 3297
rect 142450 3232 142456 3296
rect 142520 3232 142536 3296
rect 142600 3232 142616 3296
rect 142680 3232 142696 3296
rect 142760 3232 142766 3296
rect 142450 3231 142766 3232
rect 41689 2954 41755 2957
rect 42609 2954 42675 2957
rect 41689 2952 42675 2954
rect 41689 2896 41694 2952
rect 41750 2896 42614 2952
rect 42670 2896 42675 2952
rect 41689 2894 42675 2896
rect 41689 2891 41755 2894
rect 42609 2891 42675 2894
rect 69933 2954 69999 2957
rect 75729 2954 75795 2957
rect 69933 2952 75795 2954
rect 69933 2896 69938 2952
rect 69994 2896 75734 2952
rect 75790 2896 75795 2952
rect 69933 2894 75795 2896
rect 69933 2891 69999 2894
rect 75729 2891 75795 2894
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 65650 2752 65966 2753
rect 65650 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65966 2752
rect 65650 2687 65966 2688
rect 96370 2752 96686 2753
rect 96370 2688 96376 2752
rect 96440 2688 96456 2752
rect 96520 2688 96536 2752
rect 96600 2688 96616 2752
rect 96680 2688 96686 2752
rect 96370 2687 96686 2688
rect 127090 2752 127406 2753
rect 127090 2688 127096 2752
rect 127160 2688 127176 2752
rect 127240 2688 127256 2752
rect 127320 2688 127336 2752
rect 127400 2688 127406 2752
rect 127090 2687 127406 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
rect 81010 2208 81326 2209
rect 81010 2144 81016 2208
rect 81080 2144 81096 2208
rect 81160 2144 81176 2208
rect 81240 2144 81256 2208
rect 81320 2144 81326 2208
rect 81010 2143 81326 2144
rect 111730 2208 112046 2209
rect 111730 2144 111736 2208
rect 111800 2144 111816 2208
rect 111880 2144 111896 2208
rect 111960 2144 111976 2208
rect 112040 2144 112046 2208
rect 111730 2143 112046 2144
rect 142450 2208 142766 2209
rect 142450 2144 142456 2208
rect 142520 2144 142536 2208
rect 142600 2144 142616 2208
rect 142680 2144 142696 2208
rect 142760 2144 142766 2208
rect 142450 2143 142766 2144
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 65656 37564 65720 37568
rect 65656 37508 65660 37564
rect 65660 37508 65716 37564
rect 65716 37508 65720 37564
rect 65656 37504 65720 37508
rect 65736 37564 65800 37568
rect 65736 37508 65740 37564
rect 65740 37508 65796 37564
rect 65796 37508 65800 37564
rect 65736 37504 65800 37508
rect 65816 37564 65880 37568
rect 65816 37508 65820 37564
rect 65820 37508 65876 37564
rect 65876 37508 65880 37564
rect 65816 37504 65880 37508
rect 65896 37564 65960 37568
rect 65896 37508 65900 37564
rect 65900 37508 65956 37564
rect 65956 37508 65960 37564
rect 65896 37504 65960 37508
rect 96376 37564 96440 37568
rect 96376 37508 96380 37564
rect 96380 37508 96436 37564
rect 96436 37508 96440 37564
rect 96376 37504 96440 37508
rect 96456 37564 96520 37568
rect 96456 37508 96460 37564
rect 96460 37508 96516 37564
rect 96516 37508 96520 37564
rect 96456 37504 96520 37508
rect 96536 37564 96600 37568
rect 96536 37508 96540 37564
rect 96540 37508 96596 37564
rect 96596 37508 96600 37564
rect 96536 37504 96600 37508
rect 96616 37564 96680 37568
rect 96616 37508 96620 37564
rect 96620 37508 96676 37564
rect 96676 37508 96680 37564
rect 96616 37504 96680 37508
rect 127096 37564 127160 37568
rect 127096 37508 127100 37564
rect 127100 37508 127156 37564
rect 127156 37508 127160 37564
rect 127096 37504 127160 37508
rect 127176 37564 127240 37568
rect 127176 37508 127180 37564
rect 127180 37508 127236 37564
rect 127236 37508 127240 37564
rect 127176 37504 127240 37508
rect 127256 37564 127320 37568
rect 127256 37508 127260 37564
rect 127260 37508 127316 37564
rect 127316 37508 127320 37564
rect 127256 37504 127320 37508
rect 127336 37564 127400 37568
rect 127336 37508 127340 37564
rect 127340 37508 127396 37564
rect 127396 37508 127400 37564
rect 127336 37504 127400 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 81016 37020 81080 37024
rect 81016 36964 81020 37020
rect 81020 36964 81076 37020
rect 81076 36964 81080 37020
rect 81016 36960 81080 36964
rect 81096 37020 81160 37024
rect 81096 36964 81100 37020
rect 81100 36964 81156 37020
rect 81156 36964 81160 37020
rect 81096 36960 81160 36964
rect 81176 37020 81240 37024
rect 81176 36964 81180 37020
rect 81180 36964 81236 37020
rect 81236 36964 81240 37020
rect 81176 36960 81240 36964
rect 81256 37020 81320 37024
rect 81256 36964 81260 37020
rect 81260 36964 81316 37020
rect 81316 36964 81320 37020
rect 81256 36960 81320 36964
rect 111736 37020 111800 37024
rect 111736 36964 111740 37020
rect 111740 36964 111796 37020
rect 111796 36964 111800 37020
rect 111736 36960 111800 36964
rect 111816 37020 111880 37024
rect 111816 36964 111820 37020
rect 111820 36964 111876 37020
rect 111876 36964 111880 37020
rect 111816 36960 111880 36964
rect 111896 37020 111960 37024
rect 111896 36964 111900 37020
rect 111900 36964 111956 37020
rect 111956 36964 111960 37020
rect 111896 36960 111960 36964
rect 111976 37020 112040 37024
rect 111976 36964 111980 37020
rect 111980 36964 112036 37020
rect 112036 36964 112040 37020
rect 111976 36960 112040 36964
rect 142456 37020 142520 37024
rect 142456 36964 142460 37020
rect 142460 36964 142516 37020
rect 142516 36964 142520 37020
rect 142456 36960 142520 36964
rect 142536 37020 142600 37024
rect 142536 36964 142540 37020
rect 142540 36964 142596 37020
rect 142596 36964 142600 37020
rect 142536 36960 142600 36964
rect 142616 37020 142680 37024
rect 142616 36964 142620 37020
rect 142620 36964 142676 37020
rect 142676 36964 142680 37020
rect 142616 36960 142680 36964
rect 142696 37020 142760 37024
rect 142696 36964 142700 37020
rect 142700 36964 142756 37020
rect 142756 36964 142760 37020
rect 142696 36960 142760 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 65656 36476 65720 36480
rect 65656 36420 65660 36476
rect 65660 36420 65716 36476
rect 65716 36420 65720 36476
rect 65656 36416 65720 36420
rect 65736 36476 65800 36480
rect 65736 36420 65740 36476
rect 65740 36420 65796 36476
rect 65796 36420 65800 36476
rect 65736 36416 65800 36420
rect 65816 36476 65880 36480
rect 65816 36420 65820 36476
rect 65820 36420 65876 36476
rect 65876 36420 65880 36476
rect 65816 36416 65880 36420
rect 65896 36476 65960 36480
rect 65896 36420 65900 36476
rect 65900 36420 65956 36476
rect 65956 36420 65960 36476
rect 65896 36416 65960 36420
rect 96376 36476 96440 36480
rect 96376 36420 96380 36476
rect 96380 36420 96436 36476
rect 96436 36420 96440 36476
rect 96376 36416 96440 36420
rect 96456 36476 96520 36480
rect 96456 36420 96460 36476
rect 96460 36420 96516 36476
rect 96516 36420 96520 36476
rect 96456 36416 96520 36420
rect 96536 36476 96600 36480
rect 96536 36420 96540 36476
rect 96540 36420 96596 36476
rect 96596 36420 96600 36476
rect 96536 36416 96600 36420
rect 96616 36476 96680 36480
rect 96616 36420 96620 36476
rect 96620 36420 96676 36476
rect 96676 36420 96680 36476
rect 96616 36416 96680 36420
rect 127096 36476 127160 36480
rect 127096 36420 127100 36476
rect 127100 36420 127156 36476
rect 127156 36420 127160 36476
rect 127096 36416 127160 36420
rect 127176 36476 127240 36480
rect 127176 36420 127180 36476
rect 127180 36420 127236 36476
rect 127236 36420 127240 36476
rect 127176 36416 127240 36420
rect 127256 36476 127320 36480
rect 127256 36420 127260 36476
rect 127260 36420 127316 36476
rect 127316 36420 127320 36476
rect 127256 36416 127320 36420
rect 127336 36476 127400 36480
rect 127336 36420 127340 36476
rect 127340 36420 127396 36476
rect 127396 36420 127400 36476
rect 127336 36416 127400 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 81016 35932 81080 35936
rect 81016 35876 81020 35932
rect 81020 35876 81076 35932
rect 81076 35876 81080 35932
rect 81016 35872 81080 35876
rect 81096 35932 81160 35936
rect 81096 35876 81100 35932
rect 81100 35876 81156 35932
rect 81156 35876 81160 35932
rect 81096 35872 81160 35876
rect 81176 35932 81240 35936
rect 81176 35876 81180 35932
rect 81180 35876 81236 35932
rect 81236 35876 81240 35932
rect 81176 35872 81240 35876
rect 81256 35932 81320 35936
rect 81256 35876 81260 35932
rect 81260 35876 81316 35932
rect 81316 35876 81320 35932
rect 81256 35872 81320 35876
rect 111736 35932 111800 35936
rect 111736 35876 111740 35932
rect 111740 35876 111796 35932
rect 111796 35876 111800 35932
rect 111736 35872 111800 35876
rect 111816 35932 111880 35936
rect 111816 35876 111820 35932
rect 111820 35876 111876 35932
rect 111876 35876 111880 35932
rect 111816 35872 111880 35876
rect 111896 35932 111960 35936
rect 111896 35876 111900 35932
rect 111900 35876 111956 35932
rect 111956 35876 111960 35932
rect 111896 35872 111960 35876
rect 111976 35932 112040 35936
rect 111976 35876 111980 35932
rect 111980 35876 112036 35932
rect 112036 35876 112040 35932
rect 111976 35872 112040 35876
rect 142456 35932 142520 35936
rect 142456 35876 142460 35932
rect 142460 35876 142516 35932
rect 142516 35876 142520 35932
rect 142456 35872 142520 35876
rect 142536 35932 142600 35936
rect 142536 35876 142540 35932
rect 142540 35876 142596 35932
rect 142596 35876 142600 35932
rect 142536 35872 142600 35876
rect 142616 35932 142680 35936
rect 142616 35876 142620 35932
rect 142620 35876 142676 35932
rect 142676 35876 142680 35932
rect 142616 35872 142680 35876
rect 142696 35932 142760 35936
rect 142696 35876 142700 35932
rect 142700 35876 142756 35932
rect 142756 35876 142760 35932
rect 142696 35872 142760 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 65656 35388 65720 35392
rect 65656 35332 65660 35388
rect 65660 35332 65716 35388
rect 65716 35332 65720 35388
rect 65656 35328 65720 35332
rect 65736 35388 65800 35392
rect 65736 35332 65740 35388
rect 65740 35332 65796 35388
rect 65796 35332 65800 35388
rect 65736 35328 65800 35332
rect 65816 35388 65880 35392
rect 65816 35332 65820 35388
rect 65820 35332 65876 35388
rect 65876 35332 65880 35388
rect 65816 35328 65880 35332
rect 65896 35388 65960 35392
rect 65896 35332 65900 35388
rect 65900 35332 65956 35388
rect 65956 35332 65960 35388
rect 65896 35328 65960 35332
rect 96376 35388 96440 35392
rect 96376 35332 96380 35388
rect 96380 35332 96436 35388
rect 96436 35332 96440 35388
rect 96376 35328 96440 35332
rect 96456 35388 96520 35392
rect 96456 35332 96460 35388
rect 96460 35332 96516 35388
rect 96516 35332 96520 35388
rect 96456 35328 96520 35332
rect 96536 35388 96600 35392
rect 96536 35332 96540 35388
rect 96540 35332 96596 35388
rect 96596 35332 96600 35388
rect 96536 35328 96600 35332
rect 96616 35388 96680 35392
rect 96616 35332 96620 35388
rect 96620 35332 96676 35388
rect 96676 35332 96680 35388
rect 96616 35328 96680 35332
rect 127096 35388 127160 35392
rect 127096 35332 127100 35388
rect 127100 35332 127156 35388
rect 127156 35332 127160 35388
rect 127096 35328 127160 35332
rect 127176 35388 127240 35392
rect 127176 35332 127180 35388
rect 127180 35332 127236 35388
rect 127236 35332 127240 35388
rect 127176 35328 127240 35332
rect 127256 35388 127320 35392
rect 127256 35332 127260 35388
rect 127260 35332 127316 35388
rect 127316 35332 127320 35388
rect 127256 35328 127320 35332
rect 127336 35388 127400 35392
rect 127336 35332 127340 35388
rect 127340 35332 127396 35388
rect 127396 35332 127400 35388
rect 127336 35328 127400 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 81016 34844 81080 34848
rect 81016 34788 81020 34844
rect 81020 34788 81076 34844
rect 81076 34788 81080 34844
rect 81016 34784 81080 34788
rect 81096 34844 81160 34848
rect 81096 34788 81100 34844
rect 81100 34788 81156 34844
rect 81156 34788 81160 34844
rect 81096 34784 81160 34788
rect 81176 34844 81240 34848
rect 81176 34788 81180 34844
rect 81180 34788 81236 34844
rect 81236 34788 81240 34844
rect 81176 34784 81240 34788
rect 81256 34844 81320 34848
rect 81256 34788 81260 34844
rect 81260 34788 81316 34844
rect 81316 34788 81320 34844
rect 81256 34784 81320 34788
rect 111736 34844 111800 34848
rect 111736 34788 111740 34844
rect 111740 34788 111796 34844
rect 111796 34788 111800 34844
rect 111736 34784 111800 34788
rect 111816 34844 111880 34848
rect 111816 34788 111820 34844
rect 111820 34788 111876 34844
rect 111876 34788 111880 34844
rect 111816 34784 111880 34788
rect 111896 34844 111960 34848
rect 111896 34788 111900 34844
rect 111900 34788 111956 34844
rect 111956 34788 111960 34844
rect 111896 34784 111960 34788
rect 111976 34844 112040 34848
rect 111976 34788 111980 34844
rect 111980 34788 112036 34844
rect 112036 34788 112040 34844
rect 111976 34784 112040 34788
rect 142456 34844 142520 34848
rect 142456 34788 142460 34844
rect 142460 34788 142516 34844
rect 142516 34788 142520 34844
rect 142456 34784 142520 34788
rect 142536 34844 142600 34848
rect 142536 34788 142540 34844
rect 142540 34788 142596 34844
rect 142596 34788 142600 34844
rect 142536 34784 142600 34788
rect 142616 34844 142680 34848
rect 142616 34788 142620 34844
rect 142620 34788 142676 34844
rect 142676 34788 142680 34844
rect 142616 34784 142680 34788
rect 142696 34844 142760 34848
rect 142696 34788 142700 34844
rect 142700 34788 142756 34844
rect 142756 34788 142760 34844
rect 142696 34784 142760 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 65656 34300 65720 34304
rect 65656 34244 65660 34300
rect 65660 34244 65716 34300
rect 65716 34244 65720 34300
rect 65656 34240 65720 34244
rect 65736 34300 65800 34304
rect 65736 34244 65740 34300
rect 65740 34244 65796 34300
rect 65796 34244 65800 34300
rect 65736 34240 65800 34244
rect 65816 34300 65880 34304
rect 65816 34244 65820 34300
rect 65820 34244 65876 34300
rect 65876 34244 65880 34300
rect 65816 34240 65880 34244
rect 65896 34300 65960 34304
rect 65896 34244 65900 34300
rect 65900 34244 65956 34300
rect 65956 34244 65960 34300
rect 65896 34240 65960 34244
rect 96376 34300 96440 34304
rect 96376 34244 96380 34300
rect 96380 34244 96436 34300
rect 96436 34244 96440 34300
rect 96376 34240 96440 34244
rect 96456 34300 96520 34304
rect 96456 34244 96460 34300
rect 96460 34244 96516 34300
rect 96516 34244 96520 34300
rect 96456 34240 96520 34244
rect 96536 34300 96600 34304
rect 96536 34244 96540 34300
rect 96540 34244 96596 34300
rect 96596 34244 96600 34300
rect 96536 34240 96600 34244
rect 96616 34300 96680 34304
rect 96616 34244 96620 34300
rect 96620 34244 96676 34300
rect 96676 34244 96680 34300
rect 96616 34240 96680 34244
rect 127096 34300 127160 34304
rect 127096 34244 127100 34300
rect 127100 34244 127156 34300
rect 127156 34244 127160 34300
rect 127096 34240 127160 34244
rect 127176 34300 127240 34304
rect 127176 34244 127180 34300
rect 127180 34244 127236 34300
rect 127236 34244 127240 34300
rect 127176 34240 127240 34244
rect 127256 34300 127320 34304
rect 127256 34244 127260 34300
rect 127260 34244 127316 34300
rect 127316 34244 127320 34300
rect 127256 34240 127320 34244
rect 127336 34300 127400 34304
rect 127336 34244 127340 34300
rect 127340 34244 127396 34300
rect 127396 34244 127400 34300
rect 127336 34240 127400 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 81016 33756 81080 33760
rect 81016 33700 81020 33756
rect 81020 33700 81076 33756
rect 81076 33700 81080 33756
rect 81016 33696 81080 33700
rect 81096 33756 81160 33760
rect 81096 33700 81100 33756
rect 81100 33700 81156 33756
rect 81156 33700 81160 33756
rect 81096 33696 81160 33700
rect 81176 33756 81240 33760
rect 81176 33700 81180 33756
rect 81180 33700 81236 33756
rect 81236 33700 81240 33756
rect 81176 33696 81240 33700
rect 81256 33756 81320 33760
rect 81256 33700 81260 33756
rect 81260 33700 81316 33756
rect 81316 33700 81320 33756
rect 81256 33696 81320 33700
rect 111736 33756 111800 33760
rect 111736 33700 111740 33756
rect 111740 33700 111796 33756
rect 111796 33700 111800 33756
rect 111736 33696 111800 33700
rect 111816 33756 111880 33760
rect 111816 33700 111820 33756
rect 111820 33700 111876 33756
rect 111876 33700 111880 33756
rect 111816 33696 111880 33700
rect 111896 33756 111960 33760
rect 111896 33700 111900 33756
rect 111900 33700 111956 33756
rect 111956 33700 111960 33756
rect 111896 33696 111960 33700
rect 111976 33756 112040 33760
rect 111976 33700 111980 33756
rect 111980 33700 112036 33756
rect 112036 33700 112040 33756
rect 111976 33696 112040 33700
rect 142456 33756 142520 33760
rect 142456 33700 142460 33756
rect 142460 33700 142516 33756
rect 142516 33700 142520 33756
rect 142456 33696 142520 33700
rect 142536 33756 142600 33760
rect 142536 33700 142540 33756
rect 142540 33700 142596 33756
rect 142596 33700 142600 33756
rect 142536 33696 142600 33700
rect 142616 33756 142680 33760
rect 142616 33700 142620 33756
rect 142620 33700 142676 33756
rect 142676 33700 142680 33756
rect 142616 33696 142680 33700
rect 142696 33756 142760 33760
rect 142696 33700 142700 33756
rect 142700 33700 142756 33756
rect 142756 33700 142760 33756
rect 142696 33696 142760 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 65656 33212 65720 33216
rect 65656 33156 65660 33212
rect 65660 33156 65716 33212
rect 65716 33156 65720 33212
rect 65656 33152 65720 33156
rect 65736 33212 65800 33216
rect 65736 33156 65740 33212
rect 65740 33156 65796 33212
rect 65796 33156 65800 33212
rect 65736 33152 65800 33156
rect 65816 33212 65880 33216
rect 65816 33156 65820 33212
rect 65820 33156 65876 33212
rect 65876 33156 65880 33212
rect 65816 33152 65880 33156
rect 65896 33212 65960 33216
rect 65896 33156 65900 33212
rect 65900 33156 65956 33212
rect 65956 33156 65960 33212
rect 65896 33152 65960 33156
rect 96376 33212 96440 33216
rect 96376 33156 96380 33212
rect 96380 33156 96436 33212
rect 96436 33156 96440 33212
rect 96376 33152 96440 33156
rect 96456 33212 96520 33216
rect 96456 33156 96460 33212
rect 96460 33156 96516 33212
rect 96516 33156 96520 33212
rect 96456 33152 96520 33156
rect 96536 33212 96600 33216
rect 96536 33156 96540 33212
rect 96540 33156 96596 33212
rect 96596 33156 96600 33212
rect 96536 33152 96600 33156
rect 96616 33212 96680 33216
rect 96616 33156 96620 33212
rect 96620 33156 96676 33212
rect 96676 33156 96680 33212
rect 96616 33152 96680 33156
rect 127096 33212 127160 33216
rect 127096 33156 127100 33212
rect 127100 33156 127156 33212
rect 127156 33156 127160 33212
rect 127096 33152 127160 33156
rect 127176 33212 127240 33216
rect 127176 33156 127180 33212
rect 127180 33156 127236 33212
rect 127236 33156 127240 33212
rect 127176 33152 127240 33156
rect 127256 33212 127320 33216
rect 127256 33156 127260 33212
rect 127260 33156 127316 33212
rect 127316 33156 127320 33212
rect 127256 33152 127320 33156
rect 127336 33212 127400 33216
rect 127336 33156 127340 33212
rect 127340 33156 127396 33212
rect 127396 33156 127400 33212
rect 127336 33152 127400 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 81016 32668 81080 32672
rect 81016 32612 81020 32668
rect 81020 32612 81076 32668
rect 81076 32612 81080 32668
rect 81016 32608 81080 32612
rect 81096 32668 81160 32672
rect 81096 32612 81100 32668
rect 81100 32612 81156 32668
rect 81156 32612 81160 32668
rect 81096 32608 81160 32612
rect 81176 32668 81240 32672
rect 81176 32612 81180 32668
rect 81180 32612 81236 32668
rect 81236 32612 81240 32668
rect 81176 32608 81240 32612
rect 81256 32668 81320 32672
rect 81256 32612 81260 32668
rect 81260 32612 81316 32668
rect 81316 32612 81320 32668
rect 81256 32608 81320 32612
rect 111736 32668 111800 32672
rect 111736 32612 111740 32668
rect 111740 32612 111796 32668
rect 111796 32612 111800 32668
rect 111736 32608 111800 32612
rect 111816 32668 111880 32672
rect 111816 32612 111820 32668
rect 111820 32612 111876 32668
rect 111876 32612 111880 32668
rect 111816 32608 111880 32612
rect 111896 32668 111960 32672
rect 111896 32612 111900 32668
rect 111900 32612 111956 32668
rect 111956 32612 111960 32668
rect 111896 32608 111960 32612
rect 111976 32668 112040 32672
rect 111976 32612 111980 32668
rect 111980 32612 112036 32668
rect 112036 32612 112040 32668
rect 111976 32608 112040 32612
rect 142456 32668 142520 32672
rect 142456 32612 142460 32668
rect 142460 32612 142516 32668
rect 142516 32612 142520 32668
rect 142456 32608 142520 32612
rect 142536 32668 142600 32672
rect 142536 32612 142540 32668
rect 142540 32612 142596 32668
rect 142596 32612 142600 32668
rect 142536 32608 142600 32612
rect 142616 32668 142680 32672
rect 142616 32612 142620 32668
rect 142620 32612 142676 32668
rect 142676 32612 142680 32668
rect 142616 32608 142680 32612
rect 142696 32668 142760 32672
rect 142696 32612 142700 32668
rect 142700 32612 142756 32668
rect 142756 32612 142760 32668
rect 142696 32608 142760 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 65656 32124 65720 32128
rect 65656 32068 65660 32124
rect 65660 32068 65716 32124
rect 65716 32068 65720 32124
rect 65656 32064 65720 32068
rect 65736 32124 65800 32128
rect 65736 32068 65740 32124
rect 65740 32068 65796 32124
rect 65796 32068 65800 32124
rect 65736 32064 65800 32068
rect 65816 32124 65880 32128
rect 65816 32068 65820 32124
rect 65820 32068 65876 32124
rect 65876 32068 65880 32124
rect 65816 32064 65880 32068
rect 65896 32124 65960 32128
rect 65896 32068 65900 32124
rect 65900 32068 65956 32124
rect 65956 32068 65960 32124
rect 65896 32064 65960 32068
rect 96376 32124 96440 32128
rect 96376 32068 96380 32124
rect 96380 32068 96436 32124
rect 96436 32068 96440 32124
rect 96376 32064 96440 32068
rect 96456 32124 96520 32128
rect 96456 32068 96460 32124
rect 96460 32068 96516 32124
rect 96516 32068 96520 32124
rect 96456 32064 96520 32068
rect 96536 32124 96600 32128
rect 96536 32068 96540 32124
rect 96540 32068 96596 32124
rect 96596 32068 96600 32124
rect 96536 32064 96600 32068
rect 96616 32124 96680 32128
rect 96616 32068 96620 32124
rect 96620 32068 96676 32124
rect 96676 32068 96680 32124
rect 96616 32064 96680 32068
rect 127096 32124 127160 32128
rect 127096 32068 127100 32124
rect 127100 32068 127156 32124
rect 127156 32068 127160 32124
rect 127096 32064 127160 32068
rect 127176 32124 127240 32128
rect 127176 32068 127180 32124
rect 127180 32068 127236 32124
rect 127236 32068 127240 32124
rect 127176 32064 127240 32068
rect 127256 32124 127320 32128
rect 127256 32068 127260 32124
rect 127260 32068 127316 32124
rect 127316 32068 127320 32124
rect 127256 32064 127320 32068
rect 127336 32124 127400 32128
rect 127336 32068 127340 32124
rect 127340 32068 127396 32124
rect 127396 32068 127400 32124
rect 127336 32064 127400 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 81016 31580 81080 31584
rect 81016 31524 81020 31580
rect 81020 31524 81076 31580
rect 81076 31524 81080 31580
rect 81016 31520 81080 31524
rect 81096 31580 81160 31584
rect 81096 31524 81100 31580
rect 81100 31524 81156 31580
rect 81156 31524 81160 31580
rect 81096 31520 81160 31524
rect 81176 31580 81240 31584
rect 81176 31524 81180 31580
rect 81180 31524 81236 31580
rect 81236 31524 81240 31580
rect 81176 31520 81240 31524
rect 81256 31580 81320 31584
rect 81256 31524 81260 31580
rect 81260 31524 81316 31580
rect 81316 31524 81320 31580
rect 81256 31520 81320 31524
rect 111736 31580 111800 31584
rect 111736 31524 111740 31580
rect 111740 31524 111796 31580
rect 111796 31524 111800 31580
rect 111736 31520 111800 31524
rect 111816 31580 111880 31584
rect 111816 31524 111820 31580
rect 111820 31524 111876 31580
rect 111876 31524 111880 31580
rect 111816 31520 111880 31524
rect 111896 31580 111960 31584
rect 111896 31524 111900 31580
rect 111900 31524 111956 31580
rect 111956 31524 111960 31580
rect 111896 31520 111960 31524
rect 111976 31580 112040 31584
rect 111976 31524 111980 31580
rect 111980 31524 112036 31580
rect 112036 31524 112040 31580
rect 111976 31520 112040 31524
rect 142456 31580 142520 31584
rect 142456 31524 142460 31580
rect 142460 31524 142516 31580
rect 142516 31524 142520 31580
rect 142456 31520 142520 31524
rect 142536 31580 142600 31584
rect 142536 31524 142540 31580
rect 142540 31524 142596 31580
rect 142596 31524 142600 31580
rect 142536 31520 142600 31524
rect 142616 31580 142680 31584
rect 142616 31524 142620 31580
rect 142620 31524 142676 31580
rect 142676 31524 142680 31580
rect 142616 31520 142680 31524
rect 142696 31580 142760 31584
rect 142696 31524 142700 31580
rect 142700 31524 142756 31580
rect 142756 31524 142760 31580
rect 142696 31520 142760 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 65656 31036 65720 31040
rect 65656 30980 65660 31036
rect 65660 30980 65716 31036
rect 65716 30980 65720 31036
rect 65656 30976 65720 30980
rect 65736 31036 65800 31040
rect 65736 30980 65740 31036
rect 65740 30980 65796 31036
rect 65796 30980 65800 31036
rect 65736 30976 65800 30980
rect 65816 31036 65880 31040
rect 65816 30980 65820 31036
rect 65820 30980 65876 31036
rect 65876 30980 65880 31036
rect 65816 30976 65880 30980
rect 65896 31036 65960 31040
rect 65896 30980 65900 31036
rect 65900 30980 65956 31036
rect 65956 30980 65960 31036
rect 65896 30976 65960 30980
rect 96376 31036 96440 31040
rect 96376 30980 96380 31036
rect 96380 30980 96436 31036
rect 96436 30980 96440 31036
rect 96376 30976 96440 30980
rect 96456 31036 96520 31040
rect 96456 30980 96460 31036
rect 96460 30980 96516 31036
rect 96516 30980 96520 31036
rect 96456 30976 96520 30980
rect 96536 31036 96600 31040
rect 96536 30980 96540 31036
rect 96540 30980 96596 31036
rect 96596 30980 96600 31036
rect 96536 30976 96600 30980
rect 96616 31036 96680 31040
rect 96616 30980 96620 31036
rect 96620 30980 96676 31036
rect 96676 30980 96680 31036
rect 96616 30976 96680 30980
rect 127096 31036 127160 31040
rect 127096 30980 127100 31036
rect 127100 30980 127156 31036
rect 127156 30980 127160 31036
rect 127096 30976 127160 30980
rect 127176 31036 127240 31040
rect 127176 30980 127180 31036
rect 127180 30980 127236 31036
rect 127236 30980 127240 31036
rect 127176 30976 127240 30980
rect 127256 31036 127320 31040
rect 127256 30980 127260 31036
rect 127260 30980 127316 31036
rect 127316 30980 127320 31036
rect 127256 30976 127320 30980
rect 127336 31036 127400 31040
rect 127336 30980 127340 31036
rect 127340 30980 127396 31036
rect 127396 30980 127400 31036
rect 127336 30976 127400 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 81016 30492 81080 30496
rect 81016 30436 81020 30492
rect 81020 30436 81076 30492
rect 81076 30436 81080 30492
rect 81016 30432 81080 30436
rect 81096 30492 81160 30496
rect 81096 30436 81100 30492
rect 81100 30436 81156 30492
rect 81156 30436 81160 30492
rect 81096 30432 81160 30436
rect 81176 30492 81240 30496
rect 81176 30436 81180 30492
rect 81180 30436 81236 30492
rect 81236 30436 81240 30492
rect 81176 30432 81240 30436
rect 81256 30492 81320 30496
rect 81256 30436 81260 30492
rect 81260 30436 81316 30492
rect 81316 30436 81320 30492
rect 81256 30432 81320 30436
rect 111736 30492 111800 30496
rect 111736 30436 111740 30492
rect 111740 30436 111796 30492
rect 111796 30436 111800 30492
rect 111736 30432 111800 30436
rect 111816 30492 111880 30496
rect 111816 30436 111820 30492
rect 111820 30436 111876 30492
rect 111876 30436 111880 30492
rect 111816 30432 111880 30436
rect 111896 30492 111960 30496
rect 111896 30436 111900 30492
rect 111900 30436 111956 30492
rect 111956 30436 111960 30492
rect 111896 30432 111960 30436
rect 111976 30492 112040 30496
rect 111976 30436 111980 30492
rect 111980 30436 112036 30492
rect 112036 30436 112040 30492
rect 111976 30432 112040 30436
rect 142456 30492 142520 30496
rect 142456 30436 142460 30492
rect 142460 30436 142516 30492
rect 142516 30436 142520 30492
rect 142456 30432 142520 30436
rect 142536 30492 142600 30496
rect 142536 30436 142540 30492
rect 142540 30436 142596 30492
rect 142596 30436 142600 30492
rect 142536 30432 142600 30436
rect 142616 30492 142680 30496
rect 142616 30436 142620 30492
rect 142620 30436 142676 30492
rect 142676 30436 142680 30492
rect 142616 30432 142680 30436
rect 142696 30492 142760 30496
rect 142696 30436 142700 30492
rect 142700 30436 142756 30492
rect 142756 30436 142760 30492
rect 142696 30432 142760 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 65656 29948 65720 29952
rect 65656 29892 65660 29948
rect 65660 29892 65716 29948
rect 65716 29892 65720 29948
rect 65656 29888 65720 29892
rect 65736 29948 65800 29952
rect 65736 29892 65740 29948
rect 65740 29892 65796 29948
rect 65796 29892 65800 29948
rect 65736 29888 65800 29892
rect 65816 29948 65880 29952
rect 65816 29892 65820 29948
rect 65820 29892 65876 29948
rect 65876 29892 65880 29948
rect 65816 29888 65880 29892
rect 65896 29948 65960 29952
rect 65896 29892 65900 29948
rect 65900 29892 65956 29948
rect 65956 29892 65960 29948
rect 65896 29888 65960 29892
rect 96376 29948 96440 29952
rect 96376 29892 96380 29948
rect 96380 29892 96436 29948
rect 96436 29892 96440 29948
rect 96376 29888 96440 29892
rect 96456 29948 96520 29952
rect 96456 29892 96460 29948
rect 96460 29892 96516 29948
rect 96516 29892 96520 29948
rect 96456 29888 96520 29892
rect 96536 29948 96600 29952
rect 96536 29892 96540 29948
rect 96540 29892 96596 29948
rect 96596 29892 96600 29948
rect 96536 29888 96600 29892
rect 96616 29948 96680 29952
rect 96616 29892 96620 29948
rect 96620 29892 96676 29948
rect 96676 29892 96680 29948
rect 96616 29888 96680 29892
rect 127096 29948 127160 29952
rect 127096 29892 127100 29948
rect 127100 29892 127156 29948
rect 127156 29892 127160 29948
rect 127096 29888 127160 29892
rect 127176 29948 127240 29952
rect 127176 29892 127180 29948
rect 127180 29892 127236 29948
rect 127236 29892 127240 29948
rect 127176 29888 127240 29892
rect 127256 29948 127320 29952
rect 127256 29892 127260 29948
rect 127260 29892 127316 29948
rect 127316 29892 127320 29948
rect 127256 29888 127320 29892
rect 127336 29948 127400 29952
rect 127336 29892 127340 29948
rect 127340 29892 127396 29948
rect 127396 29892 127400 29948
rect 127336 29888 127400 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 81016 29404 81080 29408
rect 81016 29348 81020 29404
rect 81020 29348 81076 29404
rect 81076 29348 81080 29404
rect 81016 29344 81080 29348
rect 81096 29404 81160 29408
rect 81096 29348 81100 29404
rect 81100 29348 81156 29404
rect 81156 29348 81160 29404
rect 81096 29344 81160 29348
rect 81176 29404 81240 29408
rect 81176 29348 81180 29404
rect 81180 29348 81236 29404
rect 81236 29348 81240 29404
rect 81176 29344 81240 29348
rect 81256 29404 81320 29408
rect 81256 29348 81260 29404
rect 81260 29348 81316 29404
rect 81316 29348 81320 29404
rect 81256 29344 81320 29348
rect 111736 29404 111800 29408
rect 111736 29348 111740 29404
rect 111740 29348 111796 29404
rect 111796 29348 111800 29404
rect 111736 29344 111800 29348
rect 111816 29404 111880 29408
rect 111816 29348 111820 29404
rect 111820 29348 111876 29404
rect 111876 29348 111880 29404
rect 111816 29344 111880 29348
rect 111896 29404 111960 29408
rect 111896 29348 111900 29404
rect 111900 29348 111956 29404
rect 111956 29348 111960 29404
rect 111896 29344 111960 29348
rect 111976 29404 112040 29408
rect 111976 29348 111980 29404
rect 111980 29348 112036 29404
rect 112036 29348 112040 29404
rect 111976 29344 112040 29348
rect 142456 29404 142520 29408
rect 142456 29348 142460 29404
rect 142460 29348 142516 29404
rect 142516 29348 142520 29404
rect 142456 29344 142520 29348
rect 142536 29404 142600 29408
rect 142536 29348 142540 29404
rect 142540 29348 142596 29404
rect 142596 29348 142600 29404
rect 142536 29344 142600 29348
rect 142616 29404 142680 29408
rect 142616 29348 142620 29404
rect 142620 29348 142676 29404
rect 142676 29348 142680 29404
rect 142616 29344 142680 29348
rect 142696 29404 142760 29408
rect 142696 29348 142700 29404
rect 142700 29348 142756 29404
rect 142756 29348 142760 29404
rect 142696 29344 142760 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 65656 28860 65720 28864
rect 65656 28804 65660 28860
rect 65660 28804 65716 28860
rect 65716 28804 65720 28860
rect 65656 28800 65720 28804
rect 65736 28860 65800 28864
rect 65736 28804 65740 28860
rect 65740 28804 65796 28860
rect 65796 28804 65800 28860
rect 65736 28800 65800 28804
rect 65816 28860 65880 28864
rect 65816 28804 65820 28860
rect 65820 28804 65876 28860
rect 65876 28804 65880 28860
rect 65816 28800 65880 28804
rect 65896 28860 65960 28864
rect 65896 28804 65900 28860
rect 65900 28804 65956 28860
rect 65956 28804 65960 28860
rect 65896 28800 65960 28804
rect 96376 28860 96440 28864
rect 96376 28804 96380 28860
rect 96380 28804 96436 28860
rect 96436 28804 96440 28860
rect 96376 28800 96440 28804
rect 96456 28860 96520 28864
rect 96456 28804 96460 28860
rect 96460 28804 96516 28860
rect 96516 28804 96520 28860
rect 96456 28800 96520 28804
rect 96536 28860 96600 28864
rect 96536 28804 96540 28860
rect 96540 28804 96596 28860
rect 96596 28804 96600 28860
rect 96536 28800 96600 28804
rect 96616 28860 96680 28864
rect 96616 28804 96620 28860
rect 96620 28804 96676 28860
rect 96676 28804 96680 28860
rect 96616 28800 96680 28804
rect 127096 28860 127160 28864
rect 127096 28804 127100 28860
rect 127100 28804 127156 28860
rect 127156 28804 127160 28860
rect 127096 28800 127160 28804
rect 127176 28860 127240 28864
rect 127176 28804 127180 28860
rect 127180 28804 127236 28860
rect 127236 28804 127240 28860
rect 127176 28800 127240 28804
rect 127256 28860 127320 28864
rect 127256 28804 127260 28860
rect 127260 28804 127316 28860
rect 127316 28804 127320 28860
rect 127256 28800 127320 28804
rect 127336 28860 127400 28864
rect 127336 28804 127340 28860
rect 127340 28804 127396 28860
rect 127396 28804 127400 28860
rect 127336 28800 127400 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 81016 28316 81080 28320
rect 81016 28260 81020 28316
rect 81020 28260 81076 28316
rect 81076 28260 81080 28316
rect 81016 28256 81080 28260
rect 81096 28316 81160 28320
rect 81096 28260 81100 28316
rect 81100 28260 81156 28316
rect 81156 28260 81160 28316
rect 81096 28256 81160 28260
rect 81176 28316 81240 28320
rect 81176 28260 81180 28316
rect 81180 28260 81236 28316
rect 81236 28260 81240 28316
rect 81176 28256 81240 28260
rect 81256 28316 81320 28320
rect 81256 28260 81260 28316
rect 81260 28260 81316 28316
rect 81316 28260 81320 28316
rect 81256 28256 81320 28260
rect 111736 28316 111800 28320
rect 111736 28260 111740 28316
rect 111740 28260 111796 28316
rect 111796 28260 111800 28316
rect 111736 28256 111800 28260
rect 111816 28316 111880 28320
rect 111816 28260 111820 28316
rect 111820 28260 111876 28316
rect 111876 28260 111880 28316
rect 111816 28256 111880 28260
rect 111896 28316 111960 28320
rect 111896 28260 111900 28316
rect 111900 28260 111956 28316
rect 111956 28260 111960 28316
rect 111896 28256 111960 28260
rect 111976 28316 112040 28320
rect 111976 28260 111980 28316
rect 111980 28260 112036 28316
rect 112036 28260 112040 28316
rect 111976 28256 112040 28260
rect 142456 28316 142520 28320
rect 142456 28260 142460 28316
rect 142460 28260 142516 28316
rect 142516 28260 142520 28316
rect 142456 28256 142520 28260
rect 142536 28316 142600 28320
rect 142536 28260 142540 28316
rect 142540 28260 142596 28316
rect 142596 28260 142600 28316
rect 142536 28256 142600 28260
rect 142616 28316 142680 28320
rect 142616 28260 142620 28316
rect 142620 28260 142676 28316
rect 142676 28260 142680 28316
rect 142616 28256 142680 28260
rect 142696 28316 142760 28320
rect 142696 28260 142700 28316
rect 142700 28260 142756 28316
rect 142756 28260 142760 28316
rect 142696 28256 142760 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 65656 27772 65720 27776
rect 65656 27716 65660 27772
rect 65660 27716 65716 27772
rect 65716 27716 65720 27772
rect 65656 27712 65720 27716
rect 65736 27772 65800 27776
rect 65736 27716 65740 27772
rect 65740 27716 65796 27772
rect 65796 27716 65800 27772
rect 65736 27712 65800 27716
rect 65816 27772 65880 27776
rect 65816 27716 65820 27772
rect 65820 27716 65876 27772
rect 65876 27716 65880 27772
rect 65816 27712 65880 27716
rect 65896 27772 65960 27776
rect 65896 27716 65900 27772
rect 65900 27716 65956 27772
rect 65956 27716 65960 27772
rect 65896 27712 65960 27716
rect 96376 27772 96440 27776
rect 96376 27716 96380 27772
rect 96380 27716 96436 27772
rect 96436 27716 96440 27772
rect 96376 27712 96440 27716
rect 96456 27772 96520 27776
rect 96456 27716 96460 27772
rect 96460 27716 96516 27772
rect 96516 27716 96520 27772
rect 96456 27712 96520 27716
rect 96536 27772 96600 27776
rect 96536 27716 96540 27772
rect 96540 27716 96596 27772
rect 96596 27716 96600 27772
rect 96536 27712 96600 27716
rect 96616 27772 96680 27776
rect 96616 27716 96620 27772
rect 96620 27716 96676 27772
rect 96676 27716 96680 27772
rect 96616 27712 96680 27716
rect 127096 27772 127160 27776
rect 127096 27716 127100 27772
rect 127100 27716 127156 27772
rect 127156 27716 127160 27772
rect 127096 27712 127160 27716
rect 127176 27772 127240 27776
rect 127176 27716 127180 27772
rect 127180 27716 127236 27772
rect 127236 27716 127240 27772
rect 127176 27712 127240 27716
rect 127256 27772 127320 27776
rect 127256 27716 127260 27772
rect 127260 27716 127316 27772
rect 127316 27716 127320 27772
rect 127256 27712 127320 27716
rect 127336 27772 127400 27776
rect 127336 27716 127340 27772
rect 127340 27716 127396 27772
rect 127396 27716 127400 27772
rect 127336 27712 127400 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 81016 27228 81080 27232
rect 81016 27172 81020 27228
rect 81020 27172 81076 27228
rect 81076 27172 81080 27228
rect 81016 27168 81080 27172
rect 81096 27228 81160 27232
rect 81096 27172 81100 27228
rect 81100 27172 81156 27228
rect 81156 27172 81160 27228
rect 81096 27168 81160 27172
rect 81176 27228 81240 27232
rect 81176 27172 81180 27228
rect 81180 27172 81236 27228
rect 81236 27172 81240 27228
rect 81176 27168 81240 27172
rect 81256 27228 81320 27232
rect 81256 27172 81260 27228
rect 81260 27172 81316 27228
rect 81316 27172 81320 27228
rect 81256 27168 81320 27172
rect 111736 27228 111800 27232
rect 111736 27172 111740 27228
rect 111740 27172 111796 27228
rect 111796 27172 111800 27228
rect 111736 27168 111800 27172
rect 111816 27228 111880 27232
rect 111816 27172 111820 27228
rect 111820 27172 111876 27228
rect 111876 27172 111880 27228
rect 111816 27168 111880 27172
rect 111896 27228 111960 27232
rect 111896 27172 111900 27228
rect 111900 27172 111956 27228
rect 111956 27172 111960 27228
rect 111896 27168 111960 27172
rect 111976 27228 112040 27232
rect 111976 27172 111980 27228
rect 111980 27172 112036 27228
rect 112036 27172 112040 27228
rect 111976 27168 112040 27172
rect 142456 27228 142520 27232
rect 142456 27172 142460 27228
rect 142460 27172 142516 27228
rect 142516 27172 142520 27228
rect 142456 27168 142520 27172
rect 142536 27228 142600 27232
rect 142536 27172 142540 27228
rect 142540 27172 142596 27228
rect 142596 27172 142600 27228
rect 142536 27168 142600 27172
rect 142616 27228 142680 27232
rect 142616 27172 142620 27228
rect 142620 27172 142676 27228
rect 142676 27172 142680 27228
rect 142616 27168 142680 27172
rect 142696 27228 142760 27232
rect 142696 27172 142700 27228
rect 142700 27172 142756 27228
rect 142756 27172 142760 27228
rect 142696 27168 142760 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 65656 26684 65720 26688
rect 65656 26628 65660 26684
rect 65660 26628 65716 26684
rect 65716 26628 65720 26684
rect 65656 26624 65720 26628
rect 65736 26684 65800 26688
rect 65736 26628 65740 26684
rect 65740 26628 65796 26684
rect 65796 26628 65800 26684
rect 65736 26624 65800 26628
rect 65816 26684 65880 26688
rect 65816 26628 65820 26684
rect 65820 26628 65876 26684
rect 65876 26628 65880 26684
rect 65816 26624 65880 26628
rect 65896 26684 65960 26688
rect 65896 26628 65900 26684
rect 65900 26628 65956 26684
rect 65956 26628 65960 26684
rect 65896 26624 65960 26628
rect 96376 26684 96440 26688
rect 96376 26628 96380 26684
rect 96380 26628 96436 26684
rect 96436 26628 96440 26684
rect 96376 26624 96440 26628
rect 96456 26684 96520 26688
rect 96456 26628 96460 26684
rect 96460 26628 96516 26684
rect 96516 26628 96520 26684
rect 96456 26624 96520 26628
rect 96536 26684 96600 26688
rect 96536 26628 96540 26684
rect 96540 26628 96596 26684
rect 96596 26628 96600 26684
rect 96536 26624 96600 26628
rect 96616 26684 96680 26688
rect 96616 26628 96620 26684
rect 96620 26628 96676 26684
rect 96676 26628 96680 26684
rect 96616 26624 96680 26628
rect 127096 26684 127160 26688
rect 127096 26628 127100 26684
rect 127100 26628 127156 26684
rect 127156 26628 127160 26684
rect 127096 26624 127160 26628
rect 127176 26684 127240 26688
rect 127176 26628 127180 26684
rect 127180 26628 127236 26684
rect 127236 26628 127240 26684
rect 127176 26624 127240 26628
rect 127256 26684 127320 26688
rect 127256 26628 127260 26684
rect 127260 26628 127316 26684
rect 127316 26628 127320 26684
rect 127256 26624 127320 26628
rect 127336 26684 127400 26688
rect 127336 26628 127340 26684
rect 127340 26628 127396 26684
rect 127396 26628 127400 26684
rect 127336 26624 127400 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 81016 26140 81080 26144
rect 81016 26084 81020 26140
rect 81020 26084 81076 26140
rect 81076 26084 81080 26140
rect 81016 26080 81080 26084
rect 81096 26140 81160 26144
rect 81096 26084 81100 26140
rect 81100 26084 81156 26140
rect 81156 26084 81160 26140
rect 81096 26080 81160 26084
rect 81176 26140 81240 26144
rect 81176 26084 81180 26140
rect 81180 26084 81236 26140
rect 81236 26084 81240 26140
rect 81176 26080 81240 26084
rect 81256 26140 81320 26144
rect 81256 26084 81260 26140
rect 81260 26084 81316 26140
rect 81316 26084 81320 26140
rect 81256 26080 81320 26084
rect 111736 26140 111800 26144
rect 111736 26084 111740 26140
rect 111740 26084 111796 26140
rect 111796 26084 111800 26140
rect 111736 26080 111800 26084
rect 111816 26140 111880 26144
rect 111816 26084 111820 26140
rect 111820 26084 111876 26140
rect 111876 26084 111880 26140
rect 111816 26080 111880 26084
rect 111896 26140 111960 26144
rect 111896 26084 111900 26140
rect 111900 26084 111956 26140
rect 111956 26084 111960 26140
rect 111896 26080 111960 26084
rect 111976 26140 112040 26144
rect 111976 26084 111980 26140
rect 111980 26084 112036 26140
rect 112036 26084 112040 26140
rect 111976 26080 112040 26084
rect 142456 26140 142520 26144
rect 142456 26084 142460 26140
rect 142460 26084 142516 26140
rect 142516 26084 142520 26140
rect 142456 26080 142520 26084
rect 142536 26140 142600 26144
rect 142536 26084 142540 26140
rect 142540 26084 142596 26140
rect 142596 26084 142600 26140
rect 142536 26080 142600 26084
rect 142616 26140 142680 26144
rect 142616 26084 142620 26140
rect 142620 26084 142676 26140
rect 142676 26084 142680 26140
rect 142616 26080 142680 26084
rect 142696 26140 142760 26144
rect 142696 26084 142700 26140
rect 142700 26084 142756 26140
rect 142756 26084 142760 26140
rect 142696 26080 142760 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 65656 25596 65720 25600
rect 65656 25540 65660 25596
rect 65660 25540 65716 25596
rect 65716 25540 65720 25596
rect 65656 25536 65720 25540
rect 65736 25596 65800 25600
rect 65736 25540 65740 25596
rect 65740 25540 65796 25596
rect 65796 25540 65800 25596
rect 65736 25536 65800 25540
rect 65816 25596 65880 25600
rect 65816 25540 65820 25596
rect 65820 25540 65876 25596
rect 65876 25540 65880 25596
rect 65816 25536 65880 25540
rect 65896 25596 65960 25600
rect 65896 25540 65900 25596
rect 65900 25540 65956 25596
rect 65956 25540 65960 25596
rect 65896 25536 65960 25540
rect 96376 25596 96440 25600
rect 96376 25540 96380 25596
rect 96380 25540 96436 25596
rect 96436 25540 96440 25596
rect 96376 25536 96440 25540
rect 96456 25596 96520 25600
rect 96456 25540 96460 25596
rect 96460 25540 96516 25596
rect 96516 25540 96520 25596
rect 96456 25536 96520 25540
rect 96536 25596 96600 25600
rect 96536 25540 96540 25596
rect 96540 25540 96596 25596
rect 96596 25540 96600 25596
rect 96536 25536 96600 25540
rect 96616 25596 96680 25600
rect 96616 25540 96620 25596
rect 96620 25540 96676 25596
rect 96676 25540 96680 25596
rect 96616 25536 96680 25540
rect 127096 25596 127160 25600
rect 127096 25540 127100 25596
rect 127100 25540 127156 25596
rect 127156 25540 127160 25596
rect 127096 25536 127160 25540
rect 127176 25596 127240 25600
rect 127176 25540 127180 25596
rect 127180 25540 127236 25596
rect 127236 25540 127240 25596
rect 127176 25536 127240 25540
rect 127256 25596 127320 25600
rect 127256 25540 127260 25596
rect 127260 25540 127316 25596
rect 127316 25540 127320 25596
rect 127256 25536 127320 25540
rect 127336 25596 127400 25600
rect 127336 25540 127340 25596
rect 127340 25540 127396 25596
rect 127396 25540 127400 25596
rect 127336 25536 127400 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 81016 25052 81080 25056
rect 81016 24996 81020 25052
rect 81020 24996 81076 25052
rect 81076 24996 81080 25052
rect 81016 24992 81080 24996
rect 81096 25052 81160 25056
rect 81096 24996 81100 25052
rect 81100 24996 81156 25052
rect 81156 24996 81160 25052
rect 81096 24992 81160 24996
rect 81176 25052 81240 25056
rect 81176 24996 81180 25052
rect 81180 24996 81236 25052
rect 81236 24996 81240 25052
rect 81176 24992 81240 24996
rect 81256 25052 81320 25056
rect 81256 24996 81260 25052
rect 81260 24996 81316 25052
rect 81316 24996 81320 25052
rect 81256 24992 81320 24996
rect 111736 25052 111800 25056
rect 111736 24996 111740 25052
rect 111740 24996 111796 25052
rect 111796 24996 111800 25052
rect 111736 24992 111800 24996
rect 111816 25052 111880 25056
rect 111816 24996 111820 25052
rect 111820 24996 111876 25052
rect 111876 24996 111880 25052
rect 111816 24992 111880 24996
rect 111896 25052 111960 25056
rect 111896 24996 111900 25052
rect 111900 24996 111956 25052
rect 111956 24996 111960 25052
rect 111896 24992 111960 24996
rect 111976 25052 112040 25056
rect 111976 24996 111980 25052
rect 111980 24996 112036 25052
rect 112036 24996 112040 25052
rect 111976 24992 112040 24996
rect 142456 25052 142520 25056
rect 142456 24996 142460 25052
rect 142460 24996 142516 25052
rect 142516 24996 142520 25052
rect 142456 24992 142520 24996
rect 142536 25052 142600 25056
rect 142536 24996 142540 25052
rect 142540 24996 142596 25052
rect 142596 24996 142600 25052
rect 142536 24992 142600 24996
rect 142616 25052 142680 25056
rect 142616 24996 142620 25052
rect 142620 24996 142676 25052
rect 142676 24996 142680 25052
rect 142616 24992 142680 24996
rect 142696 25052 142760 25056
rect 142696 24996 142700 25052
rect 142700 24996 142756 25052
rect 142756 24996 142760 25052
rect 142696 24992 142760 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 65656 24508 65720 24512
rect 65656 24452 65660 24508
rect 65660 24452 65716 24508
rect 65716 24452 65720 24508
rect 65656 24448 65720 24452
rect 65736 24508 65800 24512
rect 65736 24452 65740 24508
rect 65740 24452 65796 24508
rect 65796 24452 65800 24508
rect 65736 24448 65800 24452
rect 65816 24508 65880 24512
rect 65816 24452 65820 24508
rect 65820 24452 65876 24508
rect 65876 24452 65880 24508
rect 65816 24448 65880 24452
rect 65896 24508 65960 24512
rect 65896 24452 65900 24508
rect 65900 24452 65956 24508
rect 65956 24452 65960 24508
rect 65896 24448 65960 24452
rect 96376 24508 96440 24512
rect 96376 24452 96380 24508
rect 96380 24452 96436 24508
rect 96436 24452 96440 24508
rect 96376 24448 96440 24452
rect 96456 24508 96520 24512
rect 96456 24452 96460 24508
rect 96460 24452 96516 24508
rect 96516 24452 96520 24508
rect 96456 24448 96520 24452
rect 96536 24508 96600 24512
rect 96536 24452 96540 24508
rect 96540 24452 96596 24508
rect 96596 24452 96600 24508
rect 96536 24448 96600 24452
rect 96616 24508 96680 24512
rect 96616 24452 96620 24508
rect 96620 24452 96676 24508
rect 96676 24452 96680 24508
rect 96616 24448 96680 24452
rect 127096 24508 127160 24512
rect 127096 24452 127100 24508
rect 127100 24452 127156 24508
rect 127156 24452 127160 24508
rect 127096 24448 127160 24452
rect 127176 24508 127240 24512
rect 127176 24452 127180 24508
rect 127180 24452 127236 24508
rect 127236 24452 127240 24508
rect 127176 24448 127240 24452
rect 127256 24508 127320 24512
rect 127256 24452 127260 24508
rect 127260 24452 127316 24508
rect 127316 24452 127320 24508
rect 127256 24448 127320 24452
rect 127336 24508 127400 24512
rect 127336 24452 127340 24508
rect 127340 24452 127396 24508
rect 127396 24452 127400 24508
rect 127336 24448 127400 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 81016 23964 81080 23968
rect 81016 23908 81020 23964
rect 81020 23908 81076 23964
rect 81076 23908 81080 23964
rect 81016 23904 81080 23908
rect 81096 23964 81160 23968
rect 81096 23908 81100 23964
rect 81100 23908 81156 23964
rect 81156 23908 81160 23964
rect 81096 23904 81160 23908
rect 81176 23964 81240 23968
rect 81176 23908 81180 23964
rect 81180 23908 81236 23964
rect 81236 23908 81240 23964
rect 81176 23904 81240 23908
rect 81256 23964 81320 23968
rect 81256 23908 81260 23964
rect 81260 23908 81316 23964
rect 81316 23908 81320 23964
rect 81256 23904 81320 23908
rect 111736 23964 111800 23968
rect 111736 23908 111740 23964
rect 111740 23908 111796 23964
rect 111796 23908 111800 23964
rect 111736 23904 111800 23908
rect 111816 23964 111880 23968
rect 111816 23908 111820 23964
rect 111820 23908 111876 23964
rect 111876 23908 111880 23964
rect 111816 23904 111880 23908
rect 111896 23964 111960 23968
rect 111896 23908 111900 23964
rect 111900 23908 111956 23964
rect 111956 23908 111960 23964
rect 111896 23904 111960 23908
rect 111976 23964 112040 23968
rect 111976 23908 111980 23964
rect 111980 23908 112036 23964
rect 112036 23908 112040 23964
rect 111976 23904 112040 23908
rect 142456 23964 142520 23968
rect 142456 23908 142460 23964
rect 142460 23908 142516 23964
rect 142516 23908 142520 23964
rect 142456 23904 142520 23908
rect 142536 23964 142600 23968
rect 142536 23908 142540 23964
rect 142540 23908 142596 23964
rect 142596 23908 142600 23964
rect 142536 23904 142600 23908
rect 142616 23964 142680 23968
rect 142616 23908 142620 23964
rect 142620 23908 142676 23964
rect 142676 23908 142680 23964
rect 142616 23904 142680 23908
rect 142696 23964 142760 23968
rect 142696 23908 142700 23964
rect 142700 23908 142756 23964
rect 142756 23908 142760 23964
rect 142696 23904 142760 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 65656 23420 65720 23424
rect 65656 23364 65660 23420
rect 65660 23364 65716 23420
rect 65716 23364 65720 23420
rect 65656 23360 65720 23364
rect 65736 23420 65800 23424
rect 65736 23364 65740 23420
rect 65740 23364 65796 23420
rect 65796 23364 65800 23420
rect 65736 23360 65800 23364
rect 65816 23420 65880 23424
rect 65816 23364 65820 23420
rect 65820 23364 65876 23420
rect 65876 23364 65880 23420
rect 65816 23360 65880 23364
rect 65896 23420 65960 23424
rect 65896 23364 65900 23420
rect 65900 23364 65956 23420
rect 65956 23364 65960 23420
rect 65896 23360 65960 23364
rect 96376 23420 96440 23424
rect 96376 23364 96380 23420
rect 96380 23364 96436 23420
rect 96436 23364 96440 23420
rect 96376 23360 96440 23364
rect 96456 23420 96520 23424
rect 96456 23364 96460 23420
rect 96460 23364 96516 23420
rect 96516 23364 96520 23420
rect 96456 23360 96520 23364
rect 96536 23420 96600 23424
rect 96536 23364 96540 23420
rect 96540 23364 96596 23420
rect 96596 23364 96600 23420
rect 96536 23360 96600 23364
rect 96616 23420 96680 23424
rect 96616 23364 96620 23420
rect 96620 23364 96676 23420
rect 96676 23364 96680 23420
rect 96616 23360 96680 23364
rect 127096 23420 127160 23424
rect 127096 23364 127100 23420
rect 127100 23364 127156 23420
rect 127156 23364 127160 23420
rect 127096 23360 127160 23364
rect 127176 23420 127240 23424
rect 127176 23364 127180 23420
rect 127180 23364 127236 23420
rect 127236 23364 127240 23420
rect 127176 23360 127240 23364
rect 127256 23420 127320 23424
rect 127256 23364 127260 23420
rect 127260 23364 127316 23420
rect 127316 23364 127320 23420
rect 127256 23360 127320 23364
rect 127336 23420 127400 23424
rect 127336 23364 127340 23420
rect 127340 23364 127396 23420
rect 127396 23364 127400 23420
rect 127336 23360 127400 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 81016 22876 81080 22880
rect 81016 22820 81020 22876
rect 81020 22820 81076 22876
rect 81076 22820 81080 22876
rect 81016 22816 81080 22820
rect 81096 22876 81160 22880
rect 81096 22820 81100 22876
rect 81100 22820 81156 22876
rect 81156 22820 81160 22876
rect 81096 22816 81160 22820
rect 81176 22876 81240 22880
rect 81176 22820 81180 22876
rect 81180 22820 81236 22876
rect 81236 22820 81240 22876
rect 81176 22816 81240 22820
rect 81256 22876 81320 22880
rect 81256 22820 81260 22876
rect 81260 22820 81316 22876
rect 81316 22820 81320 22876
rect 81256 22816 81320 22820
rect 111736 22876 111800 22880
rect 111736 22820 111740 22876
rect 111740 22820 111796 22876
rect 111796 22820 111800 22876
rect 111736 22816 111800 22820
rect 111816 22876 111880 22880
rect 111816 22820 111820 22876
rect 111820 22820 111876 22876
rect 111876 22820 111880 22876
rect 111816 22816 111880 22820
rect 111896 22876 111960 22880
rect 111896 22820 111900 22876
rect 111900 22820 111956 22876
rect 111956 22820 111960 22876
rect 111896 22816 111960 22820
rect 111976 22876 112040 22880
rect 111976 22820 111980 22876
rect 111980 22820 112036 22876
rect 112036 22820 112040 22876
rect 111976 22816 112040 22820
rect 142456 22876 142520 22880
rect 142456 22820 142460 22876
rect 142460 22820 142516 22876
rect 142516 22820 142520 22876
rect 142456 22816 142520 22820
rect 142536 22876 142600 22880
rect 142536 22820 142540 22876
rect 142540 22820 142596 22876
rect 142596 22820 142600 22876
rect 142536 22816 142600 22820
rect 142616 22876 142680 22880
rect 142616 22820 142620 22876
rect 142620 22820 142676 22876
rect 142676 22820 142680 22876
rect 142616 22816 142680 22820
rect 142696 22876 142760 22880
rect 142696 22820 142700 22876
rect 142700 22820 142756 22876
rect 142756 22820 142760 22876
rect 142696 22816 142760 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 65656 22332 65720 22336
rect 65656 22276 65660 22332
rect 65660 22276 65716 22332
rect 65716 22276 65720 22332
rect 65656 22272 65720 22276
rect 65736 22332 65800 22336
rect 65736 22276 65740 22332
rect 65740 22276 65796 22332
rect 65796 22276 65800 22332
rect 65736 22272 65800 22276
rect 65816 22332 65880 22336
rect 65816 22276 65820 22332
rect 65820 22276 65876 22332
rect 65876 22276 65880 22332
rect 65816 22272 65880 22276
rect 65896 22332 65960 22336
rect 65896 22276 65900 22332
rect 65900 22276 65956 22332
rect 65956 22276 65960 22332
rect 65896 22272 65960 22276
rect 96376 22332 96440 22336
rect 96376 22276 96380 22332
rect 96380 22276 96436 22332
rect 96436 22276 96440 22332
rect 96376 22272 96440 22276
rect 96456 22332 96520 22336
rect 96456 22276 96460 22332
rect 96460 22276 96516 22332
rect 96516 22276 96520 22332
rect 96456 22272 96520 22276
rect 96536 22332 96600 22336
rect 96536 22276 96540 22332
rect 96540 22276 96596 22332
rect 96596 22276 96600 22332
rect 96536 22272 96600 22276
rect 96616 22332 96680 22336
rect 96616 22276 96620 22332
rect 96620 22276 96676 22332
rect 96676 22276 96680 22332
rect 96616 22272 96680 22276
rect 127096 22332 127160 22336
rect 127096 22276 127100 22332
rect 127100 22276 127156 22332
rect 127156 22276 127160 22332
rect 127096 22272 127160 22276
rect 127176 22332 127240 22336
rect 127176 22276 127180 22332
rect 127180 22276 127236 22332
rect 127236 22276 127240 22332
rect 127176 22272 127240 22276
rect 127256 22332 127320 22336
rect 127256 22276 127260 22332
rect 127260 22276 127316 22332
rect 127316 22276 127320 22332
rect 127256 22272 127320 22276
rect 127336 22332 127400 22336
rect 127336 22276 127340 22332
rect 127340 22276 127396 22332
rect 127396 22276 127400 22332
rect 127336 22272 127400 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 81016 21788 81080 21792
rect 81016 21732 81020 21788
rect 81020 21732 81076 21788
rect 81076 21732 81080 21788
rect 81016 21728 81080 21732
rect 81096 21788 81160 21792
rect 81096 21732 81100 21788
rect 81100 21732 81156 21788
rect 81156 21732 81160 21788
rect 81096 21728 81160 21732
rect 81176 21788 81240 21792
rect 81176 21732 81180 21788
rect 81180 21732 81236 21788
rect 81236 21732 81240 21788
rect 81176 21728 81240 21732
rect 81256 21788 81320 21792
rect 81256 21732 81260 21788
rect 81260 21732 81316 21788
rect 81316 21732 81320 21788
rect 81256 21728 81320 21732
rect 111736 21788 111800 21792
rect 111736 21732 111740 21788
rect 111740 21732 111796 21788
rect 111796 21732 111800 21788
rect 111736 21728 111800 21732
rect 111816 21788 111880 21792
rect 111816 21732 111820 21788
rect 111820 21732 111876 21788
rect 111876 21732 111880 21788
rect 111816 21728 111880 21732
rect 111896 21788 111960 21792
rect 111896 21732 111900 21788
rect 111900 21732 111956 21788
rect 111956 21732 111960 21788
rect 111896 21728 111960 21732
rect 111976 21788 112040 21792
rect 111976 21732 111980 21788
rect 111980 21732 112036 21788
rect 112036 21732 112040 21788
rect 111976 21728 112040 21732
rect 142456 21788 142520 21792
rect 142456 21732 142460 21788
rect 142460 21732 142516 21788
rect 142516 21732 142520 21788
rect 142456 21728 142520 21732
rect 142536 21788 142600 21792
rect 142536 21732 142540 21788
rect 142540 21732 142596 21788
rect 142596 21732 142600 21788
rect 142536 21728 142600 21732
rect 142616 21788 142680 21792
rect 142616 21732 142620 21788
rect 142620 21732 142676 21788
rect 142676 21732 142680 21788
rect 142616 21728 142680 21732
rect 142696 21788 142760 21792
rect 142696 21732 142700 21788
rect 142700 21732 142756 21788
rect 142756 21732 142760 21788
rect 142696 21728 142760 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 65656 21244 65720 21248
rect 65656 21188 65660 21244
rect 65660 21188 65716 21244
rect 65716 21188 65720 21244
rect 65656 21184 65720 21188
rect 65736 21244 65800 21248
rect 65736 21188 65740 21244
rect 65740 21188 65796 21244
rect 65796 21188 65800 21244
rect 65736 21184 65800 21188
rect 65816 21244 65880 21248
rect 65816 21188 65820 21244
rect 65820 21188 65876 21244
rect 65876 21188 65880 21244
rect 65816 21184 65880 21188
rect 65896 21244 65960 21248
rect 65896 21188 65900 21244
rect 65900 21188 65956 21244
rect 65956 21188 65960 21244
rect 65896 21184 65960 21188
rect 96376 21244 96440 21248
rect 96376 21188 96380 21244
rect 96380 21188 96436 21244
rect 96436 21188 96440 21244
rect 96376 21184 96440 21188
rect 96456 21244 96520 21248
rect 96456 21188 96460 21244
rect 96460 21188 96516 21244
rect 96516 21188 96520 21244
rect 96456 21184 96520 21188
rect 96536 21244 96600 21248
rect 96536 21188 96540 21244
rect 96540 21188 96596 21244
rect 96596 21188 96600 21244
rect 96536 21184 96600 21188
rect 96616 21244 96680 21248
rect 96616 21188 96620 21244
rect 96620 21188 96676 21244
rect 96676 21188 96680 21244
rect 96616 21184 96680 21188
rect 127096 21244 127160 21248
rect 127096 21188 127100 21244
rect 127100 21188 127156 21244
rect 127156 21188 127160 21244
rect 127096 21184 127160 21188
rect 127176 21244 127240 21248
rect 127176 21188 127180 21244
rect 127180 21188 127236 21244
rect 127236 21188 127240 21244
rect 127176 21184 127240 21188
rect 127256 21244 127320 21248
rect 127256 21188 127260 21244
rect 127260 21188 127316 21244
rect 127316 21188 127320 21244
rect 127256 21184 127320 21188
rect 127336 21244 127400 21248
rect 127336 21188 127340 21244
rect 127340 21188 127396 21244
rect 127396 21188 127400 21244
rect 127336 21184 127400 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 81016 20700 81080 20704
rect 81016 20644 81020 20700
rect 81020 20644 81076 20700
rect 81076 20644 81080 20700
rect 81016 20640 81080 20644
rect 81096 20700 81160 20704
rect 81096 20644 81100 20700
rect 81100 20644 81156 20700
rect 81156 20644 81160 20700
rect 81096 20640 81160 20644
rect 81176 20700 81240 20704
rect 81176 20644 81180 20700
rect 81180 20644 81236 20700
rect 81236 20644 81240 20700
rect 81176 20640 81240 20644
rect 81256 20700 81320 20704
rect 81256 20644 81260 20700
rect 81260 20644 81316 20700
rect 81316 20644 81320 20700
rect 81256 20640 81320 20644
rect 111736 20700 111800 20704
rect 111736 20644 111740 20700
rect 111740 20644 111796 20700
rect 111796 20644 111800 20700
rect 111736 20640 111800 20644
rect 111816 20700 111880 20704
rect 111816 20644 111820 20700
rect 111820 20644 111876 20700
rect 111876 20644 111880 20700
rect 111816 20640 111880 20644
rect 111896 20700 111960 20704
rect 111896 20644 111900 20700
rect 111900 20644 111956 20700
rect 111956 20644 111960 20700
rect 111896 20640 111960 20644
rect 111976 20700 112040 20704
rect 111976 20644 111980 20700
rect 111980 20644 112036 20700
rect 112036 20644 112040 20700
rect 111976 20640 112040 20644
rect 142456 20700 142520 20704
rect 142456 20644 142460 20700
rect 142460 20644 142516 20700
rect 142516 20644 142520 20700
rect 142456 20640 142520 20644
rect 142536 20700 142600 20704
rect 142536 20644 142540 20700
rect 142540 20644 142596 20700
rect 142596 20644 142600 20700
rect 142536 20640 142600 20644
rect 142616 20700 142680 20704
rect 142616 20644 142620 20700
rect 142620 20644 142676 20700
rect 142676 20644 142680 20700
rect 142616 20640 142680 20644
rect 142696 20700 142760 20704
rect 142696 20644 142700 20700
rect 142700 20644 142756 20700
rect 142756 20644 142760 20700
rect 142696 20640 142760 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 65656 20156 65720 20160
rect 65656 20100 65660 20156
rect 65660 20100 65716 20156
rect 65716 20100 65720 20156
rect 65656 20096 65720 20100
rect 65736 20156 65800 20160
rect 65736 20100 65740 20156
rect 65740 20100 65796 20156
rect 65796 20100 65800 20156
rect 65736 20096 65800 20100
rect 65816 20156 65880 20160
rect 65816 20100 65820 20156
rect 65820 20100 65876 20156
rect 65876 20100 65880 20156
rect 65816 20096 65880 20100
rect 65896 20156 65960 20160
rect 65896 20100 65900 20156
rect 65900 20100 65956 20156
rect 65956 20100 65960 20156
rect 65896 20096 65960 20100
rect 96376 20156 96440 20160
rect 96376 20100 96380 20156
rect 96380 20100 96436 20156
rect 96436 20100 96440 20156
rect 96376 20096 96440 20100
rect 96456 20156 96520 20160
rect 96456 20100 96460 20156
rect 96460 20100 96516 20156
rect 96516 20100 96520 20156
rect 96456 20096 96520 20100
rect 96536 20156 96600 20160
rect 96536 20100 96540 20156
rect 96540 20100 96596 20156
rect 96596 20100 96600 20156
rect 96536 20096 96600 20100
rect 96616 20156 96680 20160
rect 96616 20100 96620 20156
rect 96620 20100 96676 20156
rect 96676 20100 96680 20156
rect 96616 20096 96680 20100
rect 127096 20156 127160 20160
rect 127096 20100 127100 20156
rect 127100 20100 127156 20156
rect 127156 20100 127160 20156
rect 127096 20096 127160 20100
rect 127176 20156 127240 20160
rect 127176 20100 127180 20156
rect 127180 20100 127236 20156
rect 127236 20100 127240 20156
rect 127176 20096 127240 20100
rect 127256 20156 127320 20160
rect 127256 20100 127260 20156
rect 127260 20100 127316 20156
rect 127316 20100 127320 20156
rect 127256 20096 127320 20100
rect 127336 20156 127400 20160
rect 127336 20100 127340 20156
rect 127340 20100 127396 20156
rect 127396 20100 127400 20156
rect 127336 20096 127400 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 81016 19612 81080 19616
rect 81016 19556 81020 19612
rect 81020 19556 81076 19612
rect 81076 19556 81080 19612
rect 81016 19552 81080 19556
rect 81096 19612 81160 19616
rect 81096 19556 81100 19612
rect 81100 19556 81156 19612
rect 81156 19556 81160 19612
rect 81096 19552 81160 19556
rect 81176 19612 81240 19616
rect 81176 19556 81180 19612
rect 81180 19556 81236 19612
rect 81236 19556 81240 19612
rect 81176 19552 81240 19556
rect 81256 19612 81320 19616
rect 81256 19556 81260 19612
rect 81260 19556 81316 19612
rect 81316 19556 81320 19612
rect 81256 19552 81320 19556
rect 111736 19612 111800 19616
rect 111736 19556 111740 19612
rect 111740 19556 111796 19612
rect 111796 19556 111800 19612
rect 111736 19552 111800 19556
rect 111816 19612 111880 19616
rect 111816 19556 111820 19612
rect 111820 19556 111876 19612
rect 111876 19556 111880 19612
rect 111816 19552 111880 19556
rect 111896 19612 111960 19616
rect 111896 19556 111900 19612
rect 111900 19556 111956 19612
rect 111956 19556 111960 19612
rect 111896 19552 111960 19556
rect 111976 19612 112040 19616
rect 111976 19556 111980 19612
rect 111980 19556 112036 19612
rect 112036 19556 112040 19612
rect 111976 19552 112040 19556
rect 142456 19612 142520 19616
rect 142456 19556 142460 19612
rect 142460 19556 142516 19612
rect 142516 19556 142520 19612
rect 142456 19552 142520 19556
rect 142536 19612 142600 19616
rect 142536 19556 142540 19612
rect 142540 19556 142596 19612
rect 142596 19556 142600 19612
rect 142536 19552 142600 19556
rect 142616 19612 142680 19616
rect 142616 19556 142620 19612
rect 142620 19556 142676 19612
rect 142676 19556 142680 19612
rect 142616 19552 142680 19556
rect 142696 19612 142760 19616
rect 142696 19556 142700 19612
rect 142700 19556 142756 19612
rect 142756 19556 142760 19612
rect 142696 19552 142760 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 65656 19068 65720 19072
rect 65656 19012 65660 19068
rect 65660 19012 65716 19068
rect 65716 19012 65720 19068
rect 65656 19008 65720 19012
rect 65736 19068 65800 19072
rect 65736 19012 65740 19068
rect 65740 19012 65796 19068
rect 65796 19012 65800 19068
rect 65736 19008 65800 19012
rect 65816 19068 65880 19072
rect 65816 19012 65820 19068
rect 65820 19012 65876 19068
rect 65876 19012 65880 19068
rect 65816 19008 65880 19012
rect 65896 19068 65960 19072
rect 65896 19012 65900 19068
rect 65900 19012 65956 19068
rect 65956 19012 65960 19068
rect 65896 19008 65960 19012
rect 96376 19068 96440 19072
rect 96376 19012 96380 19068
rect 96380 19012 96436 19068
rect 96436 19012 96440 19068
rect 96376 19008 96440 19012
rect 96456 19068 96520 19072
rect 96456 19012 96460 19068
rect 96460 19012 96516 19068
rect 96516 19012 96520 19068
rect 96456 19008 96520 19012
rect 96536 19068 96600 19072
rect 96536 19012 96540 19068
rect 96540 19012 96596 19068
rect 96596 19012 96600 19068
rect 96536 19008 96600 19012
rect 96616 19068 96680 19072
rect 96616 19012 96620 19068
rect 96620 19012 96676 19068
rect 96676 19012 96680 19068
rect 96616 19008 96680 19012
rect 127096 19068 127160 19072
rect 127096 19012 127100 19068
rect 127100 19012 127156 19068
rect 127156 19012 127160 19068
rect 127096 19008 127160 19012
rect 127176 19068 127240 19072
rect 127176 19012 127180 19068
rect 127180 19012 127236 19068
rect 127236 19012 127240 19068
rect 127176 19008 127240 19012
rect 127256 19068 127320 19072
rect 127256 19012 127260 19068
rect 127260 19012 127316 19068
rect 127316 19012 127320 19068
rect 127256 19008 127320 19012
rect 127336 19068 127400 19072
rect 127336 19012 127340 19068
rect 127340 19012 127396 19068
rect 127396 19012 127400 19068
rect 127336 19008 127400 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 81016 18524 81080 18528
rect 81016 18468 81020 18524
rect 81020 18468 81076 18524
rect 81076 18468 81080 18524
rect 81016 18464 81080 18468
rect 81096 18524 81160 18528
rect 81096 18468 81100 18524
rect 81100 18468 81156 18524
rect 81156 18468 81160 18524
rect 81096 18464 81160 18468
rect 81176 18524 81240 18528
rect 81176 18468 81180 18524
rect 81180 18468 81236 18524
rect 81236 18468 81240 18524
rect 81176 18464 81240 18468
rect 81256 18524 81320 18528
rect 81256 18468 81260 18524
rect 81260 18468 81316 18524
rect 81316 18468 81320 18524
rect 81256 18464 81320 18468
rect 111736 18524 111800 18528
rect 111736 18468 111740 18524
rect 111740 18468 111796 18524
rect 111796 18468 111800 18524
rect 111736 18464 111800 18468
rect 111816 18524 111880 18528
rect 111816 18468 111820 18524
rect 111820 18468 111876 18524
rect 111876 18468 111880 18524
rect 111816 18464 111880 18468
rect 111896 18524 111960 18528
rect 111896 18468 111900 18524
rect 111900 18468 111956 18524
rect 111956 18468 111960 18524
rect 111896 18464 111960 18468
rect 111976 18524 112040 18528
rect 111976 18468 111980 18524
rect 111980 18468 112036 18524
rect 112036 18468 112040 18524
rect 111976 18464 112040 18468
rect 142456 18524 142520 18528
rect 142456 18468 142460 18524
rect 142460 18468 142516 18524
rect 142516 18468 142520 18524
rect 142456 18464 142520 18468
rect 142536 18524 142600 18528
rect 142536 18468 142540 18524
rect 142540 18468 142596 18524
rect 142596 18468 142600 18524
rect 142536 18464 142600 18468
rect 142616 18524 142680 18528
rect 142616 18468 142620 18524
rect 142620 18468 142676 18524
rect 142676 18468 142680 18524
rect 142616 18464 142680 18468
rect 142696 18524 142760 18528
rect 142696 18468 142700 18524
rect 142700 18468 142756 18524
rect 142756 18468 142760 18524
rect 142696 18464 142760 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 65656 17980 65720 17984
rect 65656 17924 65660 17980
rect 65660 17924 65716 17980
rect 65716 17924 65720 17980
rect 65656 17920 65720 17924
rect 65736 17980 65800 17984
rect 65736 17924 65740 17980
rect 65740 17924 65796 17980
rect 65796 17924 65800 17980
rect 65736 17920 65800 17924
rect 65816 17980 65880 17984
rect 65816 17924 65820 17980
rect 65820 17924 65876 17980
rect 65876 17924 65880 17980
rect 65816 17920 65880 17924
rect 65896 17980 65960 17984
rect 65896 17924 65900 17980
rect 65900 17924 65956 17980
rect 65956 17924 65960 17980
rect 65896 17920 65960 17924
rect 96376 17980 96440 17984
rect 96376 17924 96380 17980
rect 96380 17924 96436 17980
rect 96436 17924 96440 17980
rect 96376 17920 96440 17924
rect 96456 17980 96520 17984
rect 96456 17924 96460 17980
rect 96460 17924 96516 17980
rect 96516 17924 96520 17980
rect 96456 17920 96520 17924
rect 96536 17980 96600 17984
rect 96536 17924 96540 17980
rect 96540 17924 96596 17980
rect 96596 17924 96600 17980
rect 96536 17920 96600 17924
rect 96616 17980 96680 17984
rect 96616 17924 96620 17980
rect 96620 17924 96676 17980
rect 96676 17924 96680 17980
rect 96616 17920 96680 17924
rect 127096 17980 127160 17984
rect 127096 17924 127100 17980
rect 127100 17924 127156 17980
rect 127156 17924 127160 17980
rect 127096 17920 127160 17924
rect 127176 17980 127240 17984
rect 127176 17924 127180 17980
rect 127180 17924 127236 17980
rect 127236 17924 127240 17980
rect 127176 17920 127240 17924
rect 127256 17980 127320 17984
rect 127256 17924 127260 17980
rect 127260 17924 127316 17980
rect 127316 17924 127320 17980
rect 127256 17920 127320 17924
rect 127336 17980 127400 17984
rect 127336 17924 127340 17980
rect 127340 17924 127396 17980
rect 127396 17924 127400 17980
rect 127336 17920 127400 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 81016 17436 81080 17440
rect 81016 17380 81020 17436
rect 81020 17380 81076 17436
rect 81076 17380 81080 17436
rect 81016 17376 81080 17380
rect 81096 17436 81160 17440
rect 81096 17380 81100 17436
rect 81100 17380 81156 17436
rect 81156 17380 81160 17436
rect 81096 17376 81160 17380
rect 81176 17436 81240 17440
rect 81176 17380 81180 17436
rect 81180 17380 81236 17436
rect 81236 17380 81240 17436
rect 81176 17376 81240 17380
rect 81256 17436 81320 17440
rect 81256 17380 81260 17436
rect 81260 17380 81316 17436
rect 81316 17380 81320 17436
rect 81256 17376 81320 17380
rect 111736 17436 111800 17440
rect 111736 17380 111740 17436
rect 111740 17380 111796 17436
rect 111796 17380 111800 17436
rect 111736 17376 111800 17380
rect 111816 17436 111880 17440
rect 111816 17380 111820 17436
rect 111820 17380 111876 17436
rect 111876 17380 111880 17436
rect 111816 17376 111880 17380
rect 111896 17436 111960 17440
rect 111896 17380 111900 17436
rect 111900 17380 111956 17436
rect 111956 17380 111960 17436
rect 111896 17376 111960 17380
rect 111976 17436 112040 17440
rect 111976 17380 111980 17436
rect 111980 17380 112036 17436
rect 112036 17380 112040 17436
rect 111976 17376 112040 17380
rect 142456 17436 142520 17440
rect 142456 17380 142460 17436
rect 142460 17380 142516 17436
rect 142516 17380 142520 17436
rect 142456 17376 142520 17380
rect 142536 17436 142600 17440
rect 142536 17380 142540 17436
rect 142540 17380 142596 17436
rect 142596 17380 142600 17436
rect 142536 17376 142600 17380
rect 142616 17436 142680 17440
rect 142616 17380 142620 17436
rect 142620 17380 142676 17436
rect 142676 17380 142680 17436
rect 142616 17376 142680 17380
rect 142696 17436 142760 17440
rect 142696 17380 142700 17436
rect 142700 17380 142756 17436
rect 142756 17380 142760 17436
rect 142696 17376 142760 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 65656 16892 65720 16896
rect 65656 16836 65660 16892
rect 65660 16836 65716 16892
rect 65716 16836 65720 16892
rect 65656 16832 65720 16836
rect 65736 16892 65800 16896
rect 65736 16836 65740 16892
rect 65740 16836 65796 16892
rect 65796 16836 65800 16892
rect 65736 16832 65800 16836
rect 65816 16892 65880 16896
rect 65816 16836 65820 16892
rect 65820 16836 65876 16892
rect 65876 16836 65880 16892
rect 65816 16832 65880 16836
rect 65896 16892 65960 16896
rect 65896 16836 65900 16892
rect 65900 16836 65956 16892
rect 65956 16836 65960 16892
rect 65896 16832 65960 16836
rect 96376 16892 96440 16896
rect 96376 16836 96380 16892
rect 96380 16836 96436 16892
rect 96436 16836 96440 16892
rect 96376 16832 96440 16836
rect 96456 16892 96520 16896
rect 96456 16836 96460 16892
rect 96460 16836 96516 16892
rect 96516 16836 96520 16892
rect 96456 16832 96520 16836
rect 96536 16892 96600 16896
rect 96536 16836 96540 16892
rect 96540 16836 96596 16892
rect 96596 16836 96600 16892
rect 96536 16832 96600 16836
rect 96616 16892 96680 16896
rect 96616 16836 96620 16892
rect 96620 16836 96676 16892
rect 96676 16836 96680 16892
rect 96616 16832 96680 16836
rect 127096 16892 127160 16896
rect 127096 16836 127100 16892
rect 127100 16836 127156 16892
rect 127156 16836 127160 16892
rect 127096 16832 127160 16836
rect 127176 16892 127240 16896
rect 127176 16836 127180 16892
rect 127180 16836 127236 16892
rect 127236 16836 127240 16892
rect 127176 16832 127240 16836
rect 127256 16892 127320 16896
rect 127256 16836 127260 16892
rect 127260 16836 127316 16892
rect 127316 16836 127320 16892
rect 127256 16832 127320 16836
rect 127336 16892 127400 16896
rect 127336 16836 127340 16892
rect 127340 16836 127396 16892
rect 127396 16836 127400 16892
rect 127336 16832 127400 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 81016 16348 81080 16352
rect 81016 16292 81020 16348
rect 81020 16292 81076 16348
rect 81076 16292 81080 16348
rect 81016 16288 81080 16292
rect 81096 16348 81160 16352
rect 81096 16292 81100 16348
rect 81100 16292 81156 16348
rect 81156 16292 81160 16348
rect 81096 16288 81160 16292
rect 81176 16348 81240 16352
rect 81176 16292 81180 16348
rect 81180 16292 81236 16348
rect 81236 16292 81240 16348
rect 81176 16288 81240 16292
rect 81256 16348 81320 16352
rect 81256 16292 81260 16348
rect 81260 16292 81316 16348
rect 81316 16292 81320 16348
rect 81256 16288 81320 16292
rect 111736 16348 111800 16352
rect 111736 16292 111740 16348
rect 111740 16292 111796 16348
rect 111796 16292 111800 16348
rect 111736 16288 111800 16292
rect 111816 16348 111880 16352
rect 111816 16292 111820 16348
rect 111820 16292 111876 16348
rect 111876 16292 111880 16348
rect 111816 16288 111880 16292
rect 111896 16348 111960 16352
rect 111896 16292 111900 16348
rect 111900 16292 111956 16348
rect 111956 16292 111960 16348
rect 111896 16288 111960 16292
rect 111976 16348 112040 16352
rect 111976 16292 111980 16348
rect 111980 16292 112036 16348
rect 112036 16292 112040 16348
rect 111976 16288 112040 16292
rect 142456 16348 142520 16352
rect 142456 16292 142460 16348
rect 142460 16292 142516 16348
rect 142516 16292 142520 16348
rect 142456 16288 142520 16292
rect 142536 16348 142600 16352
rect 142536 16292 142540 16348
rect 142540 16292 142596 16348
rect 142596 16292 142600 16348
rect 142536 16288 142600 16292
rect 142616 16348 142680 16352
rect 142616 16292 142620 16348
rect 142620 16292 142676 16348
rect 142676 16292 142680 16348
rect 142616 16288 142680 16292
rect 142696 16348 142760 16352
rect 142696 16292 142700 16348
rect 142700 16292 142756 16348
rect 142756 16292 142760 16348
rect 142696 16288 142760 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 65656 15804 65720 15808
rect 65656 15748 65660 15804
rect 65660 15748 65716 15804
rect 65716 15748 65720 15804
rect 65656 15744 65720 15748
rect 65736 15804 65800 15808
rect 65736 15748 65740 15804
rect 65740 15748 65796 15804
rect 65796 15748 65800 15804
rect 65736 15744 65800 15748
rect 65816 15804 65880 15808
rect 65816 15748 65820 15804
rect 65820 15748 65876 15804
rect 65876 15748 65880 15804
rect 65816 15744 65880 15748
rect 65896 15804 65960 15808
rect 65896 15748 65900 15804
rect 65900 15748 65956 15804
rect 65956 15748 65960 15804
rect 65896 15744 65960 15748
rect 96376 15804 96440 15808
rect 96376 15748 96380 15804
rect 96380 15748 96436 15804
rect 96436 15748 96440 15804
rect 96376 15744 96440 15748
rect 96456 15804 96520 15808
rect 96456 15748 96460 15804
rect 96460 15748 96516 15804
rect 96516 15748 96520 15804
rect 96456 15744 96520 15748
rect 96536 15804 96600 15808
rect 96536 15748 96540 15804
rect 96540 15748 96596 15804
rect 96596 15748 96600 15804
rect 96536 15744 96600 15748
rect 96616 15804 96680 15808
rect 96616 15748 96620 15804
rect 96620 15748 96676 15804
rect 96676 15748 96680 15804
rect 96616 15744 96680 15748
rect 127096 15804 127160 15808
rect 127096 15748 127100 15804
rect 127100 15748 127156 15804
rect 127156 15748 127160 15804
rect 127096 15744 127160 15748
rect 127176 15804 127240 15808
rect 127176 15748 127180 15804
rect 127180 15748 127236 15804
rect 127236 15748 127240 15804
rect 127176 15744 127240 15748
rect 127256 15804 127320 15808
rect 127256 15748 127260 15804
rect 127260 15748 127316 15804
rect 127316 15748 127320 15804
rect 127256 15744 127320 15748
rect 127336 15804 127400 15808
rect 127336 15748 127340 15804
rect 127340 15748 127396 15804
rect 127396 15748 127400 15804
rect 127336 15744 127400 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 81016 15260 81080 15264
rect 81016 15204 81020 15260
rect 81020 15204 81076 15260
rect 81076 15204 81080 15260
rect 81016 15200 81080 15204
rect 81096 15260 81160 15264
rect 81096 15204 81100 15260
rect 81100 15204 81156 15260
rect 81156 15204 81160 15260
rect 81096 15200 81160 15204
rect 81176 15260 81240 15264
rect 81176 15204 81180 15260
rect 81180 15204 81236 15260
rect 81236 15204 81240 15260
rect 81176 15200 81240 15204
rect 81256 15260 81320 15264
rect 81256 15204 81260 15260
rect 81260 15204 81316 15260
rect 81316 15204 81320 15260
rect 81256 15200 81320 15204
rect 111736 15260 111800 15264
rect 111736 15204 111740 15260
rect 111740 15204 111796 15260
rect 111796 15204 111800 15260
rect 111736 15200 111800 15204
rect 111816 15260 111880 15264
rect 111816 15204 111820 15260
rect 111820 15204 111876 15260
rect 111876 15204 111880 15260
rect 111816 15200 111880 15204
rect 111896 15260 111960 15264
rect 111896 15204 111900 15260
rect 111900 15204 111956 15260
rect 111956 15204 111960 15260
rect 111896 15200 111960 15204
rect 111976 15260 112040 15264
rect 111976 15204 111980 15260
rect 111980 15204 112036 15260
rect 112036 15204 112040 15260
rect 111976 15200 112040 15204
rect 142456 15260 142520 15264
rect 142456 15204 142460 15260
rect 142460 15204 142516 15260
rect 142516 15204 142520 15260
rect 142456 15200 142520 15204
rect 142536 15260 142600 15264
rect 142536 15204 142540 15260
rect 142540 15204 142596 15260
rect 142596 15204 142600 15260
rect 142536 15200 142600 15204
rect 142616 15260 142680 15264
rect 142616 15204 142620 15260
rect 142620 15204 142676 15260
rect 142676 15204 142680 15260
rect 142616 15200 142680 15204
rect 142696 15260 142760 15264
rect 142696 15204 142700 15260
rect 142700 15204 142756 15260
rect 142756 15204 142760 15260
rect 142696 15200 142760 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 65656 14716 65720 14720
rect 65656 14660 65660 14716
rect 65660 14660 65716 14716
rect 65716 14660 65720 14716
rect 65656 14656 65720 14660
rect 65736 14716 65800 14720
rect 65736 14660 65740 14716
rect 65740 14660 65796 14716
rect 65796 14660 65800 14716
rect 65736 14656 65800 14660
rect 65816 14716 65880 14720
rect 65816 14660 65820 14716
rect 65820 14660 65876 14716
rect 65876 14660 65880 14716
rect 65816 14656 65880 14660
rect 65896 14716 65960 14720
rect 65896 14660 65900 14716
rect 65900 14660 65956 14716
rect 65956 14660 65960 14716
rect 65896 14656 65960 14660
rect 96376 14716 96440 14720
rect 96376 14660 96380 14716
rect 96380 14660 96436 14716
rect 96436 14660 96440 14716
rect 96376 14656 96440 14660
rect 96456 14716 96520 14720
rect 96456 14660 96460 14716
rect 96460 14660 96516 14716
rect 96516 14660 96520 14716
rect 96456 14656 96520 14660
rect 96536 14716 96600 14720
rect 96536 14660 96540 14716
rect 96540 14660 96596 14716
rect 96596 14660 96600 14716
rect 96536 14656 96600 14660
rect 96616 14716 96680 14720
rect 96616 14660 96620 14716
rect 96620 14660 96676 14716
rect 96676 14660 96680 14716
rect 96616 14656 96680 14660
rect 127096 14716 127160 14720
rect 127096 14660 127100 14716
rect 127100 14660 127156 14716
rect 127156 14660 127160 14716
rect 127096 14656 127160 14660
rect 127176 14716 127240 14720
rect 127176 14660 127180 14716
rect 127180 14660 127236 14716
rect 127236 14660 127240 14716
rect 127176 14656 127240 14660
rect 127256 14716 127320 14720
rect 127256 14660 127260 14716
rect 127260 14660 127316 14716
rect 127316 14660 127320 14716
rect 127256 14656 127320 14660
rect 127336 14716 127400 14720
rect 127336 14660 127340 14716
rect 127340 14660 127396 14716
rect 127396 14660 127400 14716
rect 127336 14656 127400 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 81016 14172 81080 14176
rect 81016 14116 81020 14172
rect 81020 14116 81076 14172
rect 81076 14116 81080 14172
rect 81016 14112 81080 14116
rect 81096 14172 81160 14176
rect 81096 14116 81100 14172
rect 81100 14116 81156 14172
rect 81156 14116 81160 14172
rect 81096 14112 81160 14116
rect 81176 14172 81240 14176
rect 81176 14116 81180 14172
rect 81180 14116 81236 14172
rect 81236 14116 81240 14172
rect 81176 14112 81240 14116
rect 81256 14172 81320 14176
rect 81256 14116 81260 14172
rect 81260 14116 81316 14172
rect 81316 14116 81320 14172
rect 81256 14112 81320 14116
rect 111736 14172 111800 14176
rect 111736 14116 111740 14172
rect 111740 14116 111796 14172
rect 111796 14116 111800 14172
rect 111736 14112 111800 14116
rect 111816 14172 111880 14176
rect 111816 14116 111820 14172
rect 111820 14116 111876 14172
rect 111876 14116 111880 14172
rect 111816 14112 111880 14116
rect 111896 14172 111960 14176
rect 111896 14116 111900 14172
rect 111900 14116 111956 14172
rect 111956 14116 111960 14172
rect 111896 14112 111960 14116
rect 111976 14172 112040 14176
rect 111976 14116 111980 14172
rect 111980 14116 112036 14172
rect 112036 14116 112040 14172
rect 111976 14112 112040 14116
rect 142456 14172 142520 14176
rect 142456 14116 142460 14172
rect 142460 14116 142516 14172
rect 142516 14116 142520 14172
rect 142456 14112 142520 14116
rect 142536 14172 142600 14176
rect 142536 14116 142540 14172
rect 142540 14116 142596 14172
rect 142596 14116 142600 14172
rect 142536 14112 142600 14116
rect 142616 14172 142680 14176
rect 142616 14116 142620 14172
rect 142620 14116 142676 14172
rect 142676 14116 142680 14172
rect 142616 14112 142680 14116
rect 142696 14172 142760 14176
rect 142696 14116 142700 14172
rect 142700 14116 142756 14172
rect 142756 14116 142760 14172
rect 142696 14112 142760 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 65656 13628 65720 13632
rect 65656 13572 65660 13628
rect 65660 13572 65716 13628
rect 65716 13572 65720 13628
rect 65656 13568 65720 13572
rect 65736 13628 65800 13632
rect 65736 13572 65740 13628
rect 65740 13572 65796 13628
rect 65796 13572 65800 13628
rect 65736 13568 65800 13572
rect 65816 13628 65880 13632
rect 65816 13572 65820 13628
rect 65820 13572 65876 13628
rect 65876 13572 65880 13628
rect 65816 13568 65880 13572
rect 65896 13628 65960 13632
rect 65896 13572 65900 13628
rect 65900 13572 65956 13628
rect 65956 13572 65960 13628
rect 65896 13568 65960 13572
rect 96376 13628 96440 13632
rect 96376 13572 96380 13628
rect 96380 13572 96436 13628
rect 96436 13572 96440 13628
rect 96376 13568 96440 13572
rect 96456 13628 96520 13632
rect 96456 13572 96460 13628
rect 96460 13572 96516 13628
rect 96516 13572 96520 13628
rect 96456 13568 96520 13572
rect 96536 13628 96600 13632
rect 96536 13572 96540 13628
rect 96540 13572 96596 13628
rect 96596 13572 96600 13628
rect 96536 13568 96600 13572
rect 96616 13628 96680 13632
rect 96616 13572 96620 13628
rect 96620 13572 96676 13628
rect 96676 13572 96680 13628
rect 96616 13568 96680 13572
rect 127096 13628 127160 13632
rect 127096 13572 127100 13628
rect 127100 13572 127156 13628
rect 127156 13572 127160 13628
rect 127096 13568 127160 13572
rect 127176 13628 127240 13632
rect 127176 13572 127180 13628
rect 127180 13572 127236 13628
rect 127236 13572 127240 13628
rect 127176 13568 127240 13572
rect 127256 13628 127320 13632
rect 127256 13572 127260 13628
rect 127260 13572 127316 13628
rect 127316 13572 127320 13628
rect 127256 13568 127320 13572
rect 127336 13628 127400 13632
rect 127336 13572 127340 13628
rect 127340 13572 127396 13628
rect 127396 13572 127400 13628
rect 127336 13568 127400 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 81016 13084 81080 13088
rect 81016 13028 81020 13084
rect 81020 13028 81076 13084
rect 81076 13028 81080 13084
rect 81016 13024 81080 13028
rect 81096 13084 81160 13088
rect 81096 13028 81100 13084
rect 81100 13028 81156 13084
rect 81156 13028 81160 13084
rect 81096 13024 81160 13028
rect 81176 13084 81240 13088
rect 81176 13028 81180 13084
rect 81180 13028 81236 13084
rect 81236 13028 81240 13084
rect 81176 13024 81240 13028
rect 81256 13084 81320 13088
rect 81256 13028 81260 13084
rect 81260 13028 81316 13084
rect 81316 13028 81320 13084
rect 81256 13024 81320 13028
rect 111736 13084 111800 13088
rect 111736 13028 111740 13084
rect 111740 13028 111796 13084
rect 111796 13028 111800 13084
rect 111736 13024 111800 13028
rect 111816 13084 111880 13088
rect 111816 13028 111820 13084
rect 111820 13028 111876 13084
rect 111876 13028 111880 13084
rect 111816 13024 111880 13028
rect 111896 13084 111960 13088
rect 111896 13028 111900 13084
rect 111900 13028 111956 13084
rect 111956 13028 111960 13084
rect 111896 13024 111960 13028
rect 111976 13084 112040 13088
rect 111976 13028 111980 13084
rect 111980 13028 112036 13084
rect 112036 13028 112040 13084
rect 111976 13024 112040 13028
rect 142456 13084 142520 13088
rect 142456 13028 142460 13084
rect 142460 13028 142516 13084
rect 142516 13028 142520 13084
rect 142456 13024 142520 13028
rect 142536 13084 142600 13088
rect 142536 13028 142540 13084
rect 142540 13028 142596 13084
rect 142596 13028 142600 13084
rect 142536 13024 142600 13028
rect 142616 13084 142680 13088
rect 142616 13028 142620 13084
rect 142620 13028 142676 13084
rect 142676 13028 142680 13084
rect 142616 13024 142680 13028
rect 142696 13084 142760 13088
rect 142696 13028 142700 13084
rect 142700 13028 142756 13084
rect 142756 13028 142760 13084
rect 142696 13024 142760 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 65656 12540 65720 12544
rect 65656 12484 65660 12540
rect 65660 12484 65716 12540
rect 65716 12484 65720 12540
rect 65656 12480 65720 12484
rect 65736 12540 65800 12544
rect 65736 12484 65740 12540
rect 65740 12484 65796 12540
rect 65796 12484 65800 12540
rect 65736 12480 65800 12484
rect 65816 12540 65880 12544
rect 65816 12484 65820 12540
rect 65820 12484 65876 12540
rect 65876 12484 65880 12540
rect 65816 12480 65880 12484
rect 65896 12540 65960 12544
rect 65896 12484 65900 12540
rect 65900 12484 65956 12540
rect 65956 12484 65960 12540
rect 65896 12480 65960 12484
rect 96376 12540 96440 12544
rect 96376 12484 96380 12540
rect 96380 12484 96436 12540
rect 96436 12484 96440 12540
rect 96376 12480 96440 12484
rect 96456 12540 96520 12544
rect 96456 12484 96460 12540
rect 96460 12484 96516 12540
rect 96516 12484 96520 12540
rect 96456 12480 96520 12484
rect 96536 12540 96600 12544
rect 96536 12484 96540 12540
rect 96540 12484 96596 12540
rect 96596 12484 96600 12540
rect 96536 12480 96600 12484
rect 96616 12540 96680 12544
rect 96616 12484 96620 12540
rect 96620 12484 96676 12540
rect 96676 12484 96680 12540
rect 96616 12480 96680 12484
rect 127096 12540 127160 12544
rect 127096 12484 127100 12540
rect 127100 12484 127156 12540
rect 127156 12484 127160 12540
rect 127096 12480 127160 12484
rect 127176 12540 127240 12544
rect 127176 12484 127180 12540
rect 127180 12484 127236 12540
rect 127236 12484 127240 12540
rect 127176 12480 127240 12484
rect 127256 12540 127320 12544
rect 127256 12484 127260 12540
rect 127260 12484 127316 12540
rect 127316 12484 127320 12540
rect 127256 12480 127320 12484
rect 127336 12540 127400 12544
rect 127336 12484 127340 12540
rect 127340 12484 127396 12540
rect 127396 12484 127400 12540
rect 127336 12480 127400 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 81016 11996 81080 12000
rect 81016 11940 81020 11996
rect 81020 11940 81076 11996
rect 81076 11940 81080 11996
rect 81016 11936 81080 11940
rect 81096 11996 81160 12000
rect 81096 11940 81100 11996
rect 81100 11940 81156 11996
rect 81156 11940 81160 11996
rect 81096 11936 81160 11940
rect 81176 11996 81240 12000
rect 81176 11940 81180 11996
rect 81180 11940 81236 11996
rect 81236 11940 81240 11996
rect 81176 11936 81240 11940
rect 81256 11996 81320 12000
rect 81256 11940 81260 11996
rect 81260 11940 81316 11996
rect 81316 11940 81320 11996
rect 81256 11936 81320 11940
rect 111736 11996 111800 12000
rect 111736 11940 111740 11996
rect 111740 11940 111796 11996
rect 111796 11940 111800 11996
rect 111736 11936 111800 11940
rect 111816 11996 111880 12000
rect 111816 11940 111820 11996
rect 111820 11940 111876 11996
rect 111876 11940 111880 11996
rect 111816 11936 111880 11940
rect 111896 11996 111960 12000
rect 111896 11940 111900 11996
rect 111900 11940 111956 11996
rect 111956 11940 111960 11996
rect 111896 11936 111960 11940
rect 111976 11996 112040 12000
rect 111976 11940 111980 11996
rect 111980 11940 112036 11996
rect 112036 11940 112040 11996
rect 111976 11936 112040 11940
rect 142456 11996 142520 12000
rect 142456 11940 142460 11996
rect 142460 11940 142516 11996
rect 142516 11940 142520 11996
rect 142456 11936 142520 11940
rect 142536 11996 142600 12000
rect 142536 11940 142540 11996
rect 142540 11940 142596 11996
rect 142596 11940 142600 11996
rect 142536 11936 142600 11940
rect 142616 11996 142680 12000
rect 142616 11940 142620 11996
rect 142620 11940 142676 11996
rect 142676 11940 142680 11996
rect 142616 11936 142680 11940
rect 142696 11996 142760 12000
rect 142696 11940 142700 11996
rect 142700 11940 142756 11996
rect 142756 11940 142760 11996
rect 142696 11936 142760 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 65656 11452 65720 11456
rect 65656 11396 65660 11452
rect 65660 11396 65716 11452
rect 65716 11396 65720 11452
rect 65656 11392 65720 11396
rect 65736 11452 65800 11456
rect 65736 11396 65740 11452
rect 65740 11396 65796 11452
rect 65796 11396 65800 11452
rect 65736 11392 65800 11396
rect 65816 11452 65880 11456
rect 65816 11396 65820 11452
rect 65820 11396 65876 11452
rect 65876 11396 65880 11452
rect 65816 11392 65880 11396
rect 65896 11452 65960 11456
rect 65896 11396 65900 11452
rect 65900 11396 65956 11452
rect 65956 11396 65960 11452
rect 65896 11392 65960 11396
rect 96376 11452 96440 11456
rect 96376 11396 96380 11452
rect 96380 11396 96436 11452
rect 96436 11396 96440 11452
rect 96376 11392 96440 11396
rect 96456 11452 96520 11456
rect 96456 11396 96460 11452
rect 96460 11396 96516 11452
rect 96516 11396 96520 11452
rect 96456 11392 96520 11396
rect 96536 11452 96600 11456
rect 96536 11396 96540 11452
rect 96540 11396 96596 11452
rect 96596 11396 96600 11452
rect 96536 11392 96600 11396
rect 96616 11452 96680 11456
rect 96616 11396 96620 11452
rect 96620 11396 96676 11452
rect 96676 11396 96680 11452
rect 96616 11392 96680 11396
rect 127096 11452 127160 11456
rect 127096 11396 127100 11452
rect 127100 11396 127156 11452
rect 127156 11396 127160 11452
rect 127096 11392 127160 11396
rect 127176 11452 127240 11456
rect 127176 11396 127180 11452
rect 127180 11396 127236 11452
rect 127236 11396 127240 11452
rect 127176 11392 127240 11396
rect 127256 11452 127320 11456
rect 127256 11396 127260 11452
rect 127260 11396 127316 11452
rect 127316 11396 127320 11452
rect 127256 11392 127320 11396
rect 127336 11452 127400 11456
rect 127336 11396 127340 11452
rect 127340 11396 127396 11452
rect 127396 11396 127400 11452
rect 127336 11392 127400 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 81016 10908 81080 10912
rect 81016 10852 81020 10908
rect 81020 10852 81076 10908
rect 81076 10852 81080 10908
rect 81016 10848 81080 10852
rect 81096 10908 81160 10912
rect 81096 10852 81100 10908
rect 81100 10852 81156 10908
rect 81156 10852 81160 10908
rect 81096 10848 81160 10852
rect 81176 10908 81240 10912
rect 81176 10852 81180 10908
rect 81180 10852 81236 10908
rect 81236 10852 81240 10908
rect 81176 10848 81240 10852
rect 81256 10908 81320 10912
rect 81256 10852 81260 10908
rect 81260 10852 81316 10908
rect 81316 10852 81320 10908
rect 81256 10848 81320 10852
rect 111736 10908 111800 10912
rect 111736 10852 111740 10908
rect 111740 10852 111796 10908
rect 111796 10852 111800 10908
rect 111736 10848 111800 10852
rect 111816 10908 111880 10912
rect 111816 10852 111820 10908
rect 111820 10852 111876 10908
rect 111876 10852 111880 10908
rect 111816 10848 111880 10852
rect 111896 10908 111960 10912
rect 111896 10852 111900 10908
rect 111900 10852 111956 10908
rect 111956 10852 111960 10908
rect 111896 10848 111960 10852
rect 111976 10908 112040 10912
rect 111976 10852 111980 10908
rect 111980 10852 112036 10908
rect 112036 10852 112040 10908
rect 111976 10848 112040 10852
rect 142456 10908 142520 10912
rect 142456 10852 142460 10908
rect 142460 10852 142516 10908
rect 142516 10852 142520 10908
rect 142456 10848 142520 10852
rect 142536 10908 142600 10912
rect 142536 10852 142540 10908
rect 142540 10852 142596 10908
rect 142596 10852 142600 10908
rect 142536 10848 142600 10852
rect 142616 10908 142680 10912
rect 142616 10852 142620 10908
rect 142620 10852 142676 10908
rect 142676 10852 142680 10908
rect 142616 10848 142680 10852
rect 142696 10908 142760 10912
rect 142696 10852 142700 10908
rect 142700 10852 142756 10908
rect 142756 10852 142760 10908
rect 142696 10848 142760 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 65656 10364 65720 10368
rect 65656 10308 65660 10364
rect 65660 10308 65716 10364
rect 65716 10308 65720 10364
rect 65656 10304 65720 10308
rect 65736 10364 65800 10368
rect 65736 10308 65740 10364
rect 65740 10308 65796 10364
rect 65796 10308 65800 10364
rect 65736 10304 65800 10308
rect 65816 10364 65880 10368
rect 65816 10308 65820 10364
rect 65820 10308 65876 10364
rect 65876 10308 65880 10364
rect 65816 10304 65880 10308
rect 65896 10364 65960 10368
rect 65896 10308 65900 10364
rect 65900 10308 65956 10364
rect 65956 10308 65960 10364
rect 65896 10304 65960 10308
rect 96376 10364 96440 10368
rect 96376 10308 96380 10364
rect 96380 10308 96436 10364
rect 96436 10308 96440 10364
rect 96376 10304 96440 10308
rect 96456 10364 96520 10368
rect 96456 10308 96460 10364
rect 96460 10308 96516 10364
rect 96516 10308 96520 10364
rect 96456 10304 96520 10308
rect 96536 10364 96600 10368
rect 96536 10308 96540 10364
rect 96540 10308 96596 10364
rect 96596 10308 96600 10364
rect 96536 10304 96600 10308
rect 96616 10364 96680 10368
rect 96616 10308 96620 10364
rect 96620 10308 96676 10364
rect 96676 10308 96680 10364
rect 96616 10304 96680 10308
rect 127096 10364 127160 10368
rect 127096 10308 127100 10364
rect 127100 10308 127156 10364
rect 127156 10308 127160 10364
rect 127096 10304 127160 10308
rect 127176 10364 127240 10368
rect 127176 10308 127180 10364
rect 127180 10308 127236 10364
rect 127236 10308 127240 10364
rect 127176 10304 127240 10308
rect 127256 10364 127320 10368
rect 127256 10308 127260 10364
rect 127260 10308 127316 10364
rect 127316 10308 127320 10364
rect 127256 10304 127320 10308
rect 127336 10364 127400 10368
rect 127336 10308 127340 10364
rect 127340 10308 127396 10364
rect 127396 10308 127400 10364
rect 127336 10304 127400 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 81016 9820 81080 9824
rect 81016 9764 81020 9820
rect 81020 9764 81076 9820
rect 81076 9764 81080 9820
rect 81016 9760 81080 9764
rect 81096 9820 81160 9824
rect 81096 9764 81100 9820
rect 81100 9764 81156 9820
rect 81156 9764 81160 9820
rect 81096 9760 81160 9764
rect 81176 9820 81240 9824
rect 81176 9764 81180 9820
rect 81180 9764 81236 9820
rect 81236 9764 81240 9820
rect 81176 9760 81240 9764
rect 81256 9820 81320 9824
rect 81256 9764 81260 9820
rect 81260 9764 81316 9820
rect 81316 9764 81320 9820
rect 81256 9760 81320 9764
rect 111736 9820 111800 9824
rect 111736 9764 111740 9820
rect 111740 9764 111796 9820
rect 111796 9764 111800 9820
rect 111736 9760 111800 9764
rect 111816 9820 111880 9824
rect 111816 9764 111820 9820
rect 111820 9764 111876 9820
rect 111876 9764 111880 9820
rect 111816 9760 111880 9764
rect 111896 9820 111960 9824
rect 111896 9764 111900 9820
rect 111900 9764 111956 9820
rect 111956 9764 111960 9820
rect 111896 9760 111960 9764
rect 111976 9820 112040 9824
rect 111976 9764 111980 9820
rect 111980 9764 112036 9820
rect 112036 9764 112040 9820
rect 111976 9760 112040 9764
rect 142456 9820 142520 9824
rect 142456 9764 142460 9820
rect 142460 9764 142516 9820
rect 142516 9764 142520 9820
rect 142456 9760 142520 9764
rect 142536 9820 142600 9824
rect 142536 9764 142540 9820
rect 142540 9764 142596 9820
rect 142596 9764 142600 9820
rect 142536 9760 142600 9764
rect 142616 9820 142680 9824
rect 142616 9764 142620 9820
rect 142620 9764 142676 9820
rect 142676 9764 142680 9820
rect 142616 9760 142680 9764
rect 142696 9820 142760 9824
rect 142696 9764 142700 9820
rect 142700 9764 142756 9820
rect 142756 9764 142760 9820
rect 142696 9760 142760 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 65656 9276 65720 9280
rect 65656 9220 65660 9276
rect 65660 9220 65716 9276
rect 65716 9220 65720 9276
rect 65656 9216 65720 9220
rect 65736 9276 65800 9280
rect 65736 9220 65740 9276
rect 65740 9220 65796 9276
rect 65796 9220 65800 9276
rect 65736 9216 65800 9220
rect 65816 9276 65880 9280
rect 65816 9220 65820 9276
rect 65820 9220 65876 9276
rect 65876 9220 65880 9276
rect 65816 9216 65880 9220
rect 65896 9276 65960 9280
rect 65896 9220 65900 9276
rect 65900 9220 65956 9276
rect 65956 9220 65960 9276
rect 65896 9216 65960 9220
rect 96376 9276 96440 9280
rect 96376 9220 96380 9276
rect 96380 9220 96436 9276
rect 96436 9220 96440 9276
rect 96376 9216 96440 9220
rect 96456 9276 96520 9280
rect 96456 9220 96460 9276
rect 96460 9220 96516 9276
rect 96516 9220 96520 9276
rect 96456 9216 96520 9220
rect 96536 9276 96600 9280
rect 96536 9220 96540 9276
rect 96540 9220 96596 9276
rect 96596 9220 96600 9276
rect 96536 9216 96600 9220
rect 96616 9276 96680 9280
rect 96616 9220 96620 9276
rect 96620 9220 96676 9276
rect 96676 9220 96680 9276
rect 96616 9216 96680 9220
rect 127096 9276 127160 9280
rect 127096 9220 127100 9276
rect 127100 9220 127156 9276
rect 127156 9220 127160 9276
rect 127096 9216 127160 9220
rect 127176 9276 127240 9280
rect 127176 9220 127180 9276
rect 127180 9220 127236 9276
rect 127236 9220 127240 9276
rect 127176 9216 127240 9220
rect 127256 9276 127320 9280
rect 127256 9220 127260 9276
rect 127260 9220 127316 9276
rect 127316 9220 127320 9276
rect 127256 9216 127320 9220
rect 127336 9276 127400 9280
rect 127336 9220 127340 9276
rect 127340 9220 127396 9276
rect 127396 9220 127400 9276
rect 127336 9216 127400 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 81016 8732 81080 8736
rect 81016 8676 81020 8732
rect 81020 8676 81076 8732
rect 81076 8676 81080 8732
rect 81016 8672 81080 8676
rect 81096 8732 81160 8736
rect 81096 8676 81100 8732
rect 81100 8676 81156 8732
rect 81156 8676 81160 8732
rect 81096 8672 81160 8676
rect 81176 8732 81240 8736
rect 81176 8676 81180 8732
rect 81180 8676 81236 8732
rect 81236 8676 81240 8732
rect 81176 8672 81240 8676
rect 81256 8732 81320 8736
rect 81256 8676 81260 8732
rect 81260 8676 81316 8732
rect 81316 8676 81320 8732
rect 81256 8672 81320 8676
rect 111736 8732 111800 8736
rect 111736 8676 111740 8732
rect 111740 8676 111796 8732
rect 111796 8676 111800 8732
rect 111736 8672 111800 8676
rect 111816 8732 111880 8736
rect 111816 8676 111820 8732
rect 111820 8676 111876 8732
rect 111876 8676 111880 8732
rect 111816 8672 111880 8676
rect 111896 8732 111960 8736
rect 111896 8676 111900 8732
rect 111900 8676 111956 8732
rect 111956 8676 111960 8732
rect 111896 8672 111960 8676
rect 111976 8732 112040 8736
rect 111976 8676 111980 8732
rect 111980 8676 112036 8732
rect 112036 8676 112040 8732
rect 111976 8672 112040 8676
rect 142456 8732 142520 8736
rect 142456 8676 142460 8732
rect 142460 8676 142516 8732
rect 142516 8676 142520 8732
rect 142456 8672 142520 8676
rect 142536 8732 142600 8736
rect 142536 8676 142540 8732
rect 142540 8676 142596 8732
rect 142596 8676 142600 8732
rect 142536 8672 142600 8676
rect 142616 8732 142680 8736
rect 142616 8676 142620 8732
rect 142620 8676 142676 8732
rect 142676 8676 142680 8732
rect 142616 8672 142680 8676
rect 142696 8732 142760 8736
rect 142696 8676 142700 8732
rect 142700 8676 142756 8732
rect 142756 8676 142760 8732
rect 142696 8672 142760 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 65656 8188 65720 8192
rect 65656 8132 65660 8188
rect 65660 8132 65716 8188
rect 65716 8132 65720 8188
rect 65656 8128 65720 8132
rect 65736 8188 65800 8192
rect 65736 8132 65740 8188
rect 65740 8132 65796 8188
rect 65796 8132 65800 8188
rect 65736 8128 65800 8132
rect 65816 8188 65880 8192
rect 65816 8132 65820 8188
rect 65820 8132 65876 8188
rect 65876 8132 65880 8188
rect 65816 8128 65880 8132
rect 65896 8188 65960 8192
rect 65896 8132 65900 8188
rect 65900 8132 65956 8188
rect 65956 8132 65960 8188
rect 65896 8128 65960 8132
rect 96376 8188 96440 8192
rect 96376 8132 96380 8188
rect 96380 8132 96436 8188
rect 96436 8132 96440 8188
rect 96376 8128 96440 8132
rect 96456 8188 96520 8192
rect 96456 8132 96460 8188
rect 96460 8132 96516 8188
rect 96516 8132 96520 8188
rect 96456 8128 96520 8132
rect 96536 8188 96600 8192
rect 96536 8132 96540 8188
rect 96540 8132 96596 8188
rect 96596 8132 96600 8188
rect 96536 8128 96600 8132
rect 96616 8188 96680 8192
rect 96616 8132 96620 8188
rect 96620 8132 96676 8188
rect 96676 8132 96680 8188
rect 96616 8128 96680 8132
rect 127096 8188 127160 8192
rect 127096 8132 127100 8188
rect 127100 8132 127156 8188
rect 127156 8132 127160 8188
rect 127096 8128 127160 8132
rect 127176 8188 127240 8192
rect 127176 8132 127180 8188
rect 127180 8132 127236 8188
rect 127236 8132 127240 8188
rect 127176 8128 127240 8132
rect 127256 8188 127320 8192
rect 127256 8132 127260 8188
rect 127260 8132 127316 8188
rect 127316 8132 127320 8188
rect 127256 8128 127320 8132
rect 127336 8188 127400 8192
rect 127336 8132 127340 8188
rect 127340 8132 127396 8188
rect 127396 8132 127400 8188
rect 127336 8128 127400 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 81016 7644 81080 7648
rect 81016 7588 81020 7644
rect 81020 7588 81076 7644
rect 81076 7588 81080 7644
rect 81016 7584 81080 7588
rect 81096 7644 81160 7648
rect 81096 7588 81100 7644
rect 81100 7588 81156 7644
rect 81156 7588 81160 7644
rect 81096 7584 81160 7588
rect 81176 7644 81240 7648
rect 81176 7588 81180 7644
rect 81180 7588 81236 7644
rect 81236 7588 81240 7644
rect 81176 7584 81240 7588
rect 81256 7644 81320 7648
rect 81256 7588 81260 7644
rect 81260 7588 81316 7644
rect 81316 7588 81320 7644
rect 81256 7584 81320 7588
rect 111736 7644 111800 7648
rect 111736 7588 111740 7644
rect 111740 7588 111796 7644
rect 111796 7588 111800 7644
rect 111736 7584 111800 7588
rect 111816 7644 111880 7648
rect 111816 7588 111820 7644
rect 111820 7588 111876 7644
rect 111876 7588 111880 7644
rect 111816 7584 111880 7588
rect 111896 7644 111960 7648
rect 111896 7588 111900 7644
rect 111900 7588 111956 7644
rect 111956 7588 111960 7644
rect 111896 7584 111960 7588
rect 111976 7644 112040 7648
rect 111976 7588 111980 7644
rect 111980 7588 112036 7644
rect 112036 7588 112040 7644
rect 111976 7584 112040 7588
rect 142456 7644 142520 7648
rect 142456 7588 142460 7644
rect 142460 7588 142516 7644
rect 142516 7588 142520 7644
rect 142456 7584 142520 7588
rect 142536 7644 142600 7648
rect 142536 7588 142540 7644
rect 142540 7588 142596 7644
rect 142596 7588 142600 7644
rect 142536 7584 142600 7588
rect 142616 7644 142680 7648
rect 142616 7588 142620 7644
rect 142620 7588 142676 7644
rect 142676 7588 142680 7644
rect 142616 7584 142680 7588
rect 142696 7644 142760 7648
rect 142696 7588 142700 7644
rect 142700 7588 142756 7644
rect 142756 7588 142760 7644
rect 142696 7584 142760 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 65656 7100 65720 7104
rect 65656 7044 65660 7100
rect 65660 7044 65716 7100
rect 65716 7044 65720 7100
rect 65656 7040 65720 7044
rect 65736 7100 65800 7104
rect 65736 7044 65740 7100
rect 65740 7044 65796 7100
rect 65796 7044 65800 7100
rect 65736 7040 65800 7044
rect 65816 7100 65880 7104
rect 65816 7044 65820 7100
rect 65820 7044 65876 7100
rect 65876 7044 65880 7100
rect 65816 7040 65880 7044
rect 65896 7100 65960 7104
rect 65896 7044 65900 7100
rect 65900 7044 65956 7100
rect 65956 7044 65960 7100
rect 65896 7040 65960 7044
rect 96376 7100 96440 7104
rect 96376 7044 96380 7100
rect 96380 7044 96436 7100
rect 96436 7044 96440 7100
rect 96376 7040 96440 7044
rect 96456 7100 96520 7104
rect 96456 7044 96460 7100
rect 96460 7044 96516 7100
rect 96516 7044 96520 7100
rect 96456 7040 96520 7044
rect 96536 7100 96600 7104
rect 96536 7044 96540 7100
rect 96540 7044 96596 7100
rect 96596 7044 96600 7100
rect 96536 7040 96600 7044
rect 96616 7100 96680 7104
rect 96616 7044 96620 7100
rect 96620 7044 96676 7100
rect 96676 7044 96680 7100
rect 96616 7040 96680 7044
rect 127096 7100 127160 7104
rect 127096 7044 127100 7100
rect 127100 7044 127156 7100
rect 127156 7044 127160 7100
rect 127096 7040 127160 7044
rect 127176 7100 127240 7104
rect 127176 7044 127180 7100
rect 127180 7044 127236 7100
rect 127236 7044 127240 7100
rect 127176 7040 127240 7044
rect 127256 7100 127320 7104
rect 127256 7044 127260 7100
rect 127260 7044 127316 7100
rect 127316 7044 127320 7100
rect 127256 7040 127320 7044
rect 127336 7100 127400 7104
rect 127336 7044 127340 7100
rect 127340 7044 127396 7100
rect 127396 7044 127400 7100
rect 127336 7040 127400 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 81016 6556 81080 6560
rect 81016 6500 81020 6556
rect 81020 6500 81076 6556
rect 81076 6500 81080 6556
rect 81016 6496 81080 6500
rect 81096 6556 81160 6560
rect 81096 6500 81100 6556
rect 81100 6500 81156 6556
rect 81156 6500 81160 6556
rect 81096 6496 81160 6500
rect 81176 6556 81240 6560
rect 81176 6500 81180 6556
rect 81180 6500 81236 6556
rect 81236 6500 81240 6556
rect 81176 6496 81240 6500
rect 81256 6556 81320 6560
rect 81256 6500 81260 6556
rect 81260 6500 81316 6556
rect 81316 6500 81320 6556
rect 81256 6496 81320 6500
rect 111736 6556 111800 6560
rect 111736 6500 111740 6556
rect 111740 6500 111796 6556
rect 111796 6500 111800 6556
rect 111736 6496 111800 6500
rect 111816 6556 111880 6560
rect 111816 6500 111820 6556
rect 111820 6500 111876 6556
rect 111876 6500 111880 6556
rect 111816 6496 111880 6500
rect 111896 6556 111960 6560
rect 111896 6500 111900 6556
rect 111900 6500 111956 6556
rect 111956 6500 111960 6556
rect 111896 6496 111960 6500
rect 111976 6556 112040 6560
rect 111976 6500 111980 6556
rect 111980 6500 112036 6556
rect 112036 6500 112040 6556
rect 111976 6496 112040 6500
rect 142456 6556 142520 6560
rect 142456 6500 142460 6556
rect 142460 6500 142516 6556
rect 142516 6500 142520 6556
rect 142456 6496 142520 6500
rect 142536 6556 142600 6560
rect 142536 6500 142540 6556
rect 142540 6500 142596 6556
rect 142596 6500 142600 6556
rect 142536 6496 142600 6500
rect 142616 6556 142680 6560
rect 142616 6500 142620 6556
rect 142620 6500 142676 6556
rect 142676 6500 142680 6556
rect 142616 6496 142680 6500
rect 142696 6556 142760 6560
rect 142696 6500 142700 6556
rect 142700 6500 142756 6556
rect 142756 6500 142760 6556
rect 142696 6496 142760 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 65656 6012 65720 6016
rect 65656 5956 65660 6012
rect 65660 5956 65716 6012
rect 65716 5956 65720 6012
rect 65656 5952 65720 5956
rect 65736 6012 65800 6016
rect 65736 5956 65740 6012
rect 65740 5956 65796 6012
rect 65796 5956 65800 6012
rect 65736 5952 65800 5956
rect 65816 6012 65880 6016
rect 65816 5956 65820 6012
rect 65820 5956 65876 6012
rect 65876 5956 65880 6012
rect 65816 5952 65880 5956
rect 65896 6012 65960 6016
rect 65896 5956 65900 6012
rect 65900 5956 65956 6012
rect 65956 5956 65960 6012
rect 65896 5952 65960 5956
rect 96376 6012 96440 6016
rect 96376 5956 96380 6012
rect 96380 5956 96436 6012
rect 96436 5956 96440 6012
rect 96376 5952 96440 5956
rect 96456 6012 96520 6016
rect 96456 5956 96460 6012
rect 96460 5956 96516 6012
rect 96516 5956 96520 6012
rect 96456 5952 96520 5956
rect 96536 6012 96600 6016
rect 96536 5956 96540 6012
rect 96540 5956 96596 6012
rect 96596 5956 96600 6012
rect 96536 5952 96600 5956
rect 96616 6012 96680 6016
rect 96616 5956 96620 6012
rect 96620 5956 96676 6012
rect 96676 5956 96680 6012
rect 96616 5952 96680 5956
rect 127096 6012 127160 6016
rect 127096 5956 127100 6012
rect 127100 5956 127156 6012
rect 127156 5956 127160 6012
rect 127096 5952 127160 5956
rect 127176 6012 127240 6016
rect 127176 5956 127180 6012
rect 127180 5956 127236 6012
rect 127236 5956 127240 6012
rect 127176 5952 127240 5956
rect 127256 6012 127320 6016
rect 127256 5956 127260 6012
rect 127260 5956 127316 6012
rect 127316 5956 127320 6012
rect 127256 5952 127320 5956
rect 127336 6012 127400 6016
rect 127336 5956 127340 6012
rect 127340 5956 127396 6012
rect 127396 5956 127400 6012
rect 127336 5952 127400 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 81016 5468 81080 5472
rect 81016 5412 81020 5468
rect 81020 5412 81076 5468
rect 81076 5412 81080 5468
rect 81016 5408 81080 5412
rect 81096 5468 81160 5472
rect 81096 5412 81100 5468
rect 81100 5412 81156 5468
rect 81156 5412 81160 5468
rect 81096 5408 81160 5412
rect 81176 5468 81240 5472
rect 81176 5412 81180 5468
rect 81180 5412 81236 5468
rect 81236 5412 81240 5468
rect 81176 5408 81240 5412
rect 81256 5468 81320 5472
rect 81256 5412 81260 5468
rect 81260 5412 81316 5468
rect 81316 5412 81320 5468
rect 81256 5408 81320 5412
rect 111736 5468 111800 5472
rect 111736 5412 111740 5468
rect 111740 5412 111796 5468
rect 111796 5412 111800 5468
rect 111736 5408 111800 5412
rect 111816 5468 111880 5472
rect 111816 5412 111820 5468
rect 111820 5412 111876 5468
rect 111876 5412 111880 5468
rect 111816 5408 111880 5412
rect 111896 5468 111960 5472
rect 111896 5412 111900 5468
rect 111900 5412 111956 5468
rect 111956 5412 111960 5468
rect 111896 5408 111960 5412
rect 111976 5468 112040 5472
rect 111976 5412 111980 5468
rect 111980 5412 112036 5468
rect 112036 5412 112040 5468
rect 111976 5408 112040 5412
rect 142456 5468 142520 5472
rect 142456 5412 142460 5468
rect 142460 5412 142516 5468
rect 142516 5412 142520 5468
rect 142456 5408 142520 5412
rect 142536 5468 142600 5472
rect 142536 5412 142540 5468
rect 142540 5412 142596 5468
rect 142596 5412 142600 5468
rect 142536 5408 142600 5412
rect 142616 5468 142680 5472
rect 142616 5412 142620 5468
rect 142620 5412 142676 5468
rect 142676 5412 142680 5468
rect 142616 5408 142680 5412
rect 142696 5468 142760 5472
rect 142696 5412 142700 5468
rect 142700 5412 142756 5468
rect 142756 5412 142760 5468
rect 142696 5408 142760 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 65656 4924 65720 4928
rect 65656 4868 65660 4924
rect 65660 4868 65716 4924
rect 65716 4868 65720 4924
rect 65656 4864 65720 4868
rect 65736 4924 65800 4928
rect 65736 4868 65740 4924
rect 65740 4868 65796 4924
rect 65796 4868 65800 4924
rect 65736 4864 65800 4868
rect 65816 4924 65880 4928
rect 65816 4868 65820 4924
rect 65820 4868 65876 4924
rect 65876 4868 65880 4924
rect 65816 4864 65880 4868
rect 65896 4924 65960 4928
rect 65896 4868 65900 4924
rect 65900 4868 65956 4924
rect 65956 4868 65960 4924
rect 65896 4864 65960 4868
rect 96376 4924 96440 4928
rect 96376 4868 96380 4924
rect 96380 4868 96436 4924
rect 96436 4868 96440 4924
rect 96376 4864 96440 4868
rect 96456 4924 96520 4928
rect 96456 4868 96460 4924
rect 96460 4868 96516 4924
rect 96516 4868 96520 4924
rect 96456 4864 96520 4868
rect 96536 4924 96600 4928
rect 96536 4868 96540 4924
rect 96540 4868 96596 4924
rect 96596 4868 96600 4924
rect 96536 4864 96600 4868
rect 96616 4924 96680 4928
rect 96616 4868 96620 4924
rect 96620 4868 96676 4924
rect 96676 4868 96680 4924
rect 96616 4864 96680 4868
rect 127096 4924 127160 4928
rect 127096 4868 127100 4924
rect 127100 4868 127156 4924
rect 127156 4868 127160 4924
rect 127096 4864 127160 4868
rect 127176 4924 127240 4928
rect 127176 4868 127180 4924
rect 127180 4868 127236 4924
rect 127236 4868 127240 4924
rect 127176 4864 127240 4868
rect 127256 4924 127320 4928
rect 127256 4868 127260 4924
rect 127260 4868 127316 4924
rect 127316 4868 127320 4924
rect 127256 4864 127320 4868
rect 127336 4924 127400 4928
rect 127336 4868 127340 4924
rect 127340 4868 127396 4924
rect 127396 4868 127400 4924
rect 127336 4864 127400 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 81016 4380 81080 4384
rect 81016 4324 81020 4380
rect 81020 4324 81076 4380
rect 81076 4324 81080 4380
rect 81016 4320 81080 4324
rect 81096 4380 81160 4384
rect 81096 4324 81100 4380
rect 81100 4324 81156 4380
rect 81156 4324 81160 4380
rect 81096 4320 81160 4324
rect 81176 4380 81240 4384
rect 81176 4324 81180 4380
rect 81180 4324 81236 4380
rect 81236 4324 81240 4380
rect 81176 4320 81240 4324
rect 81256 4380 81320 4384
rect 81256 4324 81260 4380
rect 81260 4324 81316 4380
rect 81316 4324 81320 4380
rect 81256 4320 81320 4324
rect 111736 4380 111800 4384
rect 111736 4324 111740 4380
rect 111740 4324 111796 4380
rect 111796 4324 111800 4380
rect 111736 4320 111800 4324
rect 111816 4380 111880 4384
rect 111816 4324 111820 4380
rect 111820 4324 111876 4380
rect 111876 4324 111880 4380
rect 111816 4320 111880 4324
rect 111896 4380 111960 4384
rect 111896 4324 111900 4380
rect 111900 4324 111956 4380
rect 111956 4324 111960 4380
rect 111896 4320 111960 4324
rect 111976 4380 112040 4384
rect 111976 4324 111980 4380
rect 111980 4324 112036 4380
rect 112036 4324 112040 4380
rect 111976 4320 112040 4324
rect 142456 4380 142520 4384
rect 142456 4324 142460 4380
rect 142460 4324 142516 4380
rect 142516 4324 142520 4380
rect 142456 4320 142520 4324
rect 142536 4380 142600 4384
rect 142536 4324 142540 4380
rect 142540 4324 142596 4380
rect 142596 4324 142600 4380
rect 142536 4320 142600 4324
rect 142616 4380 142680 4384
rect 142616 4324 142620 4380
rect 142620 4324 142676 4380
rect 142676 4324 142680 4380
rect 142616 4320 142680 4324
rect 142696 4380 142760 4384
rect 142696 4324 142700 4380
rect 142700 4324 142756 4380
rect 142756 4324 142760 4380
rect 142696 4320 142760 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 65656 3836 65720 3840
rect 65656 3780 65660 3836
rect 65660 3780 65716 3836
rect 65716 3780 65720 3836
rect 65656 3776 65720 3780
rect 65736 3836 65800 3840
rect 65736 3780 65740 3836
rect 65740 3780 65796 3836
rect 65796 3780 65800 3836
rect 65736 3776 65800 3780
rect 65816 3836 65880 3840
rect 65816 3780 65820 3836
rect 65820 3780 65876 3836
rect 65876 3780 65880 3836
rect 65816 3776 65880 3780
rect 65896 3836 65960 3840
rect 65896 3780 65900 3836
rect 65900 3780 65956 3836
rect 65956 3780 65960 3836
rect 65896 3776 65960 3780
rect 96376 3836 96440 3840
rect 96376 3780 96380 3836
rect 96380 3780 96436 3836
rect 96436 3780 96440 3836
rect 96376 3776 96440 3780
rect 96456 3836 96520 3840
rect 96456 3780 96460 3836
rect 96460 3780 96516 3836
rect 96516 3780 96520 3836
rect 96456 3776 96520 3780
rect 96536 3836 96600 3840
rect 96536 3780 96540 3836
rect 96540 3780 96596 3836
rect 96596 3780 96600 3836
rect 96536 3776 96600 3780
rect 96616 3836 96680 3840
rect 96616 3780 96620 3836
rect 96620 3780 96676 3836
rect 96676 3780 96680 3836
rect 96616 3776 96680 3780
rect 127096 3836 127160 3840
rect 127096 3780 127100 3836
rect 127100 3780 127156 3836
rect 127156 3780 127160 3836
rect 127096 3776 127160 3780
rect 127176 3836 127240 3840
rect 127176 3780 127180 3836
rect 127180 3780 127236 3836
rect 127236 3780 127240 3836
rect 127176 3776 127240 3780
rect 127256 3836 127320 3840
rect 127256 3780 127260 3836
rect 127260 3780 127316 3836
rect 127316 3780 127320 3836
rect 127256 3776 127320 3780
rect 127336 3836 127400 3840
rect 127336 3780 127340 3836
rect 127340 3780 127396 3836
rect 127396 3780 127400 3836
rect 127336 3776 127400 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 81016 3292 81080 3296
rect 81016 3236 81020 3292
rect 81020 3236 81076 3292
rect 81076 3236 81080 3292
rect 81016 3232 81080 3236
rect 81096 3292 81160 3296
rect 81096 3236 81100 3292
rect 81100 3236 81156 3292
rect 81156 3236 81160 3292
rect 81096 3232 81160 3236
rect 81176 3292 81240 3296
rect 81176 3236 81180 3292
rect 81180 3236 81236 3292
rect 81236 3236 81240 3292
rect 81176 3232 81240 3236
rect 81256 3292 81320 3296
rect 81256 3236 81260 3292
rect 81260 3236 81316 3292
rect 81316 3236 81320 3292
rect 81256 3232 81320 3236
rect 111736 3292 111800 3296
rect 111736 3236 111740 3292
rect 111740 3236 111796 3292
rect 111796 3236 111800 3292
rect 111736 3232 111800 3236
rect 111816 3292 111880 3296
rect 111816 3236 111820 3292
rect 111820 3236 111876 3292
rect 111876 3236 111880 3292
rect 111816 3232 111880 3236
rect 111896 3292 111960 3296
rect 111896 3236 111900 3292
rect 111900 3236 111956 3292
rect 111956 3236 111960 3292
rect 111896 3232 111960 3236
rect 111976 3292 112040 3296
rect 111976 3236 111980 3292
rect 111980 3236 112036 3292
rect 112036 3236 112040 3292
rect 111976 3232 112040 3236
rect 142456 3292 142520 3296
rect 142456 3236 142460 3292
rect 142460 3236 142516 3292
rect 142516 3236 142520 3292
rect 142456 3232 142520 3236
rect 142536 3292 142600 3296
rect 142536 3236 142540 3292
rect 142540 3236 142596 3292
rect 142596 3236 142600 3292
rect 142536 3232 142600 3236
rect 142616 3292 142680 3296
rect 142616 3236 142620 3292
rect 142620 3236 142676 3292
rect 142676 3236 142680 3292
rect 142616 3232 142680 3236
rect 142696 3292 142760 3296
rect 142696 3236 142700 3292
rect 142700 3236 142756 3292
rect 142756 3236 142760 3292
rect 142696 3232 142760 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 65656 2748 65720 2752
rect 65656 2692 65660 2748
rect 65660 2692 65716 2748
rect 65716 2692 65720 2748
rect 65656 2688 65720 2692
rect 65736 2748 65800 2752
rect 65736 2692 65740 2748
rect 65740 2692 65796 2748
rect 65796 2692 65800 2748
rect 65736 2688 65800 2692
rect 65816 2748 65880 2752
rect 65816 2692 65820 2748
rect 65820 2692 65876 2748
rect 65876 2692 65880 2748
rect 65816 2688 65880 2692
rect 65896 2748 65960 2752
rect 65896 2692 65900 2748
rect 65900 2692 65956 2748
rect 65956 2692 65960 2748
rect 65896 2688 65960 2692
rect 96376 2748 96440 2752
rect 96376 2692 96380 2748
rect 96380 2692 96436 2748
rect 96436 2692 96440 2748
rect 96376 2688 96440 2692
rect 96456 2748 96520 2752
rect 96456 2692 96460 2748
rect 96460 2692 96516 2748
rect 96516 2692 96520 2748
rect 96456 2688 96520 2692
rect 96536 2748 96600 2752
rect 96536 2692 96540 2748
rect 96540 2692 96596 2748
rect 96596 2692 96600 2748
rect 96536 2688 96600 2692
rect 96616 2748 96680 2752
rect 96616 2692 96620 2748
rect 96620 2692 96676 2748
rect 96676 2692 96680 2748
rect 96616 2688 96680 2692
rect 127096 2748 127160 2752
rect 127096 2692 127100 2748
rect 127100 2692 127156 2748
rect 127156 2692 127160 2748
rect 127096 2688 127160 2692
rect 127176 2748 127240 2752
rect 127176 2692 127180 2748
rect 127180 2692 127236 2748
rect 127236 2692 127240 2748
rect 127176 2688 127240 2692
rect 127256 2748 127320 2752
rect 127256 2692 127260 2748
rect 127260 2692 127316 2748
rect 127316 2692 127320 2748
rect 127256 2688 127320 2692
rect 127336 2748 127400 2752
rect 127336 2692 127340 2748
rect 127340 2692 127396 2748
rect 127396 2692 127400 2748
rect 127336 2688 127400 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
rect 81016 2204 81080 2208
rect 81016 2148 81020 2204
rect 81020 2148 81076 2204
rect 81076 2148 81080 2204
rect 81016 2144 81080 2148
rect 81096 2204 81160 2208
rect 81096 2148 81100 2204
rect 81100 2148 81156 2204
rect 81156 2148 81160 2204
rect 81096 2144 81160 2148
rect 81176 2204 81240 2208
rect 81176 2148 81180 2204
rect 81180 2148 81236 2204
rect 81236 2148 81240 2204
rect 81176 2144 81240 2148
rect 81256 2204 81320 2208
rect 81256 2148 81260 2204
rect 81260 2148 81316 2204
rect 81316 2148 81320 2204
rect 81256 2144 81320 2148
rect 111736 2204 111800 2208
rect 111736 2148 111740 2204
rect 111740 2148 111796 2204
rect 111796 2148 111800 2204
rect 111736 2144 111800 2148
rect 111816 2204 111880 2208
rect 111816 2148 111820 2204
rect 111820 2148 111876 2204
rect 111876 2148 111880 2204
rect 111816 2144 111880 2148
rect 111896 2204 111960 2208
rect 111896 2148 111900 2204
rect 111900 2148 111956 2204
rect 111956 2148 111960 2204
rect 111896 2144 111960 2148
rect 111976 2204 112040 2208
rect 111976 2148 111980 2204
rect 111980 2148 112036 2204
rect 112036 2148 112040 2204
rect 111976 2144 112040 2148
rect 142456 2204 142520 2208
rect 142456 2148 142460 2204
rect 142460 2148 142516 2204
rect 142516 2148 142520 2204
rect 142456 2144 142520 2148
rect 142536 2204 142600 2208
rect 142536 2148 142540 2204
rect 142540 2148 142596 2204
rect 142596 2148 142600 2204
rect 142536 2144 142600 2148
rect 142616 2204 142680 2208
rect 142616 2148 142620 2204
rect 142620 2148 142676 2204
rect 142676 2148 142680 2204
rect 142616 2144 142680 2148
rect 142696 2204 142760 2208
rect 142696 2148 142700 2204
rect 142700 2148 142756 2204
rect 142756 2148 142760 2204
rect 142696 2144 142760 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 37024 50608 37584
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
rect 65648 37568 65968 37584
rect 65648 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65968 37568
rect 65648 36480 65968 37504
rect 65648 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65968 36480
rect 65648 35392 65968 36416
rect 65648 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65968 35392
rect 65648 34304 65968 35328
rect 65648 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65968 34304
rect 65648 33216 65968 34240
rect 65648 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65968 33216
rect 65648 32128 65968 33152
rect 65648 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65968 32128
rect 65648 31040 65968 32064
rect 65648 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65968 31040
rect 65648 29952 65968 30976
rect 65648 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65968 29952
rect 65648 28864 65968 29888
rect 65648 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65968 28864
rect 65648 27776 65968 28800
rect 65648 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65968 27776
rect 65648 26688 65968 27712
rect 65648 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65968 26688
rect 65648 25600 65968 26624
rect 65648 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65968 25600
rect 65648 24512 65968 25536
rect 65648 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65968 24512
rect 65648 23424 65968 24448
rect 65648 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65968 23424
rect 65648 22336 65968 23360
rect 65648 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65968 22336
rect 65648 21248 65968 22272
rect 65648 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65968 21248
rect 65648 20160 65968 21184
rect 65648 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65968 20160
rect 65648 19072 65968 20096
rect 65648 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65968 19072
rect 65648 17984 65968 19008
rect 65648 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65968 17984
rect 65648 16896 65968 17920
rect 65648 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65968 16896
rect 65648 15808 65968 16832
rect 65648 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65968 15808
rect 65648 14720 65968 15744
rect 65648 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65968 14720
rect 65648 13632 65968 14656
rect 65648 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65968 13632
rect 65648 12544 65968 13568
rect 65648 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65968 12544
rect 65648 11456 65968 12480
rect 65648 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65968 11456
rect 65648 10368 65968 11392
rect 65648 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65968 10368
rect 65648 9280 65968 10304
rect 65648 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65968 9280
rect 65648 8192 65968 9216
rect 65648 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65968 8192
rect 65648 7104 65968 8128
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 6016 65968 7040
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 4928 65968 5952
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 65648 3840 65968 4864
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 2752 65968 3776
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 65648 2128 65968 2688
rect 81008 37024 81328 37584
rect 81008 36960 81016 37024
rect 81080 36960 81096 37024
rect 81160 36960 81176 37024
rect 81240 36960 81256 37024
rect 81320 36960 81328 37024
rect 81008 35936 81328 36960
rect 81008 35872 81016 35936
rect 81080 35872 81096 35936
rect 81160 35872 81176 35936
rect 81240 35872 81256 35936
rect 81320 35872 81328 35936
rect 81008 34848 81328 35872
rect 81008 34784 81016 34848
rect 81080 34784 81096 34848
rect 81160 34784 81176 34848
rect 81240 34784 81256 34848
rect 81320 34784 81328 34848
rect 81008 33760 81328 34784
rect 81008 33696 81016 33760
rect 81080 33696 81096 33760
rect 81160 33696 81176 33760
rect 81240 33696 81256 33760
rect 81320 33696 81328 33760
rect 81008 32672 81328 33696
rect 81008 32608 81016 32672
rect 81080 32608 81096 32672
rect 81160 32608 81176 32672
rect 81240 32608 81256 32672
rect 81320 32608 81328 32672
rect 81008 31584 81328 32608
rect 81008 31520 81016 31584
rect 81080 31520 81096 31584
rect 81160 31520 81176 31584
rect 81240 31520 81256 31584
rect 81320 31520 81328 31584
rect 81008 30496 81328 31520
rect 81008 30432 81016 30496
rect 81080 30432 81096 30496
rect 81160 30432 81176 30496
rect 81240 30432 81256 30496
rect 81320 30432 81328 30496
rect 81008 29408 81328 30432
rect 81008 29344 81016 29408
rect 81080 29344 81096 29408
rect 81160 29344 81176 29408
rect 81240 29344 81256 29408
rect 81320 29344 81328 29408
rect 81008 28320 81328 29344
rect 81008 28256 81016 28320
rect 81080 28256 81096 28320
rect 81160 28256 81176 28320
rect 81240 28256 81256 28320
rect 81320 28256 81328 28320
rect 81008 27232 81328 28256
rect 81008 27168 81016 27232
rect 81080 27168 81096 27232
rect 81160 27168 81176 27232
rect 81240 27168 81256 27232
rect 81320 27168 81328 27232
rect 81008 26144 81328 27168
rect 81008 26080 81016 26144
rect 81080 26080 81096 26144
rect 81160 26080 81176 26144
rect 81240 26080 81256 26144
rect 81320 26080 81328 26144
rect 81008 25056 81328 26080
rect 81008 24992 81016 25056
rect 81080 24992 81096 25056
rect 81160 24992 81176 25056
rect 81240 24992 81256 25056
rect 81320 24992 81328 25056
rect 81008 23968 81328 24992
rect 81008 23904 81016 23968
rect 81080 23904 81096 23968
rect 81160 23904 81176 23968
rect 81240 23904 81256 23968
rect 81320 23904 81328 23968
rect 81008 22880 81328 23904
rect 81008 22816 81016 22880
rect 81080 22816 81096 22880
rect 81160 22816 81176 22880
rect 81240 22816 81256 22880
rect 81320 22816 81328 22880
rect 81008 21792 81328 22816
rect 81008 21728 81016 21792
rect 81080 21728 81096 21792
rect 81160 21728 81176 21792
rect 81240 21728 81256 21792
rect 81320 21728 81328 21792
rect 81008 20704 81328 21728
rect 81008 20640 81016 20704
rect 81080 20640 81096 20704
rect 81160 20640 81176 20704
rect 81240 20640 81256 20704
rect 81320 20640 81328 20704
rect 81008 19616 81328 20640
rect 81008 19552 81016 19616
rect 81080 19552 81096 19616
rect 81160 19552 81176 19616
rect 81240 19552 81256 19616
rect 81320 19552 81328 19616
rect 81008 18528 81328 19552
rect 81008 18464 81016 18528
rect 81080 18464 81096 18528
rect 81160 18464 81176 18528
rect 81240 18464 81256 18528
rect 81320 18464 81328 18528
rect 81008 17440 81328 18464
rect 81008 17376 81016 17440
rect 81080 17376 81096 17440
rect 81160 17376 81176 17440
rect 81240 17376 81256 17440
rect 81320 17376 81328 17440
rect 81008 16352 81328 17376
rect 81008 16288 81016 16352
rect 81080 16288 81096 16352
rect 81160 16288 81176 16352
rect 81240 16288 81256 16352
rect 81320 16288 81328 16352
rect 81008 15264 81328 16288
rect 81008 15200 81016 15264
rect 81080 15200 81096 15264
rect 81160 15200 81176 15264
rect 81240 15200 81256 15264
rect 81320 15200 81328 15264
rect 81008 14176 81328 15200
rect 81008 14112 81016 14176
rect 81080 14112 81096 14176
rect 81160 14112 81176 14176
rect 81240 14112 81256 14176
rect 81320 14112 81328 14176
rect 81008 13088 81328 14112
rect 81008 13024 81016 13088
rect 81080 13024 81096 13088
rect 81160 13024 81176 13088
rect 81240 13024 81256 13088
rect 81320 13024 81328 13088
rect 81008 12000 81328 13024
rect 81008 11936 81016 12000
rect 81080 11936 81096 12000
rect 81160 11936 81176 12000
rect 81240 11936 81256 12000
rect 81320 11936 81328 12000
rect 81008 10912 81328 11936
rect 81008 10848 81016 10912
rect 81080 10848 81096 10912
rect 81160 10848 81176 10912
rect 81240 10848 81256 10912
rect 81320 10848 81328 10912
rect 81008 9824 81328 10848
rect 81008 9760 81016 9824
rect 81080 9760 81096 9824
rect 81160 9760 81176 9824
rect 81240 9760 81256 9824
rect 81320 9760 81328 9824
rect 81008 8736 81328 9760
rect 81008 8672 81016 8736
rect 81080 8672 81096 8736
rect 81160 8672 81176 8736
rect 81240 8672 81256 8736
rect 81320 8672 81328 8736
rect 81008 7648 81328 8672
rect 81008 7584 81016 7648
rect 81080 7584 81096 7648
rect 81160 7584 81176 7648
rect 81240 7584 81256 7648
rect 81320 7584 81328 7648
rect 81008 6560 81328 7584
rect 81008 6496 81016 6560
rect 81080 6496 81096 6560
rect 81160 6496 81176 6560
rect 81240 6496 81256 6560
rect 81320 6496 81328 6560
rect 81008 5472 81328 6496
rect 81008 5408 81016 5472
rect 81080 5408 81096 5472
rect 81160 5408 81176 5472
rect 81240 5408 81256 5472
rect 81320 5408 81328 5472
rect 81008 4384 81328 5408
rect 81008 4320 81016 4384
rect 81080 4320 81096 4384
rect 81160 4320 81176 4384
rect 81240 4320 81256 4384
rect 81320 4320 81328 4384
rect 81008 3296 81328 4320
rect 81008 3232 81016 3296
rect 81080 3232 81096 3296
rect 81160 3232 81176 3296
rect 81240 3232 81256 3296
rect 81320 3232 81328 3296
rect 81008 2208 81328 3232
rect 81008 2144 81016 2208
rect 81080 2144 81096 2208
rect 81160 2144 81176 2208
rect 81240 2144 81256 2208
rect 81320 2144 81328 2208
rect 81008 2128 81328 2144
rect 96368 37568 96688 37584
rect 96368 37504 96376 37568
rect 96440 37504 96456 37568
rect 96520 37504 96536 37568
rect 96600 37504 96616 37568
rect 96680 37504 96688 37568
rect 96368 36480 96688 37504
rect 96368 36416 96376 36480
rect 96440 36416 96456 36480
rect 96520 36416 96536 36480
rect 96600 36416 96616 36480
rect 96680 36416 96688 36480
rect 96368 35392 96688 36416
rect 96368 35328 96376 35392
rect 96440 35328 96456 35392
rect 96520 35328 96536 35392
rect 96600 35328 96616 35392
rect 96680 35328 96688 35392
rect 96368 34304 96688 35328
rect 96368 34240 96376 34304
rect 96440 34240 96456 34304
rect 96520 34240 96536 34304
rect 96600 34240 96616 34304
rect 96680 34240 96688 34304
rect 96368 33216 96688 34240
rect 96368 33152 96376 33216
rect 96440 33152 96456 33216
rect 96520 33152 96536 33216
rect 96600 33152 96616 33216
rect 96680 33152 96688 33216
rect 96368 32128 96688 33152
rect 96368 32064 96376 32128
rect 96440 32064 96456 32128
rect 96520 32064 96536 32128
rect 96600 32064 96616 32128
rect 96680 32064 96688 32128
rect 96368 31040 96688 32064
rect 96368 30976 96376 31040
rect 96440 30976 96456 31040
rect 96520 30976 96536 31040
rect 96600 30976 96616 31040
rect 96680 30976 96688 31040
rect 96368 29952 96688 30976
rect 96368 29888 96376 29952
rect 96440 29888 96456 29952
rect 96520 29888 96536 29952
rect 96600 29888 96616 29952
rect 96680 29888 96688 29952
rect 96368 28864 96688 29888
rect 96368 28800 96376 28864
rect 96440 28800 96456 28864
rect 96520 28800 96536 28864
rect 96600 28800 96616 28864
rect 96680 28800 96688 28864
rect 96368 27776 96688 28800
rect 96368 27712 96376 27776
rect 96440 27712 96456 27776
rect 96520 27712 96536 27776
rect 96600 27712 96616 27776
rect 96680 27712 96688 27776
rect 96368 26688 96688 27712
rect 96368 26624 96376 26688
rect 96440 26624 96456 26688
rect 96520 26624 96536 26688
rect 96600 26624 96616 26688
rect 96680 26624 96688 26688
rect 96368 25600 96688 26624
rect 96368 25536 96376 25600
rect 96440 25536 96456 25600
rect 96520 25536 96536 25600
rect 96600 25536 96616 25600
rect 96680 25536 96688 25600
rect 96368 24512 96688 25536
rect 96368 24448 96376 24512
rect 96440 24448 96456 24512
rect 96520 24448 96536 24512
rect 96600 24448 96616 24512
rect 96680 24448 96688 24512
rect 96368 23424 96688 24448
rect 96368 23360 96376 23424
rect 96440 23360 96456 23424
rect 96520 23360 96536 23424
rect 96600 23360 96616 23424
rect 96680 23360 96688 23424
rect 96368 22336 96688 23360
rect 96368 22272 96376 22336
rect 96440 22272 96456 22336
rect 96520 22272 96536 22336
rect 96600 22272 96616 22336
rect 96680 22272 96688 22336
rect 96368 21248 96688 22272
rect 96368 21184 96376 21248
rect 96440 21184 96456 21248
rect 96520 21184 96536 21248
rect 96600 21184 96616 21248
rect 96680 21184 96688 21248
rect 96368 20160 96688 21184
rect 96368 20096 96376 20160
rect 96440 20096 96456 20160
rect 96520 20096 96536 20160
rect 96600 20096 96616 20160
rect 96680 20096 96688 20160
rect 96368 19072 96688 20096
rect 96368 19008 96376 19072
rect 96440 19008 96456 19072
rect 96520 19008 96536 19072
rect 96600 19008 96616 19072
rect 96680 19008 96688 19072
rect 96368 17984 96688 19008
rect 96368 17920 96376 17984
rect 96440 17920 96456 17984
rect 96520 17920 96536 17984
rect 96600 17920 96616 17984
rect 96680 17920 96688 17984
rect 96368 16896 96688 17920
rect 96368 16832 96376 16896
rect 96440 16832 96456 16896
rect 96520 16832 96536 16896
rect 96600 16832 96616 16896
rect 96680 16832 96688 16896
rect 96368 15808 96688 16832
rect 96368 15744 96376 15808
rect 96440 15744 96456 15808
rect 96520 15744 96536 15808
rect 96600 15744 96616 15808
rect 96680 15744 96688 15808
rect 96368 14720 96688 15744
rect 96368 14656 96376 14720
rect 96440 14656 96456 14720
rect 96520 14656 96536 14720
rect 96600 14656 96616 14720
rect 96680 14656 96688 14720
rect 96368 13632 96688 14656
rect 96368 13568 96376 13632
rect 96440 13568 96456 13632
rect 96520 13568 96536 13632
rect 96600 13568 96616 13632
rect 96680 13568 96688 13632
rect 96368 12544 96688 13568
rect 96368 12480 96376 12544
rect 96440 12480 96456 12544
rect 96520 12480 96536 12544
rect 96600 12480 96616 12544
rect 96680 12480 96688 12544
rect 96368 11456 96688 12480
rect 96368 11392 96376 11456
rect 96440 11392 96456 11456
rect 96520 11392 96536 11456
rect 96600 11392 96616 11456
rect 96680 11392 96688 11456
rect 96368 10368 96688 11392
rect 96368 10304 96376 10368
rect 96440 10304 96456 10368
rect 96520 10304 96536 10368
rect 96600 10304 96616 10368
rect 96680 10304 96688 10368
rect 96368 9280 96688 10304
rect 96368 9216 96376 9280
rect 96440 9216 96456 9280
rect 96520 9216 96536 9280
rect 96600 9216 96616 9280
rect 96680 9216 96688 9280
rect 96368 8192 96688 9216
rect 96368 8128 96376 8192
rect 96440 8128 96456 8192
rect 96520 8128 96536 8192
rect 96600 8128 96616 8192
rect 96680 8128 96688 8192
rect 96368 7104 96688 8128
rect 96368 7040 96376 7104
rect 96440 7040 96456 7104
rect 96520 7040 96536 7104
rect 96600 7040 96616 7104
rect 96680 7040 96688 7104
rect 96368 6016 96688 7040
rect 96368 5952 96376 6016
rect 96440 5952 96456 6016
rect 96520 5952 96536 6016
rect 96600 5952 96616 6016
rect 96680 5952 96688 6016
rect 96368 4928 96688 5952
rect 96368 4864 96376 4928
rect 96440 4864 96456 4928
rect 96520 4864 96536 4928
rect 96600 4864 96616 4928
rect 96680 4864 96688 4928
rect 96368 3840 96688 4864
rect 96368 3776 96376 3840
rect 96440 3776 96456 3840
rect 96520 3776 96536 3840
rect 96600 3776 96616 3840
rect 96680 3776 96688 3840
rect 96368 2752 96688 3776
rect 96368 2688 96376 2752
rect 96440 2688 96456 2752
rect 96520 2688 96536 2752
rect 96600 2688 96616 2752
rect 96680 2688 96688 2752
rect 96368 2128 96688 2688
rect 111728 37024 112048 37584
rect 111728 36960 111736 37024
rect 111800 36960 111816 37024
rect 111880 36960 111896 37024
rect 111960 36960 111976 37024
rect 112040 36960 112048 37024
rect 111728 35936 112048 36960
rect 111728 35872 111736 35936
rect 111800 35872 111816 35936
rect 111880 35872 111896 35936
rect 111960 35872 111976 35936
rect 112040 35872 112048 35936
rect 111728 34848 112048 35872
rect 111728 34784 111736 34848
rect 111800 34784 111816 34848
rect 111880 34784 111896 34848
rect 111960 34784 111976 34848
rect 112040 34784 112048 34848
rect 111728 33760 112048 34784
rect 111728 33696 111736 33760
rect 111800 33696 111816 33760
rect 111880 33696 111896 33760
rect 111960 33696 111976 33760
rect 112040 33696 112048 33760
rect 111728 32672 112048 33696
rect 111728 32608 111736 32672
rect 111800 32608 111816 32672
rect 111880 32608 111896 32672
rect 111960 32608 111976 32672
rect 112040 32608 112048 32672
rect 111728 31584 112048 32608
rect 111728 31520 111736 31584
rect 111800 31520 111816 31584
rect 111880 31520 111896 31584
rect 111960 31520 111976 31584
rect 112040 31520 112048 31584
rect 111728 30496 112048 31520
rect 111728 30432 111736 30496
rect 111800 30432 111816 30496
rect 111880 30432 111896 30496
rect 111960 30432 111976 30496
rect 112040 30432 112048 30496
rect 111728 29408 112048 30432
rect 111728 29344 111736 29408
rect 111800 29344 111816 29408
rect 111880 29344 111896 29408
rect 111960 29344 111976 29408
rect 112040 29344 112048 29408
rect 111728 28320 112048 29344
rect 111728 28256 111736 28320
rect 111800 28256 111816 28320
rect 111880 28256 111896 28320
rect 111960 28256 111976 28320
rect 112040 28256 112048 28320
rect 111728 27232 112048 28256
rect 111728 27168 111736 27232
rect 111800 27168 111816 27232
rect 111880 27168 111896 27232
rect 111960 27168 111976 27232
rect 112040 27168 112048 27232
rect 111728 26144 112048 27168
rect 111728 26080 111736 26144
rect 111800 26080 111816 26144
rect 111880 26080 111896 26144
rect 111960 26080 111976 26144
rect 112040 26080 112048 26144
rect 111728 25056 112048 26080
rect 111728 24992 111736 25056
rect 111800 24992 111816 25056
rect 111880 24992 111896 25056
rect 111960 24992 111976 25056
rect 112040 24992 112048 25056
rect 111728 23968 112048 24992
rect 111728 23904 111736 23968
rect 111800 23904 111816 23968
rect 111880 23904 111896 23968
rect 111960 23904 111976 23968
rect 112040 23904 112048 23968
rect 111728 22880 112048 23904
rect 111728 22816 111736 22880
rect 111800 22816 111816 22880
rect 111880 22816 111896 22880
rect 111960 22816 111976 22880
rect 112040 22816 112048 22880
rect 111728 21792 112048 22816
rect 111728 21728 111736 21792
rect 111800 21728 111816 21792
rect 111880 21728 111896 21792
rect 111960 21728 111976 21792
rect 112040 21728 112048 21792
rect 111728 20704 112048 21728
rect 111728 20640 111736 20704
rect 111800 20640 111816 20704
rect 111880 20640 111896 20704
rect 111960 20640 111976 20704
rect 112040 20640 112048 20704
rect 111728 19616 112048 20640
rect 111728 19552 111736 19616
rect 111800 19552 111816 19616
rect 111880 19552 111896 19616
rect 111960 19552 111976 19616
rect 112040 19552 112048 19616
rect 111728 18528 112048 19552
rect 111728 18464 111736 18528
rect 111800 18464 111816 18528
rect 111880 18464 111896 18528
rect 111960 18464 111976 18528
rect 112040 18464 112048 18528
rect 111728 17440 112048 18464
rect 111728 17376 111736 17440
rect 111800 17376 111816 17440
rect 111880 17376 111896 17440
rect 111960 17376 111976 17440
rect 112040 17376 112048 17440
rect 111728 16352 112048 17376
rect 111728 16288 111736 16352
rect 111800 16288 111816 16352
rect 111880 16288 111896 16352
rect 111960 16288 111976 16352
rect 112040 16288 112048 16352
rect 111728 15264 112048 16288
rect 111728 15200 111736 15264
rect 111800 15200 111816 15264
rect 111880 15200 111896 15264
rect 111960 15200 111976 15264
rect 112040 15200 112048 15264
rect 111728 14176 112048 15200
rect 111728 14112 111736 14176
rect 111800 14112 111816 14176
rect 111880 14112 111896 14176
rect 111960 14112 111976 14176
rect 112040 14112 112048 14176
rect 111728 13088 112048 14112
rect 111728 13024 111736 13088
rect 111800 13024 111816 13088
rect 111880 13024 111896 13088
rect 111960 13024 111976 13088
rect 112040 13024 112048 13088
rect 111728 12000 112048 13024
rect 111728 11936 111736 12000
rect 111800 11936 111816 12000
rect 111880 11936 111896 12000
rect 111960 11936 111976 12000
rect 112040 11936 112048 12000
rect 111728 10912 112048 11936
rect 111728 10848 111736 10912
rect 111800 10848 111816 10912
rect 111880 10848 111896 10912
rect 111960 10848 111976 10912
rect 112040 10848 112048 10912
rect 111728 9824 112048 10848
rect 111728 9760 111736 9824
rect 111800 9760 111816 9824
rect 111880 9760 111896 9824
rect 111960 9760 111976 9824
rect 112040 9760 112048 9824
rect 111728 8736 112048 9760
rect 111728 8672 111736 8736
rect 111800 8672 111816 8736
rect 111880 8672 111896 8736
rect 111960 8672 111976 8736
rect 112040 8672 112048 8736
rect 111728 7648 112048 8672
rect 111728 7584 111736 7648
rect 111800 7584 111816 7648
rect 111880 7584 111896 7648
rect 111960 7584 111976 7648
rect 112040 7584 112048 7648
rect 111728 6560 112048 7584
rect 111728 6496 111736 6560
rect 111800 6496 111816 6560
rect 111880 6496 111896 6560
rect 111960 6496 111976 6560
rect 112040 6496 112048 6560
rect 111728 5472 112048 6496
rect 111728 5408 111736 5472
rect 111800 5408 111816 5472
rect 111880 5408 111896 5472
rect 111960 5408 111976 5472
rect 112040 5408 112048 5472
rect 111728 4384 112048 5408
rect 111728 4320 111736 4384
rect 111800 4320 111816 4384
rect 111880 4320 111896 4384
rect 111960 4320 111976 4384
rect 112040 4320 112048 4384
rect 111728 3296 112048 4320
rect 111728 3232 111736 3296
rect 111800 3232 111816 3296
rect 111880 3232 111896 3296
rect 111960 3232 111976 3296
rect 112040 3232 112048 3296
rect 111728 2208 112048 3232
rect 111728 2144 111736 2208
rect 111800 2144 111816 2208
rect 111880 2144 111896 2208
rect 111960 2144 111976 2208
rect 112040 2144 112048 2208
rect 111728 2128 112048 2144
rect 127088 37568 127408 37584
rect 127088 37504 127096 37568
rect 127160 37504 127176 37568
rect 127240 37504 127256 37568
rect 127320 37504 127336 37568
rect 127400 37504 127408 37568
rect 127088 36480 127408 37504
rect 127088 36416 127096 36480
rect 127160 36416 127176 36480
rect 127240 36416 127256 36480
rect 127320 36416 127336 36480
rect 127400 36416 127408 36480
rect 127088 35392 127408 36416
rect 127088 35328 127096 35392
rect 127160 35328 127176 35392
rect 127240 35328 127256 35392
rect 127320 35328 127336 35392
rect 127400 35328 127408 35392
rect 127088 34304 127408 35328
rect 127088 34240 127096 34304
rect 127160 34240 127176 34304
rect 127240 34240 127256 34304
rect 127320 34240 127336 34304
rect 127400 34240 127408 34304
rect 127088 33216 127408 34240
rect 127088 33152 127096 33216
rect 127160 33152 127176 33216
rect 127240 33152 127256 33216
rect 127320 33152 127336 33216
rect 127400 33152 127408 33216
rect 127088 32128 127408 33152
rect 127088 32064 127096 32128
rect 127160 32064 127176 32128
rect 127240 32064 127256 32128
rect 127320 32064 127336 32128
rect 127400 32064 127408 32128
rect 127088 31040 127408 32064
rect 127088 30976 127096 31040
rect 127160 30976 127176 31040
rect 127240 30976 127256 31040
rect 127320 30976 127336 31040
rect 127400 30976 127408 31040
rect 127088 29952 127408 30976
rect 127088 29888 127096 29952
rect 127160 29888 127176 29952
rect 127240 29888 127256 29952
rect 127320 29888 127336 29952
rect 127400 29888 127408 29952
rect 127088 28864 127408 29888
rect 127088 28800 127096 28864
rect 127160 28800 127176 28864
rect 127240 28800 127256 28864
rect 127320 28800 127336 28864
rect 127400 28800 127408 28864
rect 127088 27776 127408 28800
rect 127088 27712 127096 27776
rect 127160 27712 127176 27776
rect 127240 27712 127256 27776
rect 127320 27712 127336 27776
rect 127400 27712 127408 27776
rect 127088 26688 127408 27712
rect 127088 26624 127096 26688
rect 127160 26624 127176 26688
rect 127240 26624 127256 26688
rect 127320 26624 127336 26688
rect 127400 26624 127408 26688
rect 127088 25600 127408 26624
rect 127088 25536 127096 25600
rect 127160 25536 127176 25600
rect 127240 25536 127256 25600
rect 127320 25536 127336 25600
rect 127400 25536 127408 25600
rect 127088 24512 127408 25536
rect 127088 24448 127096 24512
rect 127160 24448 127176 24512
rect 127240 24448 127256 24512
rect 127320 24448 127336 24512
rect 127400 24448 127408 24512
rect 127088 23424 127408 24448
rect 127088 23360 127096 23424
rect 127160 23360 127176 23424
rect 127240 23360 127256 23424
rect 127320 23360 127336 23424
rect 127400 23360 127408 23424
rect 127088 22336 127408 23360
rect 127088 22272 127096 22336
rect 127160 22272 127176 22336
rect 127240 22272 127256 22336
rect 127320 22272 127336 22336
rect 127400 22272 127408 22336
rect 127088 21248 127408 22272
rect 127088 21184 127096 21248
rect 127160 21184 127176 21248
rect 127240 21184 127256 21248
rect 127320 21184 127336 21248
rect 127400 21184 127408 21248
rect 127088 20160 127408 21184
rect 127088 20096 127096 20160
rect 127160 20096 127176 20160
rect 127240 20096 127256 20160
rect 127320 20096 127336 20160
rect 127400 20096 127408 20160
rect 127088 19072 127408 20096
rect 127088 19008 127096 19072
rect 127160 19008 127176 19072
rect 127240 19008 127256 19072
rect 127320 19008 127336 19072
rect 127400 19008 127408 19072
rect 127088 17984 127408 19008
rect 127088 17920 127096 17984
rect 127160 17920 127176 17984
rect 127240 17920 127256 17984
rect 127320 17920 127336 17984
rect 127400 17920 127408 17984
rect 127088 16896 127408 17920
rect 127088 16832 127096 16896
rect 127160 16832 127176 16896
rect 127240 16832 127256 16896
rect 127320 16832 127336 16896
rect 127400 16832 127408 16896
rect 127088 15808 127408 16832
rect 127088 15744 127096 15808
rect 127160 15744 127176 15808
rect 127240 15744 127256 15808
rect 127320 15744 127336 15808
rect 127400 15744 127408 15808
rect 127088 14720 127408 15744
rect 127088 14656 127096 14720
rect 127160 14656 127176 14720
rect 127240 14656 127256 14720
rect 127320 14656 127336 14720
rect 127400 14656 127408 14720
rect 127088 13632 127408 14656
rect 127088 13568 127096 13632
rect 127160 13568 127176 13632
rect 127240 13568 127256 13632
rect 127320 13568 127336 13632
rect 127400 13568 127408 13632
rect 127088 12544 127408 13568
rect 127088 12480 127096 12544
rect 127160 12480 127176 12544
rect 127240 12480 127256 12544
rect 127320 12480 127336 12544
rect 127400 12480 127408 12544
rect 127088 11456 127408 12480
rect 127088 11392 127096 11456
rect 127160 11392 127176 11456
rect 127240 11392 127256 11456
rect 127320 11392 127336 11456
rect 127400 11392 127408 11456
rect 127088 10368 127408 11392
rect 127088 10304 127096 10368
rect 127160 10304 127176 10368
rect 127240 10304 127256 10368
rect 127320 10304 127336 10368
rect 127400 10304 127408 10368
rect 127088 9280 127408 10304
rect 127088 9216 127096 9280
rect 127160 9216 127176 9280
rect 127240 9216 127256 9280
rect 127320 9216 127336 9280
rect 127400 9216 127408 9280
rect 127088 8192 127408 9216
rect 127088 8128 127096 8192
rect 127160 8128 127176 8192
rect 127240 8128 127256 8192
rect 127320 8128 127336 8192
rect 127400 8128 127408 8192
rect 127088 7104 127408 8128
rect 127088 7040 127096 7104
rect 127160 7040 127176 7104
rect 127240 7040 127256 7104
rect 127320 7040 127336 7104
rect 127400 7040 127408 7104
rect 127088 6016 127408 7040
rect 127088 5952 127096 6016
rect 127160 5952 127176 6016
rect 127240 5952 127256 6016
rect 127320 5952 127336 6016
rect 127400 5952 127408 6016
rect 127088 4928 127408 5952
rect 127088 4864 127096 4928
rect 127160 4864 127176 4928
rect 127240 4864 127256 4928
rect 127320 4864 127336 4928
rect 127400 4864 127408 4928
rect 127088 3840 127408 4864
rect 127088 3776 127096 3840
rect 127160 3776 127176 3840
rect 127240 3776 127256 3840
rect 127320 3776 127336 3840
rect 127400 3776 127408 3840
rect 127088 2752 127408 3776
rect 127088 2688 127096 2752
rect 127160 2688 127176 2752
rect 127240 2688 127256 2752
rect 127320 2688 127336 2752
rect 127400 2688 127408 2752
rect 127088 2128 127408 2688
rect 142448 37024 142768 37584
rect 142448 36960 142456 37024
rect 142520 36960 142536 37024
rect 142600 36960 142616 37024
rect 142680 36960 142696 37024
rect 142760 36960 142768 37024
rect 142448 35936 142768 36960
rect 142448 35872 142456 35936
rect 142520 35872 142536 35936
rect 142600 35872 142616 35936
rect 142680 35872 142696 35936
rect 142760 35872 142768 35936
rect 142448 34848 142768 35872
rect 142448 34784 142456 34848
rect 142520 34784 142536 34848
rect 142600 34784 142616 34848
rect 142680 34784 142696 34848
rect 142760 34784 142768 34848
rect 142448 33760 142768 34784
rect 142448 33696 142456 33760
rect 142520 33696 142536 33760
rect 142600 33696 142616 33760
rect 142680 33696 142696 33760
rect 142760 33696 142768 33760
rect 142448 32672 142768 33696
rect 142448 32608 142456 32672
rect 142520 32608 142536 32672
rect 142600 32608 142616 32672
rect 142680 32608 142696 32672
rect 142760 32608 142768 32672
rect 142448 31584 142768 32608
rect 142448 31520 142456 31584
rect 142520 31520 142536 31584
rect 142600 31520 142616 31584
rect 142680 31520 142696 31584
rect 142760 31520 142768 31584
rect 142448 30496 142768 31520
rect 142448 30432 142456 30496
rect 142520 30432 142536 30496
rect 142600 30432 142616 30496
rect 142680 30432 142696 30496
rect 142760 30432 142768 30496
rect 142448 29408 142768 30432
rect 142448 29344 142456 29408
rect 142520 29344 142536 29408
rect 142600 29344 142616 29408
rect 142680 29344 142696 29408
rect 142760 29344 142768 29408
rect 142448 28320 142768 29344
rect 142448 28256 142456 28320
rect 142520 28256 142536 28320
rect 142600 28256 142616 28320
rect 142680 28256 142696 28320
rect 142760 28256 142768 28320
rect 142448 27232 142768 28256
rect 142448 27168 142456 27232
rect 142520 27168 142536 27232
rect 142600 27168 142616 27232
rect 142680 27168 142696 27232
rect 142760 27168 142768 27232
rect 142448 26144 142768 27168
rect 142448 26080 142456 26144
rect 142520 26080 142536 26144
rect 142600 26080 142616 26144
rect 142680 26080 142696 26144
rect 142760 26080 142768 26144
rect 142448 25056 142768 26080
rect 142448 24992 142456 25056
rect 142520 24992 142536 25056
rect 142600 24992 142616 25056
rect 142680 24992 142696 25056
rect 142760 24992 142768 25056
rect 142448 23968 142768 24992
rect 142448 23904 142456 23968
rect 142520 23904 142536 23968
rect 142600 23904 142616 23968
rect 142680 23904 142696 23968
rect 142760 23904 142768 23968
rect 142448 22880 142768 23904
rect 142448 22816 142456 22880
rect 142520 22816 142536 22880
rect 142600 22816 142616 22880
rect 142680 22816 142696 22880
rect 142760 22816 142768 22880
rect 142448 21792 142768 22816
rect 142448 21728 142456 21792
rect 142520 21728 142536 21792
rect 142600 21728 142616 21792
rect 142680 21728 142696 21792
rect 142760 21728 142768 21792
rect 142448 20704 142768 21728
rect 142448 20640 142456 20704
rect 142520 20640 142536 20704
rect 142600 20640 142616 20704
rect 142680 20640 142696 20704
rect 142760 20640 142768 20704
rect 142448 19616 142768 20640
rect 142448 19552 142456 19616
rect 142520 19552 142536 19616
rect 142600 19552 142616 19616
rect 142680 19552 142696 19616
rect 142760 19552 142768 19616
rect 142448 18528 142768 19552
rect 142448 18464 142456 18528
rect 142520 18464 142536 18528
rect 142600 18464 142616 18528
rect 142680 18464 142696 18528
rect 142760 18464 142768 18528
rect 142448 17440 142768 18464
rect 142448 17376 142456 17440
rect 142520 17376 142536 17440
rect 142600 17376 142616 17440
rect 142680 17376 142696 17440
rect 142760 17376 142768 17440
rect 142448 16352 142768 17376
rect 142448 16288 142456 16352
rect 142520 16288 142536 16352
rect 142600 16288 142616 16352
rect 142680 16288 142696 16352
rect 142760 16288 142768 16352
rect 142448 15264 142768 16288
rect 142448 15200 142456 15264
rect 142520 15200 142536 15264
rect 142600 15200 142616 15264
rect 142680 15200 142696 15264
rect 142760 15200 142768 15264
rect 142448 14176 142768 15200
rect 142448 14112 142456 14176
rect 142520 14112 142536 14176
rect 142600 14112 142616 14176
rect 142680 14112 142696 14176
rect 142760 14112 142768 14176
rect 142448 13088 142768 14112
rect 142448 13024 142456 13088
rect 142520 13024 142536 13088
rect 142600 13024 142616 13088
rect 142680 13024 142696 13088
rect 142760 13024 142768 13088
rect 142448 12000 142768 13024
rect 142448 11936 142456 12000
rect 142520 11936 142536 12000
rect 142600 11936 142616 12000
rect 142680 11936 142696 12000
rect 142760 11936 142768 12000
rect 142448 10912 142768 11936
rect 142448 10848 142456 10912
rect 142520 10848 142536 10912
rect 142600 10848 142616 10912
rect 142680 10848 142696 10912
rect 142760 10848 142768 10912
rect 142448 9824 142768 10848
rect 142448 9760 142456 9824
rect 142520 9760 142536 9824
rect 142600 9760 142616 9824
rect 142680 9760 142696 9824
rect 142760 9760 142768 9824
rect 142448 8736 142768 9760
rect 142448 8672 142456 8736
rect 142520 8672 142536 8736
rect 142600 8672 142616 8736
rect 142680 8672 142696 8736
rect 142760 8672 142768 8736
rect 142448 7648 142768 8672
rect 142448 7584 142456 7648
rect 142520 7584 142536 7648
rect 142600 7584 142616 7648
rect 142680 7584 142696 7648
rect 142760 7584 142768 7648
rect 142448 6560 142768 7584
rect 142448 6496 142456 6560
rect 142520 6496 142536 6560
rect 142600 6496 142616 6560
rect 142680 6496 142696 6560
rect 142760 6496 142768 6560
rect 142448 5472 142768 6496
rect 142448 5408 142456 5472
rect 142520 5408 142536 5472
rect 142600 5408 142616 5472
rect 142680 5408 142696 5472
rect 142760 5408 142768 5472
rect 142448 4384 142768 5408
rect 142448 4320 142456 4384
rect 142520 4320 142536 4384
rect 142600 4320 142616 4384
rect 142680 4320 142696 4384
rect 142760 4320 142768 4384
rect 142448 3296 142768 4320
rect 142448 3232 142456 3296
rect 142520 3232 142536 3296
rect 142600 3232 142616 3296
rect 142680 3232 142696 3296
rect 142760 3232 142768 3296
rect 142448 2208 142768 3232
rect 142448 2144 142456 2208
rect 142520 2144 142536 2208
rect 142600 2144 142616 2208
rect 142680 2144 142696 2208
rect 142760 2144 142768 2208
rect 142448 2128 142768 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 61732 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A1
timestamp 1666464484
transform -1 0 77832 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__S
timestamp 1666464484
transform 1 0 77096 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__A
timestamp 1666464484
transform -1 0 63664 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__A0
timestamp 1666464484
transform -1 0 76268 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__A1
timestamp 1666464484
transform 1 0 75624 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__S
timestamp 1666464484
transform 1 0 74612 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A1
timestamp 1666464484
transform -1 0 80224 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__S
timestamp 1666464484
transform 1 0 78844 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A0
timestamp 1666464484
transform -1 0 77740 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A1
timestamp 1666464484
transform 1 0 78108 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__S
timestamp 1666464484
transform 1 0 77096 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A1
timestamp 1666464484
transform -1 0 83168 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__S
timestamp 1666464484
transform -1 0 81420 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A0
timestamp 1666464484
transform 1 0 84456 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A1
timestamp 1666464484
transform -1 0 84364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__S
timestamp 1666464484
transform -1 0 85192 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__A1
timestamp 1666464484
transform -1 0 82432 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__S
timestamp 1666464484
transform 1 0 81696 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A0
timestamp 1666464484
transform -1 0 82616 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A1
timestamp 1666464484
transform -1 0 83996 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__S
timestamp 1666464484
transform -1 0 83168 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__A1
timestamp 1666464484
transform -1 0 84824 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__S
timestamp 1666464484
transform -1 0 82524 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__161__A0
timestamp 1666464484
transform 1 0 82616 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__161__A1
timestamp 1666464484
transform -1 0 83260 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__161__S
timestamp 1666464484
transform 1 0 83168 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__A1
timestamp 1666464484
transform -1 0 83720 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__S
timestamp 1666464484
transform -1 0 81972 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__164__A0
timestamp 1666464484
transform -1 0 83812 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__164__A1
timestamp 1666464484
transform -1 0 84916 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__164__S
timestamp 1666464484
transform 1 0 83628 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__166__A1
timestamp 1666464484
transform -1 0 80776 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__166__S
timestamp 1666464484
transform -1 0 79672 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__167__A0
timestamp 1666464484
transform -1 0 80776 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__167__A1
timestamp 1666464484
transform -1 0 80224 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__167__S
timestamp 1666464484
transform 1 0 78660 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__A1
timestamp 1666464484
transform -1 0 71760 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__S
timestamp 1666464484
transform 1 0 70932 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__A0
timestamp 1666464484
transform -1 0 72312 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__A1
timestamp 1666464484
transform -1 0 71944 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__S
timestamp 1666464484
transform 1 0 70932 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__172__A
timestamp 1666464484
transform 1 0 61456 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__173__A1
timestamp 1666464484
transform -1 0 69368 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A0
timestamp 1666464484
transform -1 0 70288 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A1
timestamp 1666464484
transform 1 0 68908 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__S
timestamp 1666464484
transform 1 0 68632 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__A1
timestamp 1666464484
transform -1 0 67344 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__A0
timestamp 1666464484
transform -1 0 67896 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__A1
timestamp 1666464484
transform 1 0 67528 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__S
timestamp 1666464484
transform 1 0 67160 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__179__A1
timestamp 1666464484
transform -1 0 65320 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__A
timestamp 1666464484
transform -1 0 54464 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A0
timestamp 1666464484
transform -1 0 65504 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A1
timestamp 1666464484
transform -1 0 66056 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__183__A1
timestamp 1666464484
transform -1 0 66056 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A0
timestamp 1666464484
transform -1 0 64952 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A1
timestamp 1666464484
transform -1 0 65964 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__A1
timestamp 1666464484
transform -1 0 58236 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__187__A0
timestamp 1666464484
transform -1 0 58604 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__187__A1
timestamp 1666464484
transform 1 0 57868 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__A1
timestamp 1666464484
transform -1 0 55660 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A0
timestamp 1666464484
transform -1 0 56672 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A1
timestamp 1666464484
transform -1 0 56028 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__A1
timestamp 1666464484
transform -1 0 59064 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A0
timestamp 1666464484
transform -1 0 59248 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A1
timestamp 1666464484
transform -1 0 59156 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__A1
timestamp 1666464484
transform -1 0 61088 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__A0
timestamp 1666464484
transform -1 0 61824 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__A1
timestamp 1666464484
transform -1 0 61272 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__198__A0
timestamp 1666464484
transform -1 0 62192 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__198__A1
timestamp 1666464484
transform -1 0 64400 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__A1
timestamp 1666464484
transform -1 0 64216 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__201__A0
timestamp 1666464484
transform -1 0 63848 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__201__A1
timestamp 1666464484
transform -1 0 64400 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__202__A1
timestamp 1666464484
transform 1 0 63664 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__204__A
timestamp 1666464484
transform 1 0 37168 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__A1
timestamp 1666464484
transform -1 0 51612 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__S
timestamp 1666464484
transform 1 0 51152 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__206__A0
timestamp 1666464484
transform -1 0 53084 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__206__A1
timestamp 1666464484
transform -1 0 53636 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__208__A1
timestamp 1666464484
transform -1 0 53912 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__208__S
timestamp 1666464484
transform 1 0 50324 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__209__A1
timestamp 1666464484
transform -1 0 53912 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__A1
timestamp 1666464484
transform -1 0 48760 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__S
timestamp 1666464484
transform 1 0 47104 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A
timestamp 1666464484
transform 1 0 29532 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__A0
timestamp 1666464484
transform -1 0 48208 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__A1
timestamp 1666464484
transform -1 0 49680 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__S
timestamp 1666464484
transform 1 0 46460 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__A1
timestamp 1666464484
transform -1 0 48208 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__S
timestamp 1666464484
transform -1 0 47840 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A1
timestamp 1666464484
transform -1 0 49128 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__S
timestamp 1666464484
transform -1 0 47288 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__A1
timestamp 1666464484
transform -1 0 43608 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__S
timestamp 1666464484
transform 1 0 41952 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__A1
timestamp 1666464484
transform -1 0 41400 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__S
timestamp 1666464484
transform 1 0 41124 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__221__A1
timestamp 1666464484
transform -1 0 43884 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__221__S
timestamp 1666464484
transform -1 0 42872 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__A1
timestamp 1666464484
transform 1 0 43424 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__S
timestamp 1666464484
transform 1 0 43148 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__A1
timestamp 1666464484
transform -1 0 41768 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__S
timestamp 1666464484
transform -1 0 40756 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__A1
timestamp 1666464484
transform 1 0 40572 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__S
timestamp 1666464484
transform 1 0 39376 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__A1
timestamp 1666464484
transform -1 0 38824 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__S
timestamp 1666464484
transform -1 0 38916 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__A1
timestamp 1666464484
transform -1 0 38456 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__S
timestamp 1666464484
transform 1 0 36708 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__A1
timestamp 1666464484
transform -1 0 37720 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__S
timestamp 1666464484
transform 1 0 36248 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__A1
timestamp 1666464484
transform 1 0 36064 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__S
timestamp 1666464484
transform 1 0 34224 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__233__A1
timestamp 1666464484
transform -1 0 36156 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__233__S
timestamp 1666464484
transform -1 0 35328 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__A1
timestamp 1666464484
transform -1 0 32476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__S
timestamp 1666464484
transform 1 0 33580 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A1
timestamp 1666464484
transform -1 0 28704 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__S
timestamp 1666464484
transform 1 0 28612 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__A1
timestamp 1666464484
transform -1 0 28520 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__S
timestamp 1666464484
transform -1 0 27692 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A1
timestamp 1666464484
transform -1 0 28796 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__S
timestamp 1666464484
transform 1 0 29072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A1
timestamp 1666464484
transform -1 0 29164 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__S
timestamp 1666464484
transform 1 0 29716 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__A1
timestamp 1666464484
transform -1 0 24932 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__S
timestamp 1666464484
transform 1 0 24656 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A1
timestamp 1666464484
transform -1 0 24748 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__S
timestamp 1666464484
transform 1 0 24012 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__A0
timestamp 1666464484
transform -1 0 22908 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__A1
timestamp 1666464484
transform -1 0 24104 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__S
timestamp 1666464484
transform 1 0 25944 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__A1
timestamp 1666464484
transform 1 0 23920 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__S
timestamp 1666464484
transform -1 0 22724 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__A_N
timestamp 1666464484
transform 1 0 4600 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A
timestamp 1666464484
transform 1 0 74060 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__B_N
timestamp 1666464484
transform 1 0 75164 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__A
timestamp 1666464484
transform 1 0 61180 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__B
timestamp 1666464484
transform -1 0 59432 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__A
timestamp 1666464484
transform 1 0 32660 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__A
timestamp 1666464484
transform 1 0 20884 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__A
timestamp 1666464484
transform -1 0 20884 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__A
timestamp 1666464484
transform 1 0 26496 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__A
timestamp 1666464484
transform 1 0 28428 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__A
timestamp 1666464484
transform 1 0 32660 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__A
timestamp 1666464484
transform -1 0 35420 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__A
timestamp 1666464484
transform -1 0 38180 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A
timestamp 1666464484
transform -1 0 40204 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__A
timestamp 1666464484
transform 1 0 44988 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__266__A
timestamp 1666464484
transform -1 0 42044 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__A
timestamp 1666464484
transform -1 0 49312 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__A
timestamp 1666464484
transform 1 0 66056 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__A
timestamp 1666464484
transform 1 0 66608 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__A
timestamp 1666464484
transform 1 0 66976 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__A
timestamp 1666464484
transform 1 0 68080 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__282__A
timestamp 1666464484
transform -1 0 69552 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__A
timestamp 1666464484
transform 1 0 69552 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__A
timestamp 1666464484
transform 1 0 78752 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__A
timestamp 1666464484
transform 1 0 85284 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__A
timestamp 1666464484
transform 1 0 82524 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__A
timestamp 1666464484
transform 1 0 81880 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__A
timestamp 1666464484
transform -1 0 86296 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__A
timestamp 1666464484
transform 1 0 74888 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__A
timestamp 1666464484
transform 1 0 73508 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__A
timestamp 1666464484
transform -1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__A
timestamp 1666464484
transform 1 0 30176 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__A
timestamp 1666464484
transform 1 0 8464 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__CLK
timestamp 1666464484
transform 1 0 23828 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__CLK
timestamp 1666464484
transform 1 0 24564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__CLK
timestamp 1666464484
transform 1 0 28980 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__297__CLK
timestamp 1666464484
transform 1 0 28060 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__298__CLK
timestamp 1666464484
transform 1 0 32384 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__299__CLK
timestamp 1666464484
transform -1 0 36892 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__300__CLK
timestamp 1666464484
transform -1 0 37628 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__301__CLK
timestamp 1666464484
transform 1 0 38732 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__302__CLK
timestamp 1666464484
transform -1 0 42780 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__303__CLK
timestamp 1666464484
transform 1 0 41308 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__304__CLK
timestamp 1666464484
transform 1 0 50324 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__305__CLK
timestamp 1666464484
transform 1 0 45264 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__306__CLK
timestamp 1666464484
transform 1 0 50324 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__CLK
timestamp 1666464484
transform 1 0 50324 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__308__CLK
timestamp 1666464484
transform -1 0 62744 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__309__CLK
timestamp 1666464484
transform -1 0 60904 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__310__CLK
timestamp 1666464484
transform 1 0 58604 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__CLK
timestamp 1666464484
transform 1 0 58604 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__CLK
timestamp 1666464484
transform 1 0 54004 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__CLK
timestamp 1666464484
transform 1 0 54556 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__314__CLK
timestamp 1666464484
transform -1 0 66608 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__315__CLK
timestamp 1666464484
transform -1 0 65228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__316__CLK
timestamp 1666464484
transform 1 0 69184 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__CLK
timestamp 1666464484
transform -1 0 70840 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__318__CLK
timestamp 1666464484
transform 1 0 71484 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__319__CLK
timestamp 1666464484
transform 1 0 76544 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__320__CLK
timestamp 1666464484
transform -1 0 85744 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__321__CLK
timestamp 1666464484
transform -1 0 79120 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__322__CLK
timestamp 1666464484
transform 1 0 78016 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__323__CLK
timestamp 1666464484
transform -1 0 79672 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__324__CLK
timestamp 1666464484
transform 1 0 76452 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__325__CLK
timestamp 1666464484
transform 1 0 73508 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__326__CLK
timestamp 1666464484
transform 1 0 6256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__326__D
timestamp 1666464484
transform -1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__327__CLK
timestamp 1666464484
transform 1 0 31832 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__327__D
timestamp 1666464484
transform -1 0 30452 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__328__CLK
timestamp 1666464484
transform 1 0 9108 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__331__A
timestamp 1666464484
transform -1 0 20792 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__332__A
timestamp 1666464484
transform 1 0 26496 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__A
timestamp 1666464484
transform -1 0 31832 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__A
timestamp 1666464484
transform 1 0 36800 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__A
timestamp 1666464484
transform -1 0 40480 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__336__A
timestamp 1666464484
transform -1 0 42136 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__A
timestamp 1666464484
transform -1 0 48208 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__338__A
timestamp 1666464484
transform -1 0 51060 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__A
timestamp 1666464484
transform -1 0 57040 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__340__A
timestamp 1666464484
transform 1 0 52900 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__A
timestamp 1666464484
transform 1 0 29532 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__A
timestamp 1666464484
transform 1 0 33120 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__A
timestamp 1666464484
transform 1 0 38088 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__344__A
timestamp 1666464484
transform 1 0 41400 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__A
timestamp 1666464484
transform 1 0 45540 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__346__A
timestamp 1666464484
transform 1 0 49864 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__347__A
timestamp 1666464484
transform 1 0 54004 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__A
timestamp 1666464484
transform 1 0 58604 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__A
timestamp 1666464484
transform 1 0 6808 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__A
timestamp 1666464484
transform 1 0 10396 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__351__A
timestamp 1666464484
transform 1 0 24104 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__352__A
timestamp 1666464484
transform 1 0 17940 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__A
timestamp 1666464484
transform -1 0 20240 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__354__A
timestamp 1666464484
transform -1 0 39928 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__A
timestamp 1666464484
transform -1 0 43516 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__356__A
timestamp 1666464484
transform -1 0 46552 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__A
timestamp 1666464484
transform 1 0 51704 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__358__A
timestamp 1666464484
transform 1 0 55936 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__359__A
timestamp 1666464484
transform -1 0 59432 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__360__A
timestamp 1666464484
transform -1 0 63848 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__A
timestamp 1666464484
transform -1 0 69920 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__362__A
timestamp 1666464484
transform -1 0 67712 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__363__A
timestamp 1666464484
transform -1 0 73692 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__A
timestamp 1666464484
transform 1 0 82800 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__365__A
timestamp 1666464484
transform 1 0 85284 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__366__A
timestamp 1666464484
transform -1 0 91172 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__367__A
timestamp 1666464484
transform 1 0 94116 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__368__A
timestamp 1666464484
transform 1 0 97796 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__369__A
timestamp 1666464484
transform 1 0 102212 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__A
timestamp 1666464484
transform 1 0 105708 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__371__A
timestamp 1666464484
transform -1 0 110400 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__372__A
timestamp 1666464484
transform 1 0 114080 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__373__A
timestamp 1666464484
transform 1 0 118588 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__A
timestamp 1666464484
transform 1 0 122636 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__375__A
timestamp 1666464484
transform 1 0 127144 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__376__A
timestamp 1666464484
transform 1 0 130916 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__377__A
timestamp 1666464484
transform 1 0 120980 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__378__A
timestamp 1666464484
transform 1 0 113160 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__379__A
timestamp 1666464484
transform 1 0 106996 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__380__A
timestamp 1666464484
transform 1 0 95312 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__381__A
timestamp 1666464484
transform 1 0 45264 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__382__A
timestamp 1666464484
transform 1 0 20976 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__383__A
timestamp 1666464484
transform -1 0 25944 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A
timestamp 1666464484
transform -1 0 31096 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__385__A
timestamp 1666464484
transform 1 0 35328 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__386__A
timestamp 1666464484
transform 1 0 40848 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__387__A
timestamp 1666464484
transform 1 0 44436 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__388__A
timestamp 1666464484
transform 1 0 48576 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__389__A
timestamp 1666464484
transform 1 0 52992 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__390__A
timestamp 1666464484
transform 1 0 56304 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__391__A
timestamp 1666464484
transform 1 0 60628 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__392__A
timestamp 1666464484
transform -1 0 65320 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__393__A
timestamp 1666464484
transform 1 0 69184 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__A
timestamp 1666464484
transform 1 0 75072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__395__A
timestamp 1666464484
transform 1 0 77832 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__A
timestamp 1666464484
transform -1 0 84548 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__397__A
timestamp 1666464484
transform -1 0 86572 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__A
timestamp 1666464484
transform 1 0 90160 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__399__A
timestamp 1666464484
transform 1 0 94668 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__400__A
timestamp 1666464484
transform 1 0 99268 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__401__A
timestamp 1666464484
transform -1 0 103592 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__402__A
timestamp 1666464484
transform -1 0 107640 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__403__A
timestamp 1666464484
transform -1 0 111596 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__A
timestamp 1666464484
transform -1 0 115828 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__405__A
timestamp 1666464484
transform -1 0 132848 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__406__A
timestamp 1666464484
transform -1 0 124016 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__407__A
timestamp 1666464484
transform -1 0 136620 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__408__A
timestamp 1666464484
transform -1 0 138460 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__A
timestamp 1666464484
transform 1 0 139472 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__410__A
timestamp 1666464484
transform -1 0 142232 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__411__A
timestamp 1666464484
transform -1 0 144440 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__412__A
timestamp 1666464484
transform 1 0 146740 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__413__A
timestamp 1666464484
transform 1 0 8832 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__414__A
timestamp 1666464484
transform -1 0 19688 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__415__A
timestamp 1666464484
transform 1 0 25392 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__416__A
timestamp 1666464484
transform -1 0 18676 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__417__A
timestamp 1666464484
transform 1 0 34224 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__418__A
timestamp 1666464484
transform 1 0 21804 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__419__A
timestamp 1666464484
transform -1 0 25944 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__420__A
timestamp 1666464484
transform 1 0 31096 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_io_wbs_clk_A
timestamp 1666464484
transform 1 0 42596 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1666464484
transform -1 0 7360 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1666464484
transform -1 0 35880 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1666464484
transform -1 0 37720 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1666464484
transform -1 0 39560 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1666464484
transform -1 0 41032 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1666464484
transform -1 0 44068 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1666464484
transform -1 0 45264 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1666464484
transform -1 0 46000 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1666464484
transform -1 0 49312 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1666464484
transform -1 0 50600 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1666464484
transform -1 0 52440 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1666464484
transform -1 0 10120 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1666464484
transform -1 0 54924 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1666464484
transform -1 0 55936 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1666464484
transform -1 0 57592 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1666464484
transform -1 0 60536 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1666464484
transform -1 0 62468 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1666464484
transform -1 0 62744 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1666464484
transform -1 0 66148 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1666464484
transform -1 0 67160 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1666464484
transform -1 0 69828 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1666464484
transform -1 0 70472 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1666464484
transform -1 0 14628 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1666464484
transform -1 0 72312 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1666464484
transform -1 0 74152 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1666464484
transform -1 0 17572 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1666464484
transform -1 0 21160 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1666464484
transform -1 0 23552 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1666464484
transform -1 0 26680 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1666464484
transform -1 0 29900 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1666464484
transform -1 0 31832 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1666464484
transform -1 0 33856 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1666464484
transform -1 0 82616 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1666464484
transform -1 0 108744 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1666464484
transform -1 0 111044 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1666464484
transform -1 0 112884 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1666464484
transform -1 0 114816 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1666464484
transform -1 0 116380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1666464484
transform -1 0 118036 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1666464484
transform -1 0 120060 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1666464484
transform -1 0 121072 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1666464484
transform -1 0 124568 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1666464484
transform -1 0 125764 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1666464484
transform -1 0 85836 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1666464484
transform -1 0 127880 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1666464484
transform -1 0 129076 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1666464484
transform -1 0 131652 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1666464484
transform -1 0 133400 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1666464484
transform -1 0 134320 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1666464484
transform -1 0 136160 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1666464484
transform -1 0 138092 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1666464484
transform -1 0 140668 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1666464484
transform -1 0 142784 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1666464484
transform -1 0 143796 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1666464484
transform -1 0 87676 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1666464484
transform -1 0 145176 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1666464484
transform -1 0 147476 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1666464484
transform -1 0 90896 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1666464484
transform -1 0 94116 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1666464484
transform -1 0 97152 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1666464484
transform -1 0 100004 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1666464484
transform -1 0 103960 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1666464484
transform -1 0 105156 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1666464484
transform -1 0 108192 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1666464484
transform -1 0 58236 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1666464484
transform -1 0 61916 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1666464484
transform -1 0 20332 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1666464484
transform -1 0 25852 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1666464484
transform -1 0 32016 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1666464484
transform -1 0 37444 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1666464484
transform -1 0 40940 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1666464484
transform -1 0 45724 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1666464484
transform -1 0 49128 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1666464484
transform -1 0 53268 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1666464484
transform -1 0 4968 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1666464484
transform -1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1666464484
transform -1 0 60168 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1666464484
transform -1 0 64400 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1666464484
transform -1 0 68540 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1666464484
transform -1 0 73140 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1666464484
transform -1 0 78844 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1666464484
transform -1 0 84548 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1666464484
transform -1 0 87124 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1666464484
transform -1 0 89148 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1666464484
transform -1 0 93656 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1666464484
transform -1 0 97796 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1666464484
transform -1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1666464484
transform -1 0 101936 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1666464484
transform -1 0 105708 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1666464484
transform -1 0 110308 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1666464484
transform -1 0 114264 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1666464484
transform -1 0 118496 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1666464484
transform -1 0 122636 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1666464484
transform -1 0 126408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1666464484
transform -1 0 130916 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1666464484
transform -1 0 134872 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1666464484
transform -1 0 138828 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 1666464484
transform -1 0 25300 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1666464484
transform -1 0 143336 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1666464484
transform -1 0 148396 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1666464484
transform -1 0 30636 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1666464484
transform -1 0 35696 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1666464484
transform -1 0 39560 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1666464484
transform -1 0 43792 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1666464484
transform -1 0 48760 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1666464484
transform -1 0 52900 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 1666464484
transform -1 0 56120 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 1666464484
transform -1 0 7360 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 1666464484
transform -1 0 15180 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 1666464484
transform -1 0 20516 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input111_A
timestamp 1666464484
transform -1 0 26128 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input112_A
timestamp 1666464484
transform -1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input113_A
timestamp 1666464484
transform -1 0 8096 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input114_A
timestamp 1666464484
transform -1 0 10304 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output116_A
timestamp 1666464484
transform -1 0 9292 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output117_A
timestamp 1666464484
transform -1 0 12512 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output118_A
timestamp 1666464484
transform 1 0 16008 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output119_A
timestamp 1666464484
transform -1 0 19964 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output120_A
timestamp 1666464484
transform -1 0 22632 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output121_A
timestamp 1666464484
transform -1 0 25392 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output122_A
timestamp 1666464484
transform -1 0 28152 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output123_A
timestamp 1666464484
transform -1 0 30912 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output124_A
timestamp 1666464484
transform -1 0 77464 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output125_A
timestamp 1666464484
transform -1 0 80592 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output126_A
timestamp 1666464484
transform -1 0 85284 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output127_A
timestamp 1666464484
transform -1 0 89792 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output128_A
timestamp 1666464484
transform -1 0 92276 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output129_A
timestamp 1666464484
transform -1 0 96600 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output130_A
timestamp 1666464484
transform -1 0 98532 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output131_A
timestamp 1666464484
transform -1 0 100740 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output132_A
timestamp 1666464484
transform 1 0 102856 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output134_A
timestamp 1666464484
transform -1 0 34592 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output135_A
timestamp 1666464484
transform -1 0 37168 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output136_A
timestamp 1666464484
transform -1 0 39376 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output137_A
timestamp 1666464484
transform -1 0 39008 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output138_A
timestamp 1666464484
transform -1 0 42872 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output139_A
timestamp 1666464484
transform -1 0 44344 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output140_A
timestamp 1666464484
transform -1 0 46184 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output141_A
timestamp 1666464484
transform -1 0 46736 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output142_A
timestamp 1666464484
transform -1 0 50508 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output143_A
timestamp 1666464484
transform -1 0 51428 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output145_A
timestamp 1666464484
transform 1 0 54096 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output146_A
timestamp 1666464484
transform -1 0 55200 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output147_A
timestamp 1666464484
transform -1 0 54280 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output148_A
timestamp 1666464484
transform -1 0 60076 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output149_A
timestamp 1666464484
transform -1 0 59984 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output150_A
timestamp 1666464484
transform -1 0 63112 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output151_A
timestamp 1666464484
transform -1 0 64952 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output152_A
timestamp 1666464484
transform -1 0 66792 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output153_A
timestamp 1666464484
transform -1 0 68632 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output154_A
timestamp 1666464484
transform -1 0 70472 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output156_A
timestamp 1666464484
transform -1 0 72680 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output157_A
timestamp 1666464484
transform -1 0 73048 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output163_A
timestamp 1666464484
transform -1 0 31832 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output164_A
timestamp 1666464484
transform -1 0 33304 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output165_A
timestamp 1666464484
transform -1 0 79304 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output166_A
timestamp 1666464484
transform -1 0 107732 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output167_A
timestamp 1666464484
transform -1 0 109756 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output168_A
timestamp 1666464484
transform -1 0 112332 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output169_A
timestamp 1666464484
transform -1 0 113620 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output170_A
timestamp 1666464484
transform 1 0 115276 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output171_A
timestamp 1666464484
transform -1 0 117300 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output172_A
timestamp 1666464484
transform -1 0 119324 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output173_A
timestamp 1666464484
transform -1 0 121716 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output174_A
timestamp 1666464484
transform -1 0 123188 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output175_A
timestamp 1666464484
transform -1 0 125212 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output176_A
timestamp 1666464484
transform -1 0 84272 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output177_A
timestamp 1666464484
transform -1 0 126500 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output178_A
timestamp 1666464484
transform -1 0 128432 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output179_A
timestamp 1666464484
transform -1 0 129720 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output187_A
timestamp 1666464484
transform -1 0 87124 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output190_A
timestamp 1666464484
transform -1 0 89240 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output191_A
timestamp 1666464484
transform -1 0 93012 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output192_A
timestamp 1666464484
transform -1 0 96048 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output193_A
timestamp 1666464484
transform -1 0 98072 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output194_A
timestamp 1666464484
transform -1 0 100832 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output195_A
timestamp 1666464484
transform -1 0 104604 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output196_A
timestamp 1666464484
transform -1 0 106444 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output200_A
timestamp 1666464484
transform 1 0 62928 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output202_A
timestamp 1666464484
transform 1 0 72312 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output205_A
timestamp 1666464484
transform -1 0 86572 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output206_A
timestamp 1666464484
transform 1 0 87584 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output207_A
timestamp 1666464484
transform 1 0 91724 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output208_A
timestamp 1666464484
transform 1 0 96048 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output210_A
timestamp 1666464484
transform 1 0 100004 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output211_A
timestamp 1666464484
transform 1 0 104512 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output212_A
timestamp 1666464484
transform 1 0 108928 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output213_A
timestamp 1666464484
transform 1 0 112424 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output214_A
timestamp 1666464484
transform 1 0 116656 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output215_A
timestamp 1666464484
transform 1 0 120704 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output216_A
timestamp 1666464484
transform 1 0 125212 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output217_A
timestamp 1666464484
transform 1 0 129536 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output218_A
timestamp 1666464484
transform 1 0 133124 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output219_A
timestamp 1666464484
transform 1 0 137264 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output221_A
timestamp 1666464484
transform 1 0 141404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output222_A
timestamp 1666464484
transform 1 0 145912 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output230_A
timestamp 1666464484
transform -1 0 4600 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output236_A
timestamp 1666464484
transform -1 0 80040 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output237_A
timestamp 1666464484
transform -1 0 83996 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output238_A
timestamp 1666464484
transform -1 0 88228 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output239_A
timestamp 1666464484
transform -1 0 91724 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33
timestamp 1666464484
transform 1 0 4140 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1666464484
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1666464484
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94
timestamp 1666464484
transform 1 0 9752 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100
timestamp 1666464484
transform 1 0 10304 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_125
timestamp 1666464484
transform 1 0 12604 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_133 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1666464484
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_149
timestamp 1666464484
transform 1 0 14812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_157
timestamp 1666464484
transform 1 0 15548 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1666464484
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_185
timestamp 1666464484
transform 1 0 18124 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_191
timestamp 1666464484
transform 1 0 18676 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1666464484
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1666464484
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_203
timestamp 1666464484
transform 1 0 19780 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_209
timestamp 1666464484
transform 1 0 20332 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_214
timestamp 1666464484
transform 1 0 20792 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1666464484
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1666464484
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_247
timestamp 1666464484
transform 1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1666464484
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_253
timestamp 1666464484
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_260
timestamp 1666464484
transform 1 0 25024 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_270
timestamp 1666464484
transform 1 0 25944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1666464484
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1666464484
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_303
timestamp 1666464484
transform 1 0 28980 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1666464484
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_309
timestamp 1666464484
transform 1 0 29532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1666464484
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1666464484
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_359
timestamp 1666464484
transform 1 0 34132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1666464484
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1666464484
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_387
timestamp 1666464484
transform 1 0 36708 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1666464484
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1666464484
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_415
timestamp 1666464484
transform 1 0 39284 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1666464484
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1666464484
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_432
timestamp 1666464484
transform 1 0 40848 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_438
timestamp 1666464484
transform 1 0 41400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1666464484
transform 1 0 42136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1666464484
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_471
timestamp 1666464484
transform 1 0 44436 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1666464484
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_477
timestamp 1666464484
transform 1 0 44988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_481
timestamp 1666464484
transform 1 0 45356 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_502
timestamp 1666464484
transform 1 0 47288 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_505
timestamp 1666464484
transform 1 0 47564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_527
timestamp 1666464484
transform 1 0 49588 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_531
timestamp 1666464484
transform 1 0 49956 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_533
timestamp 1666464484
transform 1 0 50140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_537
timestamp 1666464484
transform 1 0 50508 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_558
timestamp 1666464484
transform 1 0 52440 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_561
timestamp 1666464484
transform 1 0 52716 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_567
timestamp 1666464484
transform 1 0 53268 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_572
timestamp 1666464484
transform 1 0 53728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_582
timestamp 1666464484
transform 1 0 54648 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_589
timestamp 1666464484
transform 1 0 55292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_614
timestamp 1666464484
transform 1 0 57592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_617
timestamp 1666464484
transform 1 0 57868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_639
timestamp 1666464484
transform 1 0 59892 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_643
timestamp 1666464484
transform 1 0 60260 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_645
timestamp 1666464484
transform 1 0 60444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_649
timestamp 1666464484
transform 1 0 60812 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_670
timestamp 1666464484
transform 1 0 62744 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_673
timestamp 1666464484
transform 1 0 63020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_695
timestamp 1666464484
transform 1 0 65044 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_699
timestamp 1666464484
transform 1 0 65412 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_701
timestamp 1666464484
transform 1 0 65596 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_724
timestamp 1666464484
transform 1 0 67712 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_729
timestamp 1666464484
transform 1 0 68172 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_735
timestamp 1666464484
transform 1 0 68724 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_740
timestamp 1666464484
transform 1 0 69184 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_747
timestamp 1666464484
transform 1 0 69828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_754
timestamp 1666464484
transform 1 0 70472 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_757
timestamp 1666464484
transform 1 0 70748 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_780
timestamp 1666464484
transform 1 0 72864 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_785
timestamp 1666464484
transform 1 0 73324 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_810
timestamp 1666464484
transform 1 0 75624 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_813
timestamp 1666464484
transform 1 0 75900 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_838
timestamp 1666464484
transform 1 0 78200 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_841
timestamp 1666464484
transform 1 0 78476 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_866
timestamp 1666464484
transform 1 0 80776 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_869
timestamp 1666464484
transform 1 0 81052 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_892
timestamp 1666464484
transform 1 0 83168 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_897
timestamp 1666464484
transform 1 0 83628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_905
timestamp 1666464484
transform 1 0 84364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_912
timestamp 1666464484
transform 1 0 85008 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_920
timestamp 1666464484
transform 1 0 85744 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_925
timestamp 1666464484
transform 1 0 86204 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_929
timestamp 1666464484
transform 1 0 86572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_935
timestamp 1666464484
transform 1 0 87124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_939
timestamp 1666464484
transform 1 0 87492 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_942
timestamp 1666464484
transform 1 0 87768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_950
timestamp 1666464484
transform 1 0 88504 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_953
timestamp 1666464484
transform 1 0 88780 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_957
timestamp 1666464484
transform 1 0 89148 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_965
timestamp 1666464484
transform 1 0 89884 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_977
timestamp 1666464484
transform 1 0 90988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_981
timestamp 1666464484
transform 1 0 91356 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_987
timestamp 1666464484
transform 1 0 91908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_995
timestamp 1666464484
transform 1 0 92644 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1003
timestamp 1666464484
transform 1 0 93380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1006
timestamp 1666464484
transform 1 0 93656 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1009
timestamp 1666464484
transform 1 0 93932 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1015
timestamp 1666464484
transform 1 0 94484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1027
timestamp 1666464484
transform 1 0 95588 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1031
timestamp 1666464484
transform 1 0 95956 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1034
timestamp 1666464484
transform 1 0 96232 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1037
timestamp 1666464484
transform 1 0 96508 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1043
timestamp 1666464484
transform 1 0 97060 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1055
timestamp 1666464484
transform 1 0 98164 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1063
timestamp 1666464484
transform 1 0 98900 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1065
timestamp 1666464484
transform 1 0 99084 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1073
timestamp 1666464484
transform 1 0 99820 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1077
timestamp 1666464484
transform 1 0 100188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1085
timestamp 1666464484
transform 1 0 100924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1091
timestamp 1666464484
transform 1 0 101476 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1093
timestamp 1666464484
transform 1 0 101660 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1100
timestamp 1666464484
transform 1 0 102304 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1112
timestamp 1666464484
transform 1 0 103408 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1121
timestamp 1666464484
transform 1 0 104236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1125
timestamp 1666464484
transform 1 0 104604 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1130
timestamp 1666464484
transform 1 0 105064 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1134
timestamp 1666464484
transform 1 0 105432 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1137
timestamp 1666464484
transform 1 0 105708 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1145
timestamp 1666464484
transform 1 0 106444 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1149
timestamp 1666464484
transform 1 0 106812 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1161
timestamp 1666464484
transform 1 0 107916 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1169
timestamp 1666464484
transform 1 0 108652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1174
timestamp 1666464484
transform 1 0 109112 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1177
timestamp 1666464484
transform 1 0 109388 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1183
timestamp 1666464484
transform 1 0 109940 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1191
timestamp 1666464484
transform 1 0 110676 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1203
timestamp 1666464484
transform 1 0 111780 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1205
timestamp 1666464484
transform 1 0 111964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1209
timestamp 1666464484
transform 1 0 112332 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1212
timestamp 1666464484
transform 1 0 112608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1220
timestamp 1666464484
transform 1 0 113344 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1230
timestamp 1666464484
transform 1 0 114264 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1233
timestamp 1666464484
transform 1 0 114540 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1239
timestamp 1666464484
transform 1 0 115092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1251
timestamp 1666464484
transform 1 0 116196 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1255
timestamp 1666464484
transform 1 0 116564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1258
timestamp 1666464484
transform 1 0 116840 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1261
timestamp 1666464484
transform 1 0 117116 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1267
timestamp 1666464484
transform 1 0 117668 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1275
timestamp 1666464484
transform 1 0 118404 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1280
timestamp 1666464484
transform 1 0 118864 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1289
timestamp 1666464484
transform 1 0 119692 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1297
timestamp 1666464484
transform 1 0 120428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1302
timestamp 1666464484
transform 1 0 120888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1310
timestamp 1666464484
transform 1 0 121624 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1317
timestamp 1666464484
transform 1 0 122268 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1325
timestamp 1666464484
transform 1 0 123004 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1337
timestamp 1666464484
transform 1 0 124108 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1343
timestamp 1666464484
transform 1 0 124660 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1345
timestamp 1666464484
transform 1 0 124844 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1355
timestamp 1666464484
transform 1 0 125764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1359
timestamp 1666464484
transform 1 0 126132 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1362
timestamp 1666464484
transform 1 0 126408 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1370
timestamp 1666464484
transform 1 0 127144 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1373
timestamp 1666464484
transform 1 0 127420 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1385
timestamp 1666464484
transform 1 0 128524 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1393
timestamp 1666464484
transform 1 0 129260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1398
timestamp 1666464484
transform 1 0 129720 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1401
timestamp 1666464484
transform 1 0 129996 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1407
timestamp 1666464484
transform 1 0 130548 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1415
timestamp 1666464484
transform 1 0 131284 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1427
timestamp 1666464484
transform 1 0 132388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1429
timestamp 1666464484
transform 1 0 132572 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1437
timestamp 1666464484
transform 1 0 133308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1445
timestamp 1666464484
transform 1 0 134044 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1451
timestamp 1666464484
transform 1 0 134596 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1454
timestamp 1666464484
transform 1 0 134872 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1457
timestamp 1666464484
transform 1 0 135148 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1463
timestamp 1666464484
transform 1 0 135700 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1475
timestamp 1666464484
transform 1 0 136804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1479
timestamp 1666464484
transform 1 0 137172 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1482
timestamp 1666464484
transform 1 0 137448 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1485
timestamp 1666464484
transform 1 0 137724 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1491
timestamp 1666464484
transform 1 0 138276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1497
timestamp 1666464484
transform 1 0 138828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1505
timestamp 1666464484
transform 1 0 139564 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1511
timestamp 1666464484
transform 1 0 140116 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1513
timestamp 1666464484
transform 1 0 140300 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1527
timestamp 1666464484
transform 1 0 141588 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1535
timestamp 1666464484
transform 1 0 142324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1539
timestamp 1666464484
transform 1 0 142692 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1541
timestamp 1666464484
transform 1 0 142876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1545
timestamp 1666464484
transform 1 0 143244 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1552
timestamp 1666464484
transform 1 0 143888 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1564
timestamp 1666464484
transform 1 0 144992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1569
timestamp 1666464484
transform 1 0 145452 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1575
timestamp 1666464484
transform 1 0 146004 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1580
timestamp 1666464484
transform 1 0 146464 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1594
timestamp 1666464484
transform 1 0 147752 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1597
timestamp 1666464484
transform 1 0 148028 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1601
timestamp 1666464484
transform 1 0 148396 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1666464484
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_27
timestamp 1666464484
transform 1 0 3588 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_35
timestamp 1666464484
transform 1 0 4324 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_40
timestamp 1666464484
transform 1 0 4784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1666464484
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_67
timestamp 1666464484
transform 1 0 7268 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_75
timestamp 1666464484
transform 1 0 8004 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_79
timestamp 1666464484
transform 1 0 8372 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_87
timestamp 1666464484
transform 1 0 9108 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_91
timestamp 1666464484
transform 1 0 9476 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_103
timestamp 1666464484
transform 1 0 10580 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1666464484
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1666464484
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1666464484
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_149
timestamp 1666464484
transform 1 0 14812 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_153
timestamp 1666464484
transform 1 0 15180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 1666464484
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1666464484
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1666464484
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_205
timestamp 1666464484
transform 1 0 19964 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_209
timestamp 1666464484
transform 1 0 20332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1666464484
transform 1 0 20884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1666464484
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1666464484
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_247
timestamp 1666464484
transform 1 0 23828 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_260
timestamp 1666464484
transform 1 0 25024 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_271
timestamp 1666464484
transform 1 0 26036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1666464484
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1666464484
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_294
timestamp 1666464484
transform 1 0 28152 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_307
timestamp 1666464484
transform 1 0 29348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_317
timestamp 1666464484
transform 1 0 30268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_325
timestamp 1666464484
transform 1 0 31004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_329
timestamp 1666464484
transform 1 0 31372 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_334
timestamp 1666464484
transform 1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1666464484
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_341
timestamp 1666464484
transform 1 0 32476 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_351
timestamp 1666464484
transform 1 0 33396 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_364
timestamp 1666464484
transform 1 0 34592 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1666464484
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1666464484
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_404
timestamp 1666464484
transform 1 0 38272 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_410
timestamp 1666464484
transform 1 0 38824 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_431
timestamp 1666464484
transform 1 0 40756 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_446
timestamp 1666464484
transform 1 0 42136 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_449
timestamp 1666464484
transform 1 0 42412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_453
timestamp 1666464484
transform 1 0 42780 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_459
timestamp 1666464484
transform 1 0 43332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_483
timestamp 1666464484
transform 1 0 45540 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_491
timestamp 1666464484
transform 1 0 46276 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_495
timestamp 1666464484
transform 1 0 46644 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_500
timestamp 1666464484
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_505
timestamp 1666464484
transform 1 0 47564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_527
timestamp 1666464484
transform 1 0 49588 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_534
timestamp 1666464484
transform 1 0 50232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_558
timestamp 1666464484
transform 1 0 52440 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_561
timestamp 1666464484
transform 1 0 52716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_572
timestamp 1666464484
transform 1 0 53728 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_599
timestamp 1666464484
transform 1 0 56212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_606
timestamp 1666464484
transform 1 0 56856 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_614
timestamp 1666464484
transform 1 0 57592 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_617
timestamp 1666464484
transform 1 0 57868 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_628
timestamp 1666464484
transform 1 0 58880 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_636
timestamp 1666464484
transform 1 0 59616 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_657
timestamp 1666464484
transform 1 0 61548 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_667
timestamp 1666464484
transform 1 0 62468 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1666464484
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_673
timestamp 1666464484
transform 1 0 63020 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_684
timestamp 1666464484
transform 1 0 64032 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_688
timestamp 1666464484
transform 1 0 64400 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_693
timestamp 1666464484
transform 1 0 64860 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_718
timestamp 1666464484
transform 1 0 67160 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_726
timestamp 1666464484
transform 1 0 67896 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_729
timestamp 1666464484
transform 1 0 68172 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_735
timestamp 1666464484
transform 1 0 68724 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_739
timestamp 1666464484
transform 1 0 69092 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_746
timestamp 1666464484
transform 1 0 69736 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_771
timestamp 1666464484
transform 1 0 72036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_779
timestamp 1666464484
transform 1 0 72772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_783
timestamp 1666464484
transform 1 0 73140 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_785
timestamp 1666464484
transform 1 0 73324 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_791
timestamp 1666464484
transform 1 0 73876 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_798
timestamp 1666464484
transform 1 0 74520 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_807
timestamp 1666464484
transform 1 0 75348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_815
timestamp 1666464484
transform 1 0 76084 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_821
timestamp 1666464484
transform 1 0 76636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_825
timestamp 1666464484
transform 1 0 77004 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_830
timestamp 1666464484
transform 1 0 77464 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_838
timestamp 1666464484
transform 1 0 78200 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_841
timestamp 1666464484
transform 1 0 78476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_845
timestamp 1666464484
transform 1 0 78844 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_872
timestamp 1666464484
transform 1 0 81328 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_885
timestamp 1666464484
transform 1 0 82524 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_893
timestamp 1666464484
transform 1 0 83260 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_897
timestamp 1666464484
transform 1 0 83628 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_902
timestamp 1666464484
transform 1 0 84088 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_908
timestamp 1666464484
transform 1 0 84640 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_914
timestamp 1666464484
transform 1 0 85192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_920
timestamp 1666464484
transform 1 0 85744 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_926
timestamp 1666464484
transform 1 0 86296 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_938
timestamp 1666464484
transform 1 0 87400 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_950
timestamp 1666464484
transform 1 0 88504 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_953
timestamp 1666464484
transform 1 0 88780 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_965
timestamp 1666464484
transform 1 0 89884 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_977
timestamp 1666464484
transform 1 0 90988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_989
timestamp 1666464484
transform 1 0 92092 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1001
timestamp 1666464484
transform 1 0 93196 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1007
timestamp 1666464484
transform 1 0 93748 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1009
timestamp 1666464484
transform 1 0 93932 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1021
timestamp 1666464484
transform 1 0 95036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1033
timestamp 1666464484
transform 1 0 96140 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1045
timestamp 1666464484
transform 1 0 97244 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1051
timestamp 1666464484
transform 1 0 97796 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1063
timestamp 1666464484
transform 1 0 98900 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1065
timestamp 1666464484
transform 1 0 99084 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1077
timestamp 1666464484
transform 1 0 100188 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1089
timestamp 1666464484
transform 1 0 101292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1093
timestamp 1666464484
transform 1 0 101660 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1096
timestamp 1666464484
transform 1 0 101936 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1108
timestamp 1666464484
transform 1 0 103040 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1121
timestamp 1666464484
transform 1 0 104236 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1126
timestamp 1666464484
transform 1 0 104696 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1138
timestamp 1666464484
transform 1 0 105800 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1150
timestamp 1666464484
transform 1 0 106904 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1162
timestamp 1666464484
transform 1 0 108008 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1174
timestamp 1666464484
transform 1 0 109112 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1177
timestamp 1666464484
transform 1 0 109388 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1187
timestamp 1666464484
transform 1 0 110308 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1199
timestamp 1666464484
transform 1 0 111412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1211
timestamp 1666464484
transform 1 0 112516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1223
timestamp 1666464484
transform 1 0 113620 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1231
timestamp 1666464484
transform 1 0 114356 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1233
timestamp 1666464484
transform 1 0 114540 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1245
timestamp 1666464484
transform 1 0 115644 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1257
timestamp 1666464484
transform 1 0 116748 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1269
timestamp 1666464484
transform 1 0 117852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1273
timestamp 1666464484
transform 1 0 118220 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1276
timestamp 1666464484
transform 1 0 118496 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1289
timestamp 1666464484
transform 1 0 119692 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1301
timestamp 1666464484
transform 1 0 120796 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1313
timestamp 1666464484
transform 1 0 121900 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1321
timestamp 1666464484
transform 1 0 122636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1333
timestamp 1666464484
transform 1 0 123740 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1341
timestamp 1666464484
transform 1 0 124476 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1345
timestamp 1666464484
transform 1 0 124844 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1351
timestamp 1666464484
transform 1 0 125396 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1363
timestamp 1666464484
transform 1 0 126500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1375
timestamp 1666464484
transform 1 0 127604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1387
timestamp 1666464484
transform 1 0 128708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1399
timestamp 1666464484
transform 1 0 129812 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1401
timestamp 1666464484
transform 1 0 129996 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1411
timestamp 1666464484
transform 1 0 130916 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1423
timestamp 1666464484
transform 1 0 132020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1435
timestamp 1666464484
transform 1 0 133124 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1447
timestamp 1666464484
transform 1 0 134228 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1455
timestamp 1666464484
transform 1 0 134964 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1457
timestamp 1666464484
transform 1 0 135148 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1469
timestamp 1666464484
transform 1 0 136252 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1481
timestamp 1666464484
transform 1 0 137356 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1493
timestamp 1666464484
transform 1 0 138460 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1505
timestamp 1666464484
transform 1 0 139564 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1511
timestamp 1666464484
transform 1 0 140116 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1513
timestamp 1666464484
transform 1 0 140300 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1525
timestamp 1666464484
transform 1 0 141404 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1537
timestamp 1666464484
transform 1 0 142508 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1543
timestamp 1666464484
transform 1 0 143060 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1546
timestamp 1666464484
transform 1 0 143336 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1558
timestamp 1666464484
transform 1 0 144440 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1566
timestamp 1666464484
transform 1 0 145176 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1569
timestamp 1666464484
transform 1 0 145452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1573
timestamp 1666464484
transform 1 0 145820 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1576
timestamp 1666464484
transform 1 0 146096 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1588
timestamp 1666464484
transform 1 0 147200 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1600
timestamp 1666464484
transform 1 0 148304 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1666464484
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1666464484
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_37
timestamp 1666464484
transform 1 0 4508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_42
timestamp 1666464484
transform 1 0 4968 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_49
timestamp 1666464484
transform 1 0 5612 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_53
timestamp 1666464484
transform 1 0 5980 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_57
timestamp 1666464484
transform 1 0 6348 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_64
timestamp 1666464484
transform 1 0 6992 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_72
timestamp 1666464484
transform 1 0 7728 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_76
timestamp 1666464484
transform 1 0 8096 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1666464484
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_89
timestamp 1666464484
transform 1 0 9292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_101
timestamp 1666464484
transform 1 0 10396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_113
timestamp 1666464484
transform 1 0 11500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_125
timestamp 1666464484
transform 1 0 12604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_137
timestamp 1666464484
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1666464484
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1666464484
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1666464484
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1666464484
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1666464484
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1666464484
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_211
timestamp 1666464484
transform 1 0 20516 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_217
timestamp 1666464484
transform 1 0 21068 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_224
timestamp 1666464484
transform 1 0 21712 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_231
timestamp 1666464484
transform 1 0 22356 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_244
timestamp 1666464484
transform 1 0 23552 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1666464484
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1666464484
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_257
timestamp 1666464484
transform 1 0 24748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_263
timestamp 1666464484
transform 1 0 25300 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_269
timestamp 1666464484
transform 1 0 25852 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_293
timestamp 1666464484
transform 1 0 28060 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_305
timestamp 1666464484
transform 1 0 29164 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_309
timestamp 1666464484
transform 1 0 29532 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_315
timestamp 1666464484
transform 1 0 30084 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_318
timestamp 1666464484
transform 1 0 30360 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_325
timestamp 1666464484
transform 1 0 31004 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_333
timestamp 1666464484
transform 1 0 31740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_336
timestamp 1666464484
transform 1 0 32016 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_342
timestamp 1666464484
transform 1 0 32568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_350
timestamp 1666464484
transform 1 0 33304 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_358
timestamp 1666464484
transform 1 0 34040 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_362
timestamp 1666464484
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_365
timestamp 1666464484
transform 1 0 34684 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_380
timestamp 1666464484
transform 1 0 36064 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_404
timestamp 1666464484
transform 1 0 38272 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_412
timestamp 1666464484
transform 1 0 39008 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_418
timestamp 1666464484
transform 1 0 39560 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1666464484
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_427
timestamp 1666464484
transform 1 0 40388 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_431
timestamp 1666464484
transform 1 0 40756 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_436
timestamp 1666464484
transform 1 0 41216 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_460
timestamp 1666464484
transform 1 0 43424 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_473
timestamp 1666464484
transform 1 0 44620 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_477
timestamp 1666464484
transform 1 0 44988 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_482
timestamp 1666464484
transform 1 0 45448 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_493
timestamp 1666464484
transform 1 0 46460 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_517
timestamp 1666464484
transform 1 0 48668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_527
timestamp 1666464484
transform 1 0 49588 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1666464484
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_533
timestamp 1666464484
transform 1 0 50140 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_537
timestamp 1666464484
transform 1 0 50508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_545
timestamp 1666464484
transform 1 0 51244 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_551
timestamp 1666464484
transform 1 0 51796 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_561
timestamp 1666464484
transform 1 0 52716 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_567
timestamp 1666464484
transform 1 0 53268 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_575
timestamp 1666464484
transform 1 0 54004 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_586
timestamp 1666464484
transform 1 0 55016 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_589
timestamp 1666464484
transform 1 0 55292 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_595
timestamp 1666464484
transform 1 0 55844 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_605
timestamp 1666464484
transform 1 0 56764 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_611
timestamp 1666464484
transform 1 0 57316 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_621
timestamp 1666464484
transform 1 0 58236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_627
timestamp 1666464484
transform 1 0 58788 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_635
timestamp 1666464484
transform 1 0 59524 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_642
timestamp 1666464484
transform 1 0 60168 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_645
timestamp 1666464484
transform 1 0 60444 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_656
timestamp 1666464484
transform 1 0 61456 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_663
timestamp 1666464484
transform 1 0 62100 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_670
timestamp 1666464484
transform 1 0 62744 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_685
timestamp 1666464484
transform 1 0 64124 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_698
timestamp 1666464484
transform 1 0 65320 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_701
timestamp 1666464484
transform 1 0 65596 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_707
timestamp 1666464484
transform 1 0 66148 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_714
timestamp 1666464484
transform 1 0 66792 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_721
timestamp 1666464484
transform 1 0 67436 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_727
timestamp 1666464484
transform 1 0 67988 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_737
timestamp 1666464484
transform 1 0 68908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_750
timestamp 1666464484
transform 1 0 70104 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_757
timestamp 1666464484
transform 1 0 70748 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_768
timestamp 1666464484
transform 1 0 71760 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_774
timestamp 1666464484
transform 1 0 72312 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_780
timestamp 1666464484
transform 1 0 72864 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_783
timestamp 1666464484
transform 1 0 73140 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_789
timestamp 1666464484
transform 1 0 73692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_796
timestamp 1666464484
transform 1 0 74336 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_800
timestamp 1666464484
transform 1 0 74704 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_810
timestamp 1666464484
transform 1 0 75624 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_813
timestamp 1666464484
transform 1 0 75900 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_817
timestamp 1666464484
transform 1 0 76268 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_824
timestamp 1666464484
transform 1 0 76912 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_837
timestamp 1666464484
transform 1 0 78108 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_862
timestamp 1666464484
transform 1 0 80408 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_869
timestamp 1666464484
transform 1 0 81052 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_880
timestamp 1666464484
transform 1 0 82064 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_893
timestamp 1666464484
transform 1 0 83260 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_899
timestamp 1666464484
transform 1 0 83812 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_905
timestamp 1666464484
transform 1 0 84364 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_911
timestamp 1666464484
transform 1 0 84916 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_917
timestamp 1666464484
transform 1 0 85468 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_923
timestamp 1666464484
transform 1 0 86020 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_925
timestamp 1666464484
transform 1 0 86204 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_937
timestamp 1666464484
transform 1 0 87308 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_949
timestamp 1666464484
transform 1 0 88412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_961
timestamp 1666464484
transform 1 0 89516 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_973
timestamp 1666464484
transform 1 0 90620 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_979
timestamp 1666464484
transform 1 0 91172 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_981
timestamp 1666464484
transform 1 0 91356 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_993
timestamp 1666464484
transform 1 0 92460 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1005
timestamp 1666464484
transform 1 0 93564 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1017
timestamp 1666464484
transform 1 0 94668 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1029
timestamp 1666464484
transform 1 0 95772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1035
timestamp 1666464484
transform 1 0 96324 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1037
timestamp 1666464484
transform 1 0 96508 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1049
timestamp 1666464484
transform 1 0 97612 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1061
timestamp 1666464484
transform 1 0 98716 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1073
timestamp 1666464484
transform 1 0 99820 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1085
timestamp 1666464484
transform 1 0 100924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1091
timestamp 1666464484
transform 1 0 101476 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1093
timestamp 1666464484
transform 1 0 101660 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1105
timestamp 1666464484
transform 1 0 102764 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1117
timestamp 1666464484
transform 1 0 103868 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1129
timestamp 1666464484
transform 1 0 104972 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1141
timestamp 1666464484
transform 1 0 106076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1147
timestamp 1666464484
transform 1 0 106628 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1149
timestamp 1666464484
transform 1 0 106812 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1161
timestamp 1666464484
transform 1 0 107916 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1173
timestamp 1666464484
transform 1 0 109020 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1185
timestamp 1666464484
transform 1 0 110124 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1197
timestamp 1666464484
transform 1 0 111228 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1203
timestamp 1666464484
transform 1 0 111780 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1205
timestamp 1666464484
transform 1 0 111964 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1217
timestamp 1666464484
transform 1 0 113068 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1229
timestamp 1666464484
transform 1 0 114172 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1241
timestamp 1666464484
transform 1 0 115276 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1253
timestamp 1666464484
transform 1 0 116380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1259
timestamp 1666464484
transform 1 0 116932 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1261
timestamp 1666464484
transform 1 0 117116 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1273
timestamp 1666464484
transform 1 0 118220 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1285
timestamp 1666464484
transform 1 0 119324 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1297
timestamp 1666464484
transform 1 0 120428 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1309
timestamp 1666464484
transform 1 0 121532 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1315
timestamp 1666464484
transform 1 0 122084 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1317
timestamp 1666464484
transform 1 0 122268 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1329
timestamp 1666464484
transform 1 0 123372 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1341
timestamp 1666464484
transform 1 0 124476 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1353
timestamp 1666464484
transform 1 0 125580 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1365
timestamp 1666464484
transform 1 0 126684 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1371
timestamp 1666464484
transform 1 0 127236 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1373
timestamp 1666464484
transform 1 0 127420 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1385
timestamp 1666464484
transform 1 0 128524 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1397
timestamp 1666464484
transform 1 0 129628 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1409
timestamp 1666464484
transform 1 0 130732 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1421
timestamp 1666464484
transform 1 0 131836 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1427
timestamp 1666464484
transform 1 0 132388 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1429
timestamp 1666464484
transform 1 0 132572 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1441
timestamp 1666464484
transform 1 0 133676 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1453
timestamp 1666464484
transform 1 0 134780 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1465
timestamp 1666464484
transform 1 0 135884 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1477
timestamp 1666464484
transform 1 0 136988 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1483
timestamp 1666464484
transform 1 0 137540 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1485
timestamp 1666464484
transform 1 0 137724 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1497
timestamp 1666464484
transform 1 0 138828 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1509
timestamp 1666464484
transform 1 0 139932 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1521
timestamp 1666464484
transform 1 0 141036 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1533
timestamp 1666464484
transform 1 0 142140 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1539
timestamp 1666464484
transform 1 0 142692 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1541
timestamp 1666464484
transform 1 0 142876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1553
timestamp 1666464484
transform 1 0 143980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1565
timestamp 1666464484
transform 1 0 145084 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1577
timestamp 1666464484
transform 1 0 146188 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1589
timestamp 1666464484
transform 1 0 147292 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1595
timestamp 1666464484
transform 1 0 147844 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1597
timestamp 1666464484
transform 1 0 148028 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1666464484
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1666464484
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1666464484
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_51
timestamp 1666464484
transform 1 0 5796 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1666464484
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_62
timestamp 1666464484
transform 1 0 6808 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_68
timestamp 1666464484
transform 1 0 7360 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_76
timestamp 1666464484
transform 1 0 8096 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_88
timestamp 1666464484
transform 1 0 9200 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_100
timestamp 1666464484
transform 1 0 10304 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1666464484
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1666464484
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1666464484
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1666464484
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1666464484
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1666464484
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1666464484
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1666464484
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1666464484
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1666464484
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_225
timestamp 1666464484
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_229
timestamp 1666464484
transform 1 0 22172 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_233
timestamp 1666464484
transform 1 0 22540 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_245
timestamp 1666464484
transform 1 0 23644 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_251
timestamp 1666464484
transform 1 0 24196 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_257
timestamp 1666464484
transform 1 0 24748 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_269
timestamp 1666464484
transform 1 0 25852 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_272
timestamp 1666464484
transform 1 0 26128 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1666464484
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1666464484
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_286
timestamp 1666464484
transform 1 0 27416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_293
timestamp 1666464484
transform 1 0 28060 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_299
timestamp 1666464484
transform 1 0 28612 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_305
timestamp 1666464484
transform 1 0 29164 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_311
timestamp 1666464484
transform 1 0 29716 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_321
timestamp 1666464484
transform 1 0 30636 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_329
timestamp 1666464484
transform 1 0 31372 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp 1666464484
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_337
timestamp 1666464484
transform 1 0 32108 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_345
timestamp 1666464484
transform 1 0 32844 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_352
timestamp 1666464484
transform 1 0 33488 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_359
timestamp 1666464484
transform 1 0 34132 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_367
timestamp 1666464484
transform 1 0 34868 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_372
timestamp 1666464484
transform 1 0 35328 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_380
timestamp 1666464484
transform 1 0 36064 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_387
timestamp 1666464484
transform 1 0 36708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1666464484
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_393
timestamp 1666464484
transform 1 0 37260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_399
timestamp 1666464484
transform 1 0 37812 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_406
timestamp 1666464484
transform 1 0 38456 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_417
timestamp 1666464484
transform 1 0 39468 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_424
timestamp 1666464484
transform 1 0 40112 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_430
timestamp 1666464484
transform 1 0 40664 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_433
timestamp 1666464484
transform 1 0 40940 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_439
timestamp 1666464484
transform 1 0 41492 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_446
timestamp 1666464484
transform 1 0 42136 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_449
timestamp 1666464484
transform 1 0 42412 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_456
timestamp 1666464484
transform 1 0 43056 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_464
timestamp 1666464484
transform 1 0 43792 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_472
timestamp 1666464484
transform 1 0 44528 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_476
timestamp 1666464484
transform 1 0 44896 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_479
timestamp 1666464484
transform 1 0 45172 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_485
timestamp 1666464484
transform 1 0 45724 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_492
timestamp 1666464484
transform 1 0 46368 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_496
timestamp 1666464484
transform 1 0 46736 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_500
timestamp 1666464484
transform 1 0 47104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_505
timestamp 1666464484
transform 1 0 47564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_516
timestamp 1666464484
transform 1 0 48576 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_522
timestamp 1666464484
transform 1 0 49128 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_530
timestamp 1666464484
transform 1 0 49864 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_534
timestamp 1666464484
transform 1 0 50232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_537
timestamp 1666464484
transform 1 0 50508 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_544
timestamp 1666464484
transform 1 0 51152 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_551
timestamp 1666464484
transform 1 0 51796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_558
timestamp 1666464484
transform 1 0 52440 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_561
timestamp 1666464484
transform 1 0 52716 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_567
timestamp 1666464484
transform 1 0 53268 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_577
timestamp 1666464484
transform 1 0 54188 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_583
timestamp 1666464484
transform 1 0 54740 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_590
timestamp 1666464484
transform 1 0 55384 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_594
timestamp 1666464484
transform 1 0 55752 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_597
timestamp 1666464484
transform 1 0 56028 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_605
timestamp 1666464484
transform 1 0 56764 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_612
timestamp 1666464484
transform 1 0 57408 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_617
timestamp 1666464484
transform 1 0 57868 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_622
timestamp 1666464484
transform 1 0 58328 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_632
timestamp 1666464484
transform 1 0 59248 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_642
timestamp 1666464484
transform 1 0 60168 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_650
timestamp 1666464484
transform 1 0 60904 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_657
timestamp 1666464484
transform 1 0 61548 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_668
timestamp 1666464484
transform 1 0 62560 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_673
timestamp 1666464484
transform 1 0 63020 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_680
timestamp 1666464484
transform 1 0 63664 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_686
timestamp 1666464484
transform 1 0 64216 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_696
timestamp 1666464484
transform 1 0 65136 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_703
timestamp 1666464484
transform 1 0 65780 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_712
timestamp 1666464484
transform 1 0 66608 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_720
timestamp 1666464484
transform 1 0 67344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_726
timestamp 1666464484
transform 1 0 67896 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_729
timestamp 1666464484
transform 1 0 68172 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_738
timestamp 1666464484
transform 1 0 69000 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_763
timestamp 1666464484
transform 1 0 71300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_767
timestamp 1666464484
transform 1 0 71668 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_770
timestamp 1666464484
transform 1 0 71944 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_776
timestamp 1666464484
transform 1 0 72496 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_785
timestamp 1666464484
transform 1 0 73324 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_789
timestamp 1666464484
transform 1 0 73692 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_797
timestamp 1666464484
transform 1 0 74428 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_801
timestamp 1666464484
transform 1 0 74796 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_809
timestamp 1666464484
transform 1 0 75532 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_812
timestamp 1666464484
transform 1 0 75808 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_822
timestamp 1666464484
transform 1 0 76728 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_828
timestamp 1666464484
transform 1 0 77280 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_834
timestamp 1666464484
transform 1 0 77832 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_838
timestamp 1666464484
transform 1 0 78200 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_841
timestamp 1666464484
transform 1 0 78476 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_847
timestamp 1666464484
transform 1 0 79028 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_869
timestamp 1666464484
transform 1 0 81052 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_882
timestamp 1666464484
transform 1 0 82248 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_888
timestamp 1666464484
transform 1 0 82800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_894
timestamp 1666464484
transform 1 0 83352 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_897
timestamp 1666464484
transform 1 0 83628 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_901
timestamp 1666464484
transform 1 0 83996 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_907
timestamp 1666464484
transform 1 0 84548 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_919
timestamp 1666464484
transform 1 0 85652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_931
timestamp 1666464484
transform 1 0 86756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_943
timestamp 1666464484
transform 1 0 87860 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_951
timestamp 1666464484
transform 1 0 88596 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_953
timestamp 1666464484
transform 1 0 88780 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_965
timestamp 1666464484
transform 1 0 89884 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_977
timestamp 1666464484
transform 1 0 90988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_989
timestamp 1666464484
transform 1 0 92092 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1001
timestamp 1666464484
transform 1 0 93196 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1007
timestamp 1666464484
transform 1 0 93748 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1009
timestamp 1666464484
transform 1 0 93932 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1021
timestamp 1666464484
transform 1 0 95036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1033
timestamp 1666464484
transform 1 0 96140 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1045
timestamp 1666464484
transform 1 0 97244 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1057
timestamp 1666464484
transform 1 0 98348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1063
timestamp 1666464484
transform 1 0 98900 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1065
timestamp 1666464484
transform 1 0 99084 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1077
timestamp 1666464484
transform 1 0 100188 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1089
timestamp 1666464484
transform 1 0 101292 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1101
timestamp 1666464484
transform 1 0 102396 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1113
timestamp 1666464484
transform 1 0 103500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1119
timestamp 1666464484
transform 1 0 104052 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1121
timestamp 1666464484
transform 1 0 104236 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1133
timestamp 1666464484
transform 1 0 105340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1145
timestamp 1666464484
transform 1 0 106444 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1157
timestamp 1666464484
transform 1 0 107548 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1169
timestamp 1666464484
transform 1 0 108652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1175
timestamp 1666464484
transform 1 0 109204 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1177
timestamp 1666464484
transform 1 0 109388 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1189
timestamp 1666464484
transform 1 0 110492 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1201
timestamp 1666464484
transform 1 0 111596 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1213
timestamp 1666464484
transform 1 0 112700 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1225
timestamp 1666464484
transform 1 0 113804 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1231
timestamp 1666464484
transform 1 0 114356 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1233
timestamp 1666464484
transform 1 0 114540 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1245
timestamp 1666464484
transform 1 0 115644 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1257
timestamp 1666464484
transform 1 0 116748 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1269
timestamp 1666464484
transform 1 0 117852 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1281
timestamp 1666464484
transform 1 0 118956 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1287
timestamp 1666464484
transform 1 0 119508 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1289
timestamp 1666464484
transform 1 0 119692 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1301
timestamp 1666464484
transform 1 0 120796 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1313
timestamp 1666464484
transform 1 0 121900 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1325
timestamp 1666464484
transform 1 0 123004 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1337
timestamp 1666464484
transform 1 0 124108 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1343
timestamp 1666464484
transform 1 0 124660 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1345
timestamp 1666464484
transform 1 0 124844 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1357
timestamp 1666464484
transform 1 0 125948 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1369
timestamp 1666464484
transform 1 0 127052 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1381
timestamp 1666464484
transform 1 0 128156 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1393
timestamp 1666464484
transform 1 0 129260 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1399
timestamp 1666464484
transform 1 0 129812 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1401
timestamp 1666464484
transform 1 0 129996 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1413
timestamp 1666464484
transform 1 0 131100 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1425
timestamp 1666464484
transform 1 0 132204 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1437
timestamp 1666464484
transform 1 0 133308 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1449
timestamp 1666464484
transform 1 0 134412 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1455
timestamp 1666464484
transform 1 0 134964 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1457
timestamp 1666464484
transform 1 0 135148 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1469
timestamp 1666464484
transform 1 0 136252 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1481
timestamp 1666464484
transform 1 0 137356 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1493
timestamp 1666464484
transform 1 0 138460 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1505
timestamp 1666464484
transform 1 0 139564 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1511
timestamp 1666464484
transform 1 0 140116 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1513
timestamp 1666464484
transform 1 0 140300 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1525
timestamp 1666464484
transform 1 0 141404 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1537
timestamp 1666464484
transform 1 0 142508 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1549
timestamp 1666464484
transform 1 0 143612 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1561
timestamp 1666464484
transform 1 0 144716 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1567
timestamp 1666464484
transform 1 0 145268 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1569
timestamp 1666464484
transform 1 0 145452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1581
timestamp 1666464484
transform 1 0 146556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1593
timestamp 1666464484
transform 1 0 147660 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1601
timestamp 1666464484
transform 1 0 148396 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1666464484
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1666464484
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1666464484
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_53
timestamp 1666464484
transform 1 0 5980 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_58
timestamp 1666464484
transform 1 0 6440 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_70
timestamp 1666464484
transform 1 0 7544 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1666464484
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1666464484
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1666464484
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1666464484
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1666464484
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1666464484
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1666464484
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1666464484
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1666464484
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1666464484
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1666464484
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1666464484
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1666464484
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1666464484
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_235
timestamp 1666464484
transform 1 0 22724 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 1666464484
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1666464484
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1666464484
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_277
timestamp 1666464484
transform 1 0 26588 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_285
timestamp 1666464484
transform 1 0 27324 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_289
timestamp 1666464484
transform 1 0 27692 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_295
timestamp 1666464484
transform 1 0 28244 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_305
timestamp 1666464484
transform 1 0 29164 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_309
timestamp 1666464484
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_313
timestamp 1666464484
transform 1 0 29900 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_319
timestamp 1666464484
transform 1 0 30452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_331
timestamp 1666464484
transform 1 0 31556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_336
timestamp 1666464484
transform 1 0 32016 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_342
timestamp 1666464484
transform 1 0 32568 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_345
timestamp 1666464484
transform 1 0 32844 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_355
timestamp 1666464484
transform 1 0 33764 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_359
timestamp 1666464484
transform 1 0 34132 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_362
timestamp 1666464484
transform 1 0 34408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_365
timestamp 1666464484
transform 1 0 34684 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_373
timestamp 1666464484
transform 1 0 35420 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_380
timestamp 1666464484
transform 1 0 36064 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_386
timestamp 1666464484
transform 1 0 36616 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_389
timestamp 1666464484
transform 1 0 36892 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_395
timestamp 1666464484
transform 1 0 37444 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_403
timestamp 1666464484
transform 1 0 38180 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_411
timestamp 1666464484
transform 1 0 38916 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_415
timestamp 1666464484
transform 1 0 39284 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_418
timestamp 1666464484
transform 1 0 39560 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_421
timestamp 1666464484
transform 1 0 39836 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_425
timestamp 1666464484
transform 1 0 40204 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_431
timestamp 1666464484
transform 1 0 40756 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_437
timestamp 1666464484
transform 1 0 41308 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_445
timestamp 1666464484
transform 1 0 42044 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_452
timestamp 1666464484
transform 1 0 42688 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_462
timestamp 1666464484
transform 1 0 43608 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_474
timestamp 1666464484
transform 1 0 44712 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_477
timestamp 1666464484
transform 1 0 44988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_482
timestamp 1666464484
transform 1 0 45448 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_490
timestamp 1666464484
transform 1 0 46184 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_495
timestamp 1666464484
transform 1 0 46644 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_508
timestamp 1666464484
transform 1 0 47840 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_516
timestamp 1666464484
transform 1 0 48576 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_522
timestamp 1666464484
transform 1 0 49128 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_528
timestamp 1666464484
transform 1 0 49680 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_533
timestamp 1666464484
transform 1 0 50140 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_537
timestamp 1666464484
transform 1 0 50508 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_552
timestamp 1666464484
transform 1 0 51888 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_560
timestamp 1666464484
transform 1 0 52624 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_563
timestamp 1666464484
transform 1 0 52900 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_571
timestamp 1666464484
transform 1 0 53636 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_574
timestamp 1666464484
transform 1 0 53912 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_580
timestamp 1666464484
transform 1 0 54464 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_589
timestamp 1666464484
transform 1 0 55292 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_595
timestamp 1666464484
transform 1 0 55844 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_598
timestamp 1666464484
transform 1 0 56120 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_604
timestamp 1666464484
transform 1 0 56672 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_611
timestamp 1666464484
transform 1 0 57316 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_619
timestamp 1666464484
transform 1 0 58052 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_625
timestamp 1666464484
transform 1 0 58604 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_631
timestamp 1666464484
transform 1 0 59156 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1666464484
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_645
timestamp 1666464484
transform 1 0 60444 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_651
timestamp 1666464484
transform 1 0 60996 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_654
timestamp 1666464484
transform 1 0 61272 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_660
timestamp 1666464484
transform 1 0 61824 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_667
timestamp 1666464484
transform 1 0 62468 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_671
timestamp 1666464484
transform 1 0 62836 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_674
timestamp 1666464484
transform 1 0 63112 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_680
timestamp 1666464484
transform 1 0 63664 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_690
timestamp 1666464484
transform 1 0 64584 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_694
timestamp 1666464484
transform 1 0 64952 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_698
timestamp 1666464484
transform 1 0 65320 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_701
timestamp 1666464484
transform 1 0 65596 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_705
timestamp 1666464484
transform 1 0 65964 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_708
timestamp 1666464484
transform 1 0 66240 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_714
timestamp 1666464484
transform 1 0 66792 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_724
timestamp 1666464484
transform 1 0 67712 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_730
timestamp 1666464484
transform 1 0 68264 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_736
timestamp 1666464484
transform 1 0 68816 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_742
timestamp 1666464484
transform 1 0 69368 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_746
timestamp 1666464484
transform 1 0 69736 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_750
timestamp 1666464484
transform 1 0 70104 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_757
timestamp 1666464484
transform 1 0 70748 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_761
timestamp 1666464484
transform 1 0 71116 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_767
timestamp 1666464484
transform 1 0 71668 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_779
timestamp 1666464484
transform 1 0 72772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_791
timestamp 1666464484
transform 1 0 73876 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_799
timestamp 1666464484
transform 1 0 74612 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_804
timestamp 1666464484
transform 1 0 75072 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_813
timestamp 1666464484
transform 1 0 75900 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_825
timestamp 1666464484
transform 1 0 77004 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_833
timestamp 1666464484
transform 1 0 77740 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_839
timestamp 1666464484
transform 1 0 78292 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_845
timestamp 1666464484
transform 1 0 78844 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_858
timestamp 1666464484
transform 1 0 80040 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_865
timestamp 1666464484
transform 1 0 80684 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_869
timestamp 1666464484
transform 1 0 81052 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_874
timestamp 1666464484
transform 1 0 81512 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_881
timestamp 1666464484
transform 1 0 82156 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_887
timestamp 1666464484
transform 1 0 82708 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_893
timestamp 1666464484
transform 1 0 83260 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_899
timestamp 1666464484
transform 1 0 83812 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_911
timestamp 1666464484
transform 1 0 84916 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_923
timestamp 1666464484
transform 1 0 86020 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_925
timestamp 1666464484
transform 1 0 86204 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_937
timestamp 1666464484
transform 1 0 87308 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_949
timestamp 1666464484
transform 1 0 88412 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_961
timestamp 1666464484
transform 1 0 89516 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_973
timestamp 1666464484
transform 1 0 90620 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_979
timestamp 1666464484
transform 1 0 91172 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_981
timestamp 1666464484
transform 1 0 91356 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_993
timestamp 1666464484
transform 1 0 92460 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1005
timestamp 1666464484
transform 1 0 93564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1017
timestamp 1666464484
transform 1 0 94668 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1029
timestamp 1666464484
transform 1 0 95772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1035
timestamp 1666464484
transform 1 0 96324 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1037
timestamp 1666464484
transform 1 0 96508 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1049
timestamp 1666464484
transform 1 0 97612 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1061
timestamp 1666464484
transform 1 0 98716 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1073
timestamp 1666464484
transform 1 0 99820 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1085
timestamp 1666464484
transform 1 0 100924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1091
timestamp 1666464484
transform 1 0 101476 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1093
timestamp 1666464484
transform 1 0 101660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1105
timestamp 1666464484
transform 1 0 102764 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1117
timestamp 1666464484
transform 1 0 103868 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1129
timestamp 1666464484
transform 1 0 104972 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1141
timestamp 1666464484
transform 1 0 106076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1147
timestamp 1666464484
transform 1 0 106628 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1149
timestamp 1666464484
transform 1 0 106812 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1161
timestamp 1666464484
transform 1 0 107916 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1173
timestamp 1666464484
transform 1 0 109020 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1185
timestamp 1666464484
transform 1 0 110124 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1197
timestamp 1666464484
transform 1 0 111228 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1203
timestamp 1666464484
transform 1 0 111780 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1205
timestamp 1666464484
transform 1 0 111964 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1217
timestamp 1666464484
transform 1 0 113068 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1229
timestamp 1666464484
transform 1 0 114172 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1241
timestamp 1666464484
transform 1 0 115276 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1253
timestamp 1666464484
transform 1 0 116380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1259
timestamp 1666464484
transform 1 0 116932 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1261
timestamp 1666464484
transform 1 0 117116 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1273
timestamp 1666464484
transform 1 0 118220 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1285
timestamp 1666464484
transform 1 0 119324 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1297
timestamp 1666464484
transform 1 0 120428 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1309
timestamp 1666464484
transform 1 0 121532 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1315
timestamp 1666464484
transform 1 0 122084 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1317
timestamp 1666464484
transform 1 0 122268 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1329
timestamp 1666464484
transform 1 0 123372 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1341
timestamp 1666464484
transform 1 0 124476 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1353
timestamp 1666464484
transform 1 0 125580 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1365
timestamp 1666464484
transform 1 0 126684 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1371
timestamp 1666464484
transform 1 0 127236 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1373
timestamp 1666464484
transform 1 0 127420 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1385
timestamp 1666464484
transform 1 0 128524 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1397
timestamp 1666464484
transform 1 0 129628 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1409
timestamp 1666464484
transform 1 0 130732 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1421
timestamp 1666464484
transform 1 0 131836 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1427
timestamp 1666464484
transform 1 0 132388 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1429
timestamp 1666464484
transform 1 0 132572 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1441
timestamp 1666464484
transform 1 0 133676 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1453
timestamp 1666464484
transform 1 0 134780 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1465
timestamp 1666464484
transform 1 0 135884 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1477
timestamp 1666464484
transform 1 0 136988 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1483
timestamp 1666464484
transform 1 0 137540 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1485
timestamp 1666464484
transform 1 0 137724 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1497
timestamp 1666464484
transform 1 0 138828 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1509
timestamp 1666464484
transform 1 0 139932 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1521
timestamp 1666464484
transform 1 0 141036 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1533
timestamp 1666464484
transform 1 0 142140 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1539
timestamp 1666464484
transform 1 0 142692 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1541
timestamp 1666464484
transform 1 0 142876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1553
timestamp 1666464484
transform 1 0 143980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1565
timestamp 1666464484
transform 1 0 145084 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1577
timestamp 1666464484
transform 1 0 146188 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1589
timestamp 1666464484
transform 1 0 147292 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1595
timestamp 1666464484
transform 1 0 147844 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1597
timestamp 1666464484
transform 1 0 148028 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1666464484
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1666464484
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1666464484
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1666464484
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1666464484
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1666464484
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1666464484
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1666464484
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1666464484
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1666464484
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1666464484
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1666464484
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1666464484
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1666464484
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1666464484
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1666464484
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1666464484
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1666464484
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1666464484
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1666464484
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1666464484
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1666464484
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1666464484
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1666464484
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1666464484
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1666464484
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1666464484
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_293
timestamp 1666464484
transform 1 0 28060 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_298
timestamp 1666464484
transform 1 0 28520 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_310
timestamp 1666464484
transform 1 0 29624 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_322
timestamp 1666464484
transform 1 0 30728 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_334
timestamp 1666464484
transform 1 0 31832 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1666464484
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1666464484
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1666464484
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_373
timestamp 1666464484
transform 1 0 35420 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_376
timestamp 1666464484
transform 1 0 35696 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_382
timestamp 1666464484
transform 1 0 36248 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_386
timestamp 1666464484
transform 1 0 36616 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_389
timestamp 1666464484
transform 1 0 36892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_393
timestamp 1666464484
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_397
timestamp 1666464484
transform 1 0 37628 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_403
timestamp 1666464484
transform 1 0 38180 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_406
timestamp 1666464484
transform 1 0 38456 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_418
timestamp 1666464484
transform 1 0 39560 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_430
timestamp 1666464484
transform 1 0 40664 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_442
timestamp 1666464484
transform 1 0 41768 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_449
timestamp 1666464484
transform 1 0 42412 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_453
timestamp 1666464484
transform 1 0 42780 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_465
timestamp 1666464484
transform 1 0 43884 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_477
timestamp 1666464484
transform 1 0 44988 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_489
timestamp 1666464484
transform 1 0 46092 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_497
timestamp 1666464484
transform 1 0 46828 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_502
timestamp 1666464484
transform 1 0 47288 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_505
timestamp 1666464484
transform 1 0 47564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_509
timestamp 1666464484
transform 1 0 47932 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_512
timestamp 1666464484
transform 1 0 48208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_518
timestamp 1666464484
transform 1 0 48760 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_524
timestamp 1666464484
transform 1 0 49312 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_536
timestamp 1666464484
transform 1 0 50416 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_548
timestamp 1666464484
transform 1 0 51520 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_561
timestamp 1666464484
transform 1 0 52716 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_565
timestamp 1666464484
transform 1 0 53084 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_571
timestamp 1666464484
transform 1 0 53636 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_583
timestamp 1666464484
transform 1 0 54740 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_595
timestamp 1666464484
transform 1 0 55844 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_607
timestamp 1666464484
transform 1 0 56948 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1666464484
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_617
timestamp 1666464484
transform 1 0 57868 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_621
timestamp 1666464484
transform 1 0 58236 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_627
timestamp 1666464484
transform 1 0 58788 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_639
timestamp 1666464484
transform 1 0 59892 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_647
timestamp 1666464484
transform 1 0 60628 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_650
timestamp 1666464484
transform 1 0 60904 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_658
timestamp 1666464484
transform 1 0 61640 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_661
timestamp 1666464484
transform 1 0 61916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_667
timestamp 1666464484
transform 1 0 62468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_670
timestamp 1666464484
transform 1 0 62744 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_673
timestamp 1666464484
transform 1 0 63020 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_679
timestamp 1666464484
transform 1 0 63572 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_682
timestamp 1666464484
transform 1 0 63848 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_688
timestamp 1666464484
transform 1 0 64400 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_694
timestamp 1666464484
transform 1 0 64952 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_700
timestamp 1666464484
transform 1 0 65504 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_706
timestamp 1666464484
transform 1 0 66056 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_712
timestamp 1666464484
transform 1 0 66608 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_718
timestamp 1666464484
transform 1 0 67160 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_726
timestamp 1666464484
transform 1 0 67896 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_729
timestamp 1666464484
transform 1 0 68172 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_733
timestamp 1666464484
transform 1 0 68540 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_739
timestamp 1666464484
transform 1 0 69092 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_743
timestamp 1666464484
transform 1 0 69460 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_746
timestamp 1666464484
transform 1 0 69736 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_752
timestamp 1666464484
transform 1 0 70288 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_758
timestamp 1666464484
transform 1 0 70840 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_770
timestamp 1666464484
transform 1 0 71944 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_782
timestamp 1666464484
transform 1 0 73048 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_785
timestamp 1666464484
transform 1 0 73324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_797
timestamp 1666464484
transform 1 0 74428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_809
timestamp 1666464484
transform 1 0 75532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_821
timestamp 1666464484
transform 1 0 76636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_833
timestamp 1666464484
transform 1 0 77740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_838
timestamp 1666464484
transform 1 0 78200 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_841
timestamp 1666464484
transform 1 0 78476 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_846
timestamp 1666464484
transform 1 0 78936 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_853
timestamp 1666464484
transform 1 0 79580 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_860
timestamp 1666464484
transform 1 0 80224 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_867
timestamp 1666464484
transform 1 0 80868 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_874
timestamp 1666464484
transform 1 0 81512 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_880
timestamp 1666464484
transform 1 0 82064 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_886
timestamp 1666464484
transform 1 0 82616 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_892
timestamp 1666464484
transform 1 0 83168 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_897
timestamp 1666464484
transform 1 0 83628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_909
timestamp 1666464484
transform 1 0 84732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_921
timestamp 1666464484
transform 1 0 85836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_933
timestamp 1666464484
transform 1 0 86940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_945
timestamp 1666464484
transform 1 0 88044 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_951
timestamp 1666464484
transform 1 0 88596 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_953
timestamp 1666464484
transform 1 0 88780 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_965
timestamp 1666464484
transform 1 0 89884 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_977
timestamp 1666464484
transform 1 0 90988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_989
timestamp 1666464484
transform 1 0 92092 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1001
timestamp 1666464484
transform 1 0 93196 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1007
timestamp 1666464484
transform 1 0 93748 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1009
timestamp 1666464484
transform 1 0 93932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1021
timestamp 1666464484
transform 1 0 95036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1033
timestamp 1666464484
transform 1 0 96140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1045
timestamp 1666464484
transform 1 0 97244 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1057
timestamp 1666464484
transform 1 0 98348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1063
timestamp 1666464484
transform 1 0 98900 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1065
timestamp 1666464484
transform 1 0 99084 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1077
timestamp 1666464484
transform 1 0 100188 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1089
timestamp 1666464484
transform 1 0 101292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1101
timestamp 1666464484
transform 1 0 102396 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1113
timestamp 1666464484
transform 1 0 103500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1119
timestamp 1666464484
transform 1 0 104052 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1121
timestamp 1666464484
transform 1 0 104236 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1133
timestamp 1666464484
transform 1 0 105340 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1145
timestamp 1666464484
transform 1 0 106444 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1157
timestamp 1666464484
transform 1 0 107548 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1169
timestamp 1666464484
transform 1 0 108652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1175
timestamp 1666464484
transform 1 0 109204 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1177
timestamp 1666464484
transform 1 0 109388 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1189
timestamp 1666464484
transform 1 0 110492 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1201
timestamp 1666464484
transform 1 0 111596 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1213
timestamp 1666464484
transform 1 0 112700 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1225
timestamp 1666464484
transform 1 0 113804 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1231
timestamp 1666464484
transform 1 0 114356 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1233
timestamp 1666464484
transform 1 0 114540 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1245
timestamp 1666464484
transform 1 0 115644 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1257
timestamp 1666464484
transform 1 0 116748 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1269
timestamp 1666464484
transform 1 0 117852 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1281
timestamp 1666464484
transform 1 0 118956 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1287
timestamp 1666464484
transform 1 0 119508 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1289
timestamp 1666464484
transform 1 0 119692 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1301
timestamp 1666464484
transform 1 0 120796 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1313
timestamp 1666464484
transform 1 0 121900 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1325
timestamp 1666464484
transform 1 0 123004 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1337
timestamp 1666464484
transform 1 0 124108 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1343
timestamp 1666464484
transform 1 0 124660 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1345
timestamp 1666464484
transform 1 0 124844 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1357
timestamp 1666464484
transform 1 0 125948 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1369
timestamp 1666464484
transform 1 0 127052 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1381
timestamp 1666464484
transform 1 0 128156 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1393
timestamp 1666464484
transform 1 0 129260 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1399
timestamp 1666464484
transform 1 0 129812 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1401
timestamp 1666464484
transform 1 0 129996 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1413
timestamp 1666464484
transform 1 0 131100 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1425
timestamp 1666464484
transform 1 0 132204 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1437
timestamp 1666464484
transform 1 0 133308 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1449
timestamp 1666464484
transform 1 0 134412 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1455
timestamp 1666464484
transform 1 0 134964 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1457
timestamp 1666464484
transform 1 0 135148 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1469
timestamp 1666464484
transform 1 0 136252 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1481
timestamp 1666464484
transform 1 0 137356 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1493
timestamp 1666464484
transform 1 0 138460 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1505
timestamp 1666464484
transform 1 0 139564 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1511
timestamp 1666464484
transform 1 0 140116 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1513
timestamp 1666464484
transform 1 0 140300 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1525
timestamp 1666464484
transform 1 0 141404 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1537
timestamp 1666464484
transform 1 0 142508 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1549
timestamp 1666464484
transform 1 0 143612 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1561
timestamp 1666464484
transform 1 0 144716 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1567
timestamp 1666464484
transform 1 0 145268 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1569
timestamp 1666464484
transform 1 0 145452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1581
timestamp 1666464484
transform 1 0 146556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1593
timestamp 1666464484
transform 1 0 147660 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1601
timestamp 1666464484
transform 1 0 148396 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1666464484
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1666464484
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1666464484
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1666464484
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1666464484
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1666464484
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1666464484
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1666464484
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1666464484
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1666464484
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1666464484
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1666464484
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1666464484
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1666464484
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1666464484
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1666464484
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1666464484
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1666464484
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1666464484
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1666464484
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1666464484
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1666464484
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1666464484
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1666464484
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1666464484
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1666464484
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1666464484
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1666464484
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1666464484
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1666464484
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1666464484
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1666464484
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1666464484
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1666464484
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1666464484
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1666464484
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1666464484
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1666464484
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1666464484
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1666464484
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1666464484
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1666464484
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1666464484
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1666464484
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1666464484
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1666464484
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1666464484
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1666464484
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1666464484
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1666464484
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1666464484
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1666464484
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1666464484
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1666464484
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1666464484
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1666464484
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1666464484
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1666464484
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1666464484
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1666464484
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1666464484
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1666464484
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_625
timestamp 1666464484
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1666464484
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1666464484
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1666464484
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1666464484
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_669
timestamp 1666464484
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_681
timestamp 1666464484
transform 1 0 63756 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_686
timestamp 1666464484
transform 1 0 64216 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_694
timestamp 1666464484
transform 1 0 64952 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_697
timestamp 1666464484
transform 1 0 65228 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_701
timestamp 1666464484
transform 1 0 65596 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_705
timestamp 1666464484
transform 1 0 65964 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_717
timestamp 1666464484
transform 1 0 67068 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_729
timestamp 1666464484
transform 1 0 68172 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_741
timestamp 1666464484
transform 1 0 69276 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_744
timestamp 1666464484
transform 1 0 69552 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_757
timestamp 1666464484
transform 1 0 70748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_769
timestamp 1666464484
transform 1 0 71852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_781
timestamp 1666464484
transform 1 0 72956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_793
timestamp 1666464484
transform 1 0 74060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_805
timestamp 1666464484
transform 1 0 75164 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_811
timestamp 1666464484
transform 1 0 75716 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_813
timestamp 1666464484
transform 1 0 75900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_825
timestamp 1666464484
transform 1 0 77004 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_837
timestamp 1666464484
transform 1 0 78108 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_845
timestamp 1666464484
transform 1 0 78844 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_848
timestamp 1666464484
transform 1 0 79120 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_854
timestamp 1666464484
transform 1 0 79672 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_860
timestamp 1666464484
transform 1 0 80224 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_866
timestamp 1666464484
transform 1 0 80776 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_869
timestamp 1666464484
transform 1 0 81052 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_881
timestamp 1666464484
transform 1 0 82156 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_893
timestamp 1666464484
transform 1 0 83260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_905
timestamp 1666464484
transform 1 0 84364 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_917
timestamp 1666464484
transform 1 0 85468 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_923
timestamp 1666464484
transform 1 0 86020 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_925
timestamp 1666464484
transform 1 0 86204 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_937
timestamp 1666464484
transform 1 0 87308 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_949
timestamp 1666464484
transform 1 0 88412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_961
timestamp 1666464484
transform 1 0 89516 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_973
timestamp 1666464484
transform 1 0 90620 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_979
timestamp 1666464484
transform 1 0 91172 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_981
timestamp 1666464484
transform 1 0 91356 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_993
timestamp 1666464484
transform 1 0 92460 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1005
timestamp 1666464484
transform 1 0 93564 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1017
timestamp 1666464484
transform 1 0 94668 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1029
timestamp 1666464484
transform 1 0 95772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1035
timestamp 1666464484
transform 1 0 96324 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1037
timestamp 1666464484
transform 1 0 96508 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1049
timestamp 1666464484
transform 1 0 97612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1061
timestamp 1666464484
transform 1 0 98716 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1073
timestamp 1666464484
transform 1 0 99820 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1085
timestamp 1666464484
transform 1 0 100924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1091
timestamp 1666464484
transform 1 0 101476 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1093
timestamp 1666464484
transform 1 0 101660 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1105
timestamp 1666464484
transform 1 0 102764 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1117
timestamp 1666464484
transform 1 0 103868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1129
timestamp 1666464484
transform 1 0 104972 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1141
timestamp 1666464484
transform 1 0 106076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1147
timestamp 1666464484
transform 1 0 106628 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1149
timestamp 1666464484
transform 1 0 106812 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1161
timestamp 1666464484
transform 1 0 107916 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1173
timestamp 1666464484
transform 1 0 109020 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1185
timestamp 1666464484
transform 1 0 110124 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1197
timestamp 1666464484
transform 1 0 111228 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1203
timestamp 1666464484
transform 1 0 111780 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1205
timestamp 1666464484
transform 1 0 111964 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1217
timestamp 1666464484
transform 1 0 113068 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1229
timestamp 1666464484
transform 1 0 114172 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1241
timestamp 1666464484
transform 1 0 115276 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1253
timestamp 1666464484
transform 1 0 116380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1259
timestamp 1666464484
transform 1 0 116932 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1261
timestamp 1666464484
transform 1 0 117116 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1273
timestamp 1666464484
transform 1 0 118220 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1285
timestamp 1666464484
transform 1 0 119324 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1297
timestamp 1666464484
transform 1 0 120428 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1309
timestamp 1666464484
transform 1 0 121532 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1315
timestamp 1666464484
transform 1 0 122084 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1317
timestamp 1666464484
transform 1 0 122268 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1329
timestamp 1666464484
transform 1 0 123372 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1341
timestamp 1666464484
transform 1 0 124476 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1353
timestamp 1666464484
transform 1 0 125580 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1365
timestamp 1666464484
transform 1 0 126684 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1371
timestamp 1666464484
transform 1 0 127236 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1373
timestamp 1666464484
transform 1 0 127420 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1385
timestamp 1666464484
transform 1 0 128524 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1397
timestamp 1666464484
transform 1 0 129628 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1409
timestamp 1666464484
transform 1 0 130732 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1421
timestamp 1666464484
transform 1 0 131836 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1427
timestamp 1666464484
transform 1 0 132388 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1429
timestamp 1666464484
transform 1 0 132572 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1441
timestamp 1666464484
transform 1 0 133676 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1453
timestamp 1666464484
transform 1 0 134780 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1465
timestamp 1666464484
transform 1 0 135884 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1477
timestamp 1666464484
transform 1 0 136988 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1483
timestamp 1666464484
transform 1 0 137540 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1485
timestamp 1666464484
transform 1 0 137724 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1497
timestamp 1666464484
transform 1 0 138828 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1509
timestamp 1666464484
transform 1 0 139932 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1521
timestamp 1666464484
transform 1 0 141036 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1533
timestamp 1666464484
transform 1 0 142140 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1539
timestamp 1666464484
transform 1 0 142692 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1541
timestamp 1666464484
transform 1 0 142876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1553
timestamp 1666464484
transform 1 0 143980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1565
timestamp 1666464484
transform 1 0 145084 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1577
timestamp 1666464484
transform 1 0 146188 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1589
timestamp 1666464484
transform 1 0 147292 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1595
timestamp 1666464484
transform 1 0 147844 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1597
timestamp 1666464484
transform 1 0 148028 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1666464484
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1666464484
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1666464484
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1666464484
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1666464484
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1666464484
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1666464484
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1666464484
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1666464484
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1666464484
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1666464484
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1666464484
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1666464484
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1666464484
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1666464484
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1666464484
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1666464484
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1666464484
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1666464484
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1666464484
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1666464484
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1666464484
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1666464484
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1666464484
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1666464484
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1666464484
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1666464484
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1666464484
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1666464484
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1666464484
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1666464484
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1666464484
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1666464484
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1666464484
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1666464484
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1666464484
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1666464484
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1666464484
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1666464484
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1666464484
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1666464484
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1666464484
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1666464484
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1666464484
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1666464484
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1666464484
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1666464484
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1666464484
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1666464484
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1666464484
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1666464484
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1666464484
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1666464484
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1666464484
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1666464484
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1666464484
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1666464484
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1666464484
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1666464484
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1666464484
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1666464484
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1666464484
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_617
timestamp 1666464484
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_629
timestamp 1666464484
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_641
timestamp 1666464484
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_653
timestamp 1666464484
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1666464484
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1666464484
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_673
timestamp 1666464484
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_685
timestamp 1666464484
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_697
timestamp 1666464484
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_709
timestamp 1666464484
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1666464484
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1666464484
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_729
timestamp 1666464484
transform 1 0 68172 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_741
timestamp 1666464484
transform 1 0 69276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_753
timestamp 1666464484
transform 1 0 70380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_765
timestamp 1666464484
transform 1 0 71484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_777
timestamp 1666464484
transform 1 0 72588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_783
timestamp 1666464484
transform 1 0 73140 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_785
timestamp 1666464484
transform 1 0 73324 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_797
timestamp 1666464484
transform 1 0 74428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_809
timestamp 1666464484
transform 1 0 75532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_821
timestamp 1666464484
transform 1 0 76636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_833
timestamp 1666464484
transform 1 0 77740 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_839
timestamp 1666464484
transform 1 0 78292 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_841
timestamp 1666464484
transform 1 0 78476 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_853
timestamp 1666464484
transform 1 0 79580 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_865
timestamp 1666464484
transform 1 0 80684 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_877
timestamp 1666464484
transform 1 0 81788 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_889
timestamp 1666464484
transform 1 0 82892 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_895
timestamp 1666464484
transform 1 0 83444 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_897
timestamp 1666464484
transform 1 0 83628 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_909
timestamp 1666464484
transform 1 0 84732 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_921
timestamp 1666464484
transform 1 0 85836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_933
timestamp 1666464484
transform 1 0 86940 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_945
timestamp 1666464484
transform 1 0 88044 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_951
timestamp 1666464484
transform 1 0 88596 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_953
timestamp 1666464484
transform 1 0 88780 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_965
timestamp 1666464484
transform 1 0 89884 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_977
timestamp 1666464484
transform 1 0 90988 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_989
timestamp 1666464484
transform 1 0 92092 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1001
timestamp 1666464484
transform 1 0 93196 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1007
timestamp 1666464484
transform 1 0 93748 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1009
timestamp 1666464484
transform 1 0 93932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1021
timestamp 1666464484
transform 1 0 95036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1033
timestamp 1666464484
transform 1 0 96140 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1045
timestamp 1666464484
transform 1 0 97244 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1057
timestamp 1666464484
transform 1 0 98348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1063
timestamp 1666464484
transform 1 0 98900 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1065
timestamp 1666464484
transform 1 0 99084 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1077
timestamp 1666464484
transform 1 0 100188 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1089
timestamp 1666464484
transform 1 0 101292 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1101
timestamp 1666464484
transform 1 0 102396 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1113
timestamp 1666464484
transform 1 0 103500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1119
timestamp 1666464484
transform 1 0 104052 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1121
timestamp 1666464484
transform 1 0 104236 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1133
timestamp 1666464484
transform 1 0 105340 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1145
timestamp 1666464484
transform 1 0 106444 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1157
timestamp 1666464484
transform 1 0 107548 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1169
timestamp 1666464484
transform 1 0 108652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1175
timestamp 1666464484
transform 1 0 109204 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1177
timestamp 1666464484
transform 1 0 109388 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1189
timestamp 1666464484
transform 1 0 110492 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1201
timestamp 1666464484
transform 1 0 111596 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1213
timestamp 1666464484
transform 1 0 112700 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1225
timestamp 1666464484
transform 1 0 113804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1231
timestamp 1666464484
transform 1 0 114356 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1233
timestamp 1666464484
transform 1 0 114540 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1245
timestamp 1666464484
transform 1 0 115644 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1257
timestamp 1666464484
transform 1 0 116748 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1269
timestamp 1666464484
transform 1 0 117852 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1281
timestamp 1666464484
transform 1 0 118956 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1287
timestamp 1666464484
transform 1 0 119508 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1289
timestamp 1666464484
transform 1 0 119692 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1301
timestamp 1666464484
transform 1 0 120796 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1313
timestamp 1666464484
transform 1 0 121900 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1325
timestamp 1666464484
transform 1 0 123004 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1337
timestamp 1666464484
transform 1 0 124108 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1343
timestamp 1666464484
transform 1 0 124660 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1345
timestamp 1666464484
transform 1 0 124844 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1357
timestamp 1666464484
transform 1 0 125948 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1369
timestamp 1666464484
transform 1 0 127052 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1381
timestamp 1666464484
transform 1 0 128156 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1393
timestamp 1666464484
transform 1 0 129260 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1399
timestamp 1666464484
transform 1 0 129812 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1401
timestamp 1666464484
transform 1 0 129996 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1413
timestamp 1666464484
transform 1 0 131100 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1425
timestamp 1666464484
transform 1 0 132204 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1437
timestamp 1666464484
transform 1 0 133308 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1449
timestamp 1666464484
transform 1 0 134412 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1455
timestamp 1666464484
transform 1 0 134964 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1457
timestamp 1666464484
transform 1 0 135148 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1469
timestamp 1666464484
transform 1 0 136252 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1481
timestamp 1666464484
transform 1 0 137356 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1493
timestamp 1666464484
transform 1 0 138460 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1505
timestamp 1666464484
transform 1 0 139564 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1511
timestamp 1666464484
transform 1 0 140116 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1513
timestamp 1666464484
transform 1 0 140300 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1525
timestamp 1666464484
transform 1 0 141404 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1537
timestamp 1666464484
transform 1 0 142508 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1549
timestamp 1666464484
transform 1 0 143612 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1561
timestamp 1666464484
transform 1 0 144716 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1567
timestamp 1666464484
transform 1 0 145268 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1569
timestamp 1666464484
transform 1 0 145452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1581
timestamp 1666464484
transform 1 0 146556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1593
timestamp 1666464484
transform 1 0 147660 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1601
timestamp 1666464484
transform 1 0 148396 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1666464484
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1666464484
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1666464484
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1666464484
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1666464484
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1666464484
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1666464484
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1666464484
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1666464484
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1666464484
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1666464484
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1666464484
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1666464484
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1666464484
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1666464484
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1666464484
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1666464484
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1666464484
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1666464484
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1666464484
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1666464484
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1666464484
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1666464484
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1666464484
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1666464484
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1666464484
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1666464484
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1666464484
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1666464484
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1666464484
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1666464484
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1666464484
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1666464484
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1666464484
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1666464484
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1666464484
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1666464484
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1666464484
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1666464484
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1666464484
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1666464484
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1666464484
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1666464484
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1666464484
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1666464484
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1666464484
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1666464484
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1666464484
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1666464484
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1666464484
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1666464484
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1666464484
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1666464484
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1666464484
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1666464484
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1666464484
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1666464484
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1666464484
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1666464484
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1666464484
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1666464484
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1666464484
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_625
timestamp 1666464484
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1666464484
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1666464484
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_645
timestamp 1666464484
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_657
timestamp 1666464484
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_669
timestamp 1666464484
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_681
timestamp 1666464484
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1666464484
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1666464484
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_701
timestamp 1666464484
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_713
timestamp 1666464484
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_725
timestamp 1666464484
transform 1 0 67804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_737
timestamp 1666464484
transform 1 0 68908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_749
timestamp 1666464484
transform 1 0 70012 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_755
timestamp 1666464484
transform 1 0 70564 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_757
timestamp 1666464484
transform 1 0 70748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_769
timestamp 1666464484
transform 1 0 71852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_781
timestamp 1666464484
transform 1 0 72956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_793
timestamp 1666464484
transform 1 0 74060 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_805
timestamp 1666464484
transform 1 0 75164 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_811
timestamp 1666464484
transform 1 0 75716 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_813
timestamp 1666464484
transform 1 0 75900 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_825
timestamp 1666464484
transform 1 0 77004 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_837
timestamp 1666464484
transform 1 0 78108 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_849
timestamp 1666464484
transform 1 0 79212 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_861
timestamp 1666464484
transform 1 0 80316 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_867
timestamp 1666464484
transform 1 0 80868 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_869
timestamp 1666464484
transform 1 0 81052 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_881
timestamp 1666464484
transform 1 0 82156 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_893
timestamp 1666464484
transform 1 0 83260 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_905
timestamp 1666464484
transform 1 0 84364 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_917
timestamp 1666464484
transform 1 0 85468 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_923
timestamp 1666464484
transform 1 0 86020 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_925
timestamp 1666464484
transform 1 0 86204 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_937
timestamp 1666464484
transform 1 0 87308 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_949
timestamp 1666464484
transform 1 0 88412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_961
timestamp 1666464484
transform 1 0 89516 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_973
timestamp 1666464484
transform 1 0 90620 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_979
timestamp 1666464484
transform 1 0 91172 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_981
timestamp 1666464484
transform 1 0 91356 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_993
timestamp 1666464484
transform 1 0 92460 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1005
timestamp 1666464484
transform 1 0 93564 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1017
timestamp 1666464484
transform 1 0 94668 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1029
timestamp 1666464484
transform 1 0 95772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1035
timestamp 1666464484
transform 1 0 96324 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1037
timestamp 1666464484
transform 1 0 96508 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1049
timestamp 1666464484
transform 1 0 97612 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1061
timestamp 1666464484
transform 1 0 98716 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1073
timestamp 1666464484
transform 1 0 99820 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1085
timestamp 1666464484
transform 1 0 100924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1091
timestamp 1666464484
transform 1 0 101476 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1093
timestamp 1666464484
transform 1 0 101660 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1105
timestamp 1666464484
transform 1 0 102764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1117
timestamp 1666464484
transform 1 0 103868 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1129
timestamp 1666464484
transform 1 0 104972 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1141
timestamp 1666464484
transform 1 0 106076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1147
timestamp 1666464484
transform 1 0 106628 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1149
timestamp 1666464484
transform 1 0 106812 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1161
timestamp 1666464484
transform 1 0 107916 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1173
timestamp 1666464484
transform 1 0 109020 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1185
timestamp 1666464484
transform 1 0 110124 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1197
timestamp 1666464484
transform 1 0 111228 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1203
timestamp 1666464484
transform 1 0 111780 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1205
timestamp 1666464484
transform 1 0 111964 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1217
timestamp 1666464484
transform 1 0 113068 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1229
timestamp 1666464484
transform 1 0 114172 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1241
timestamp 1666464484
transform 1 0 115276 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1253
timestamp 1666464484
transform 1 0 116380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1259
timestamp 1666464484
transform 1 0 116932 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1261
timestamp 1666464484
transform 1 0 117116 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1273
timestamp 1666464484
transform 1 0 118220 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1285
timestamp 1666464484
transform 1 0 119324 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1297
timestamp 1666464484
transform 1 0 120428 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1309
timestamp 1666464484
transform 1 0 121532 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1315
timestamp 1666464484
transform 1 0 122084 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1317
timestamp 1666464484
transform 1 0 122268 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1329
timestamp 1666464484
transform 1 0 123372 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1341
timestamp 1666464484
transform 1 0 124476 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1353
timestamp 1666464484
transform 1 0 125580 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1365
timestamp 1666464484
transform 1 0 126684 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1371
timestamp 1666464484
transform 1 0 127236 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1373
timestamp 1666464484
transform 1 0 127420 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1385
timestamp 1666464484
transform 1 0 128524 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1397
timestamp 1666464484
transform 1 0 129628 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1409
timestamp 1666464484
transform 1 0 130732 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1421
timestamp 1666464484
transform 1 0 131836 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1427
timestamp 1666464484
transform 1 0 132388 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1429
timestamp 1666464484
transform 1 0 132572 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1441
timestamp 1666464484
transform 1 0 133676 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1453
timestamp 1666464484
transform 1 0 134780 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1465
timestamp 1666464484
transform 1 0 135884 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1477
timestamp 1666464484
transform 1 0 136988 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1483
timestamp 1666464484
transform 1 0 137540 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1485
timestamp 1666464484
transform 1 0 137724 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1497
timestamp 1666464484
transform 1 0 138828 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1509
timestamp 1666464484
transform 1 0 139932 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1521
timestamp 1666464484
transform 1 0 141036 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1533
timestamp 1666464484
transform 1 0 142140 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1539
timestamp 1666464484
transform 1 0 142692 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1541
timestamp 1666464484
transform 1 0 142876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1553
timestamp 1666464484
transform 1 0 143980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1565
timestamp 1666464484
transform 1 0 145084 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1577
timestamp 1666464484
transform 1 0 146188 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1589
timestamp 1666464484
transform 1 0 147292 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1595
timestamp 1666464484
transform 1 0 147844 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1597
timestamp 1666464484
transform 1 0 148028 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1666464484
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1666464484
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1666464484
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1666464484
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1666464484
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1666464484
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1666464484
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1666464484
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1666464484
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1666464484
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1666464484
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1666464484
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1666464484
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1666464484
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1666464484
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1666464484
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1666464484
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1666464484
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1666464484
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1666464484
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1666464484
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1666464484
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1666464484
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1666464484
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1666464484
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1666464484
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1666464484
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1666464484
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1666464484
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1666464484
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1666464484
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1666464484
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1666464484
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1666464484
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1666464484
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1666464484
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1666464484
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1666464484
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1666464484
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1666464484
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1666464484
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1666464484
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1666464484
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1666464484
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1666464484
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1666464484
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1666464484
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1666464484
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1666464484
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1666464484
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1666464484
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1666464484
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1666464484
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1666464484
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1666464484
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1666464484
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1666464484
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1666464484
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1666464484
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1666464484
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1666464484
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1666464484
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_617
timestamp 1666464484
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_629
timestamp 1666464484
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_641
timestamp 1666464484
transform 1 0 60076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_653
timestamp 1666464484
transform 1 0 61180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_665
timestamp 1666464484
transform 1 0 62284 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_671
timestamp 1666464484
transform 1 0 62836 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_673
timestamp 1666464484
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_685
timestamp 1666464484
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_697
timestamp 1666464484
transform 1 0 65228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_709
timestamp 1666464484
transform 1 0 66332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_721
timestamp 1666464484
transform 1 0 67436 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_727
timestamp 1666464484
transform 1 0 67988 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_729
timestamp 1666464484
transform 1 0 68172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_741
timestamp 1666464484
transform 1 0 69276 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_753
timestamp 1666464484
transform 1 0 70380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_765
timestamp 1666464484
transform 1 0 71484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_777
timestamp 1666464484
transform 1 0 72588 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_783
timestamp 1666464484
transform 1 0 73140 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_785
timestamp 1666464484
transform 1 0 73324 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_797
timestamp 1666464484
transform 1 0 74428 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_809
timestamp 1666464484
transform 1 0 75532 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_821
timestamp 1666464484
transform 1 0 76636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_833
timestamp 1666464484
transform 1 0 77740 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_839
timestamp 1666464484
transform 1 0 78292 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_841
timestamp 1666464484
transform 1 0 78476 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_853
timestamp 1666464484
transform 1 0 79580 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_865
timestamp 1666464484
transform 1 0 80684 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_877
timestamp 1666464484
transform 1 0 81788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_889
timestamp 1666464484
transform 1 0 82892 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_895
timestamp 1666464484
transform 1 0 83444 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_897
timestamp 1666464484
transform 1 0 83628 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_909
timestamp 1666464484
transform 1 0 84732 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_921
timestamp 1666464484
transform 1 0 85836 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_933
timestamp 1666464484
transform 1 0 86940 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_945
timestamp 1666464484
transform 1 0 88044 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_951
timestamp 1666464484
transform 1 0 88596 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_953
timestamp 1666464484
transform 1 0 88780 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_965
timestamp 1666464484
transform 1 0 89884 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_977
timestamp 1666464484
transform 1 0 90988 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_989
timestamp 1666464484
transform 1 0 92092 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1001
timestamp 1666464484
transform 1 0 93196 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1007
timestamp 1666464484
transform 1 0 93748 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1009
timestamp 1666464484
transform 1 0 93932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1021
timestamp 1666464484
transform 1 0 95036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1033
timestamp 1666464484
transform 1 0 96140 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1045
timestamp 1666464484
transform 1 0 97244 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1057
timestamp 1666464484
transform 1 0 98348 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1063
timestamp 1666464484
transform 1 0 98900 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1065
timestamp 1666464484
transform 1 0 99084 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1077
timestamp 1666464484
transform 1 0 100188 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1089
timestamp 1666464484
transform 1 0 101292 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1101
timestamp 1666464484
transform 1 0 102396 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1113
timestamp 1666464484
transform 1 0 103500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1119
timestamp 1666464484
transform 1 0 104052 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1121
timestamp 1666464484
transform 1 0 104236 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1133
timestamp 1666464484
transform 1 0 105340 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1145
timestamp 1666464484
transform 1 0 106444 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1157
timestamp 1666464484
transform 1 0 107548 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1169
timestamp 1666464484
transform 1 0 108652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1175
timestamp 1666464484
transform 1 0 109204 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1177
timestamp 1666464484
transform 1 0 109388 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1189
timestamp 1666464484
transform 1 0 110492 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1201
timestamp 1666464484
transform 1 0 111596 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1213
timestamp 1666464484
transform 1 0 112700 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1225
timestamp 1666464484
transform 1 0 113804 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1231
timestamp 1666464484
transform 1 0 114356 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1233
timestamp 1666464484
transform 1 0 114540 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1245
timestamp 1666464484
transform 1 0 115644 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1257
timestamp 1666464484
transform 1 0 116748 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1269
timestamp 1666464484
transform 1 0 117852 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1281
timestamp 1666464484
transform 1 0 118956 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1287
timestamp 1666464484
transform 1 0 119508 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1289
timestamp 1666464484
transform 1 0 119692 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1301
timestamp 1666464484
transform 1 0 120796 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1313
timestamp 1666464484
transform 1 0 121900 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1325
timestamp 1666464484
transform 1 0 123004 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1337
timestamp 1666464484
transform 1 0 124108 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1343
timestamp 1666464484
transform 1 0 124660 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1345
timestamp 1666464484
transform 1 0 124844 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1357
timestamp 1666464484
transform 1 0 125948 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1369
timestamp 1666464484
transform 1 0 127052 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1381
timestamp 1666464484
transform 1 0 128156 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1393
timestamp 1666464484
transform 1 0 129260 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1399
timestamp 1666464484
transform 1 0 129812 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1401
timestamp 1666464484
transform 1 0 129996 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1413
timestamp 1666464484
transform 1 0 131100 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1425
timestamp 1666464484
transform 1 0 132204 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1437
timestamp 1666464484
transform 1 0 133308 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1449
timestamp 1666464484
transform 1 0 134412 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1455
timestamp 1666464484
transform 1 0 134964 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1457
timestamp 1666464484
transform 1 0 135148 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1469
timestamp 1666464484
transform 1 0 136252 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1481
timestamp 1666464484
transform 1 0 137356 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1493
timestamp 1666464484
transform 1 0 138460 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1505
timestamp 1666464484
transform 1 0 139564 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1511
timestamp 1666464484
transform 1 0 140116 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1513
timestamp 1666464484
transform 1 0 140300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1525
timestamp 1666464484
transform 1 0 141404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1537
timestamp 1666464484
transform 1 0 142508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1549
timestamp 1666464484
transform 1 0 143612 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1561
timestamp 1666464484
transform 1 0 144716 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1567
timestamp 1666464484
transform 1 0 145268 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1569
timestamp 1666464484
transform 1 0 145452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1581
timestamp 1666464484
transform 1 0 146556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1593
timestamp 1666464484
transform 1 0 147660 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1601
timestamp 1666464484
transform 1 0 148396 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1666464484
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1666464484
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1666464484
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1666464484
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1666464484
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1666464484
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1666464484
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1666464484
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1666464484
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1666464484
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1666464484
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1666464484
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1666464484
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1666464484
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1666464484
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1666464484
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1666464484
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1666464484
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1666464484
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1666464484
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1666464484
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1666464484
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1666464484
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1666464484
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1666464484
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1666464484
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1666464484
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1666464484
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1666464484
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1666464484
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1666464484
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1666464484
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1666464484
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1666464484
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1666464484
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1666464484
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1666464484
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1666464484
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1666464484
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1666464484
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1666464484
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1666464484
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1666464484
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1666464484
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1666464484
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1666464484
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1666464484
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1666464484
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1666464484
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1666464484
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1666464484
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1666464484
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1666464484
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1666464484
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1666464484
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1666464484
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1666464484
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1666464484
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1666464484
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1666464484
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_601
timestamp 1666464484
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_613
timestamp 1666464484
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_625
timestamp 1666464484
transform 1 0 58604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_637
timestamp 1666464484
transform 1 0 59708 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_643
timestamp 1666464484
transform 1 0 60260 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_645
timestamp 1666464484
transform 1 0 60444 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_657
timestamp 1666464484
transform 1 0 61548 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_669
timestamp 1666464484
transform 1 0 62652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_681
timestamp 1666464484
transform 1 0 63756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_693
timestamp 1666464484
transform 1 0 64860 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_699
timestamp 1666464484
transform 1 0 65412 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_701
timestamp 1666464484
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_713
timestamp 1666464484
transform 1 0 66700 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_725
timestamp 1666464484
transform 1 0 67804 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_737
timestamp 1666464484
transform 1 0 68908 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_749
timestamp 1666464484
transform 1 0 70012 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_755
timestamp 1666464484
transform 1 0 70564 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_757
timestamp 1666464484
transform 1 0 70748 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_769
timestamp 1666464484
transform 1 0 71852 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_781
timestamp 1666464484
transform 1 0 72956 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_793
timestamp 1666464484
transform 1 0 74060 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_805
timestamp 1666464484
transform 1 0 75164 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_811
timestamp 1666464484
transform 1 0 75716 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_813
timestamp 1666464484
transform 1 0 75900 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_825
timestamp 1666464484
transform 1 0 77004 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_837
timestamp 1666464484
transform 1 0 78108 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_849
timestamp 1666464484
transform 1 0 79212 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_861
timestamp 1666464484
transform 1 0 80316 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_867
timestamp 1666464484
transform 1 0 80868 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_869
timestamp 1666464484
transform 1 0 81052 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_881
timestamp 1666464484
transform 1 0 82156 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_893
timestamp 1666464484
transform 1 0 83260 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_905
timestamp 1666464484
transform 1 0 84364 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_917
timestamp 1666464484
transform 1 0 85468 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_923
timestamp 1666464484
transform 1 0 86020 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_925
timestamp 1666464484
transform 1 0 86204 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_937
timestamp 1666464484
transform 1 0 87308 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_949
timestamp 1666464484
transform 1 0 88412 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_961
timestamp 1666464484
transform 1 0 89516 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_973
timestamp 1666464484
transform 1 0 90620 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_979
timestamp 1666464484
transform 1 0 91172 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_981
timestamp 1666464484
transform 1 0 91356 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_993
timestamp 1666464484
transform 1 0 92460 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1005
timestamp 1666464484
transform 1 0 93564 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1017
timestamp 1666464484
transform 1 0 94668 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1029
timestamp 1666464484
transform 1 0 95772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1035
timestamp 1666464484
transform 1 0 96324 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1037
timestamp 1666464484
transform 1 0 96508 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1049
timestamp 1666464484
transform 1 0 97612 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1061
timestamp 1666464484
transform 1 0 98716 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1073
timestamp 1666464484
transform 1 0 99820 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1085
timestamp 1666464484
transform 1 0 100924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1091
timestamp 1666464484
transform 1 0 101476 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1093
timestamp 1666464484
transform 1 0 101660 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1105
timestamp 1666464484
transform 1 0 102764 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1117
timestamp 1666464484
transform 1 0 103868 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1129
timestamp 1666464484
transform 1 0 104972 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1141
timestamp 1666464484
transform 1 0 106076 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1147
timestamp 1666464484
transform 1 0 106628 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1149
timestamp 1666464484
transform 1 0 106812 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1161
timestamp 1666464484
transform 1 0 107916 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1173
timestamp 1666464484
transform 1 0 109020 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1185
timestamp 1666464484
transform 1 0 110124 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1197
timestamp 1666464484
transform 1 0 111228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1203
timestamp 1666464484
transform 1 0 111780 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1205
timestamp 1666464484
transform 1 0 111964 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1217
timestamp 1666464484
transform 1 0 113068 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1229
timestamp 1666464484
transform 1 0 114172 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1241
timestamp 1666464484
transform 1 0 115276 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1253
timestamp 1666464484
transform 1 0 116380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1259
timestamp 1666464484
transform 1 0 116932 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1261
timestamp 1666464484
transform 1 0 117116 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1273
timestamp 1666464484
transform 1 0 118220 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1285
timestamp 1666464484
transform 1 0 119324 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1297
timestamp 1666464484
transform 1 0 120428 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1309
timestamp 1666464484
transform 1 0 121532 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1315
timestamp 1666464484
transform 1 0 122084 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1317
timestamp 1666464484
transform 1 0 122268 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1329
timestamp 1666464484
transform 1 0 123372 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1341
timestamp 1666464484
transform 1 0 124476 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1353
timestamp 1666464484
transform 1 0 125580 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1365
timestamp 1666464484
transform 1 0 126684 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1371
timestamp 1666464484
transform 1 0 127236 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1373
timestamp 1666464484
transform 1 0 127420 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1385
timestamp 1666464484
transform 1 0 128524 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1397
timestamp 1666464484
transform 1 0 129628 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1409
timestamp 1666464484
transform 1 0 130732 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1421
timestamp 1666464484
transform 1 0 131836 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1427
timestamp 1666464484
transform 1 0 132388 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1429
timestamp 1666464484
transform 1 0 132572 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1441
timestamp 1666464484
transform 1 0 133676 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1453
timestamp 1666464484
transform 1 0 134780 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1465
timestamp 1666464484
transform 1 0 135884 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1477
timestamp 1666464484
transform 1 0 136988 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1483
timestamp 1666464484
transform 1 0 137540 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1485
timestamp 1666464484
transform 1 0 137724 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1497
timestamp 1666464484
transform 1 0 138828 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1509
timestamp 1666464484
transform 1 0 139932 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1521
timestamp 1666464484
transform 1 0 141036 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1533
timestamp 1666464484
transform 1 0 142140 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1539
timestamp 1666464484
transform 1 0 142692 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1541
timestamp 1666464484
transform 1 0 142876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1553
timestamp 1666464484
transform 1 0 143980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1565
timestamp 1666464484
transform 1 0 145084 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1577
timestamp 1666464484
transform 1 0 146188 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1589
timestamp 1666464484
transform 1 0 147292 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1595
timestamp 1666464484
transform 1 0 147844 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1597
timestamp 1666464484
transform 1 0 148028 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1666464484
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1666464484
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1666464484
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1666464484
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1666464484
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1666464484
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1666464484
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1666464484
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1666464484
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1666464484
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1666464484
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1666464484
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1666464484
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1666464484
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1666464484
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1666464484
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1666464484
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1666464484
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1666464484
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1666464484
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1666464484
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1666464484
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1666464484
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1666464484
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1666464484
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1666464484
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1666464484
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1666464484
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1666464484
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1666464484
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1666464484
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1666464484
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1666464484
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1666464484
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1666464484
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1666464484
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1666464484
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1666464484
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1666464484
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1666464484
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1666464484
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1666464484
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1666464484
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1666464484
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1666464484
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1666464484
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1666464484
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1666464484
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1666464484
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1666464484
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1666464484
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1666464484
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1666464484
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1666464484
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1666464484
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1666464484
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1666464484
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1666464484
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1666464484
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1666464484
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_597
timestamp 1666464484
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1666464484
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1666464484
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_617
timestamp 1666464484
transform 1 0 57868 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_629
timestamp 1666464484
transform 1 0 58972 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_641
timestamp 1666464484
transform 1 0 60076 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_653
timestamp 1666464484
transform 1 0 61180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_665
timestamp 1666464484
transform 1 0 62284 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_671
timestamp 1666464484
transform 1 0 62836 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_673
timestamp 1666464484
transform 1 0 63020 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_685
timestamp 1666464484
transform 1 0 64124 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_697
timestamp 1666464484
transform 1 0 65228 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_709
timestamp 1666464484
transform 1 0 66332 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_721
timestamp 1666464484
transform 1 0 67436 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_727
timestamp 1666464484
transform 1 0 67988 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_729
timestamp 1666464484
transform 1 0 68172 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_741
timestamp 1666464484
transform 1 0 69276 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_753
timestamp 1666464484
transform 1 0 70380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_765
timestamp 1666464484
transform 1 0 71484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_777
timestamp 1666464484
transform 1 0 72588 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_783
timestamp 1666464484
transform 1 0 73140 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_785
timestamp 1666464484
transform 1 0 73324 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_797
timestamp 1666464484
transform 1 0 74428 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_809
timestamp 1666464484
transform 1 0 75532 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_821
timestamp 1666464484
transform 1 0 76636 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_833
timestamp 1666464484
transform 1 0 77740 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_839
timestamp 1666464484
transform 1 0 78292 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_841
timestamp 1666464484
transform 1 0 78476 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_853
timestamp 1666464484
transform 1 0 79580 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_865
timestamp 1666464484
transform 1 0 80684 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_877
timestamp 1666464484
transform 1 0 81788 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_889
timestamp 1666464484
transform 1 0 82892 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_895
timestamp 1666464484
transform 1 0 83444 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_897
timestamp 1666464484
transform 1 0 83628 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_909
timestamp 1666464484
transform 1 0 84732 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_921
timestamp 1666464484
transform 1 0 85836 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_933
timestamp 1666464484
transform 1 0 86940 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_945
timestamp 1666464484
transform 1 0 88044 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_951
timestamp 1666464484
transform 1 0 88596 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_953
timestamp 1666464484
transform 1 0 88780 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_965
timestamp 1666464484
transform 1 0 89884 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_977
timestamp 1666464484
transform 1 0 90988 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_989
timestamp 1666464484
transform 1 0 92092 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1001
timestamp 1666464484
transform 1 0 93196 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1007
timestamp 1666464484
transform 1 0 93748 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1009
timestamp 1666464484
transform 1 0 93932 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1021
timestamp 1666464484
transform 1 0 95036 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1033
timestamp 1666464484
transform 1 0 96140 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1045
timestamp 1666464484
transform 1 0 97244 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1057
timestamp 1666464484
transform 1 0 98348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1063
timestamp 1666464484
transform 1 0 98900 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1065
timestamp 1666464484
transform 1 0 99084 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1077
timestamp 1666464484
transform 1 0 100188 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1089
timestamp 1666464484
transform 1 0 101292 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1101
timestamp 1666464484
transform 1 0 102396 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1113
timestamp 1666464484
transform 1 0 103500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1119
timestamp 1666464484
transform 1 0 104052 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1121
timestamp 1666464484
transform 1 0 104236 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1133
timestamp 1666464484
transform 1 0 105340 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1145
timestamp 1666464484
transform 1 0 106444 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1157
timestamp 1666464484
transform 1 0 107548 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1169
timestamp 1666464484
transform 1 0 108652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1175
timestamp 1666464484
transform 1 0 109204 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1177
timestamp 1666464484
transform 1 0 109388 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1189
timestamp 1666464484
transform 1 0 110492 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1201
timestamp 1666464484
transform 1 0 111596 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1213
timestamp 1666464484
transform 1 0 112700 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1225
timestamp 1666464484
transform 1 0 113804 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1231
timestamp 1666464484
transform 1 0 114356 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1233
timestamp 1666464484
transform 1 0 114540 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1245
timestamp 1666464484
transform 1 0 115644 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1257
timestamp 1666464484
transform 1 0 116748 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1269
timestamp 1666464484
transform 1 0 117852 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1281
timestamp 1666464484
transform 1 0 118956 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1287
timestamp 1666464484
transform 1 0 119508 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1289
timestamp 1666464484
transform 1 0 119692 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1301
timestamp 1666464484
transform 1 0 120796 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1313
timestamp 1666464484
transform 1 0 121900 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1325
timestamp 1666464484
transform 1 0 123004 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1337
timestamp 1666464484
transform 1 0 124108 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1343
timestamp 1666464484
transform 1 0 124660 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1345
timestamp 1666464484
transform 1 0 124844 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1357
timestamp 1666464484
transform 1 0 125948 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1369
timestamp 1666464484
transform 1 0 127052 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1381
timestamp 1666464484
transform 1 0 128156 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1393
timestamp 1666464484
transform 1 0 129260 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1399
timestamp 1666464484
transform 1 0 129812 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1401
timestamp 1666464484
transform 1 0 129996 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1413
timestamp 1666464484
transform 1 0 131100 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1425
timestamp 1666464484
transform 1 0 132204 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1437
timestamp 1666464484
transform 1 0 133308 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1449
timestamp 1666464484
transform 1 0 134412 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1455
timestamp 1666464484
transform 1 0 134964 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1457
timestamp 1666464484
transform 1 0 135148 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1469
timestamp 1666464484
transform 1 0 136252 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1481
timestamp 1666464484
transform 1 0 137356 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1493
timestamp 1666464484
transform 1 0 138460 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1505
timestamp 1666464484
transform 1 0 139564 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1511
timestamp 1666464484
transform 1 0 140116 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1513
timestamp 1666464484
transform 1 0 140300 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1525
timestamp 1666464484
transform 1 0 141404 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1537
timestamp 1666464484
transform 1 0 142508 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1549
timestamp 1666464484
transform 1 0 143612 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1561
timestamp 1666464484
transform 1 0 144716 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1567
timestamp 1666464484
transform 1 0 145268 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1569
timestamp 1666464484
transform 1 0 145452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1581
timestamp 1666464484
transform 1 0 146556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1593
timestamp 1666464484
transform 1 0 147660 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1601
timestamp 1666464484
transform 1 0 148396 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1666464484
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1666464484
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1666464484
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1666464484
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1666464484
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1666464484
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1666464484
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1666464484
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1666464484
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1666464484
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1666464484
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1666464484
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1666464484
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1666464484
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1666464484
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1666464484
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1666464484
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1666464484
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1666464484
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1666464484
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1666464484
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1666464484
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1666464484
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1666464484
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1666464484
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1666464484
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1666464484
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1666464484
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1666464484
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1666464484
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1666464484
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1666464484
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1666464484
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1666464484
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1666464484
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1666464484
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1666464484
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1666464484
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1666464484
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1666464484
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1666464484
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1666464484
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1666464484
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1666464484
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1666464484
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1666464484
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1666464484
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1666464484
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1666464484
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1666464484
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1666464484
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1666464484
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1666464484
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1666464484
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1666464484
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1666464484
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1666464484
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1666464484
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1666464484
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1666464484
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_601
timestamp 1666464484
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_613
timestamp 1666464484
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_625
timestamp 1666464484
transform 1 0 58604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_637
timestamp 1666464484
transform 1 0 59708 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_643
timestamp 1666464484
transform 1 0 60260 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_645
timestamp 1666464484
transform 1 0 60444 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_657
timestamp 1666464484
transform 1 0 61548 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_669
timestamp 1666464484
transform 1 0 62652 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_681
timestamp 1666464484
transform 1 0 63756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_693
timestamp 1666464484
transform 1 0 64860 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_699
timestamp 1666464484
transform 1 0 65412 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_701
timestamp 1666464484
transform 1 0 65596 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_713
timestamp 1666464484
transform 1 0 66700 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_725
timestamp 1666464484
transform 1 0 67804 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_737
timestamp 1666464484
transform 1 0 68908 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_749
timestamp 1666464484
transform 1 0 70012 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_755
timestamp 1666464484
transform 1 0 70564 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_757
timestamp 1666464484
transform 1 0 70748 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_769
timestamp 1666464484
transform 1 0 71852 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_781
timestamp 1666464484
transform 1 0 72956 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_793
timestamp 1666464484
transform 1 0 74060 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_805
timestamp 1666464484
transform 1 0 75164 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_811
timestamp 1666464484
transform 1 0 75716 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_813
timestamp 1666464484
transform 1 0 75900 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_825
timestamp 1666464484
transform 1 0 77004 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_837
timestamp 1666464484
transform 1 0 78108 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_849
timestamp 1666464484
transform 1 0 79212 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_861
timestamp 1666464484
transform 1 0 80316 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_867
timestamp 1666464484
transform 1 0 80868 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_869
timestamp 1666464484
transform 1 0 81052 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_881
timestamp 1666464484
transform 1 0 82156 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_893
timestamp 1666464484
transform 1 0 83260 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_905
timestamp 1666464484
transform 1 0 84364 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_917
timestamp 1666464484
transform 1 0 85468 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_923
timestamp 1666464484
transform 1 0 86020 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_925
timestamp 1666464484
transform 1 0 86204 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_937
timestamp 1666464484
transform 1 0 87308 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_949
timestamp 1666464484
transform 1 0 88412 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_961
timestamp 1666464484
transform 1 0 89516 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_973
timestamp 1666464484
transform 1 0 90620 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_979
timestamp 1666464484
transform 1 0 91172 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_981
timestamp 1666464484
transform 1 0 91356 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_993
timestamp 1666464484
transform 1 0 92460 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1005
timestamp 1666464484
transform 1 0 93564 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1017
timestamp 1666464484
transform 1 0 94668 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1029
timestamp 1666464484
transform 1 0 95772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1035
timestamp 1666464484
transform 1 0 96324 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1037
timestamp 1666464484
transform 1 0 96508 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1049
timestamp 1666464484
transform 1 0 97612 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1061
timestamp 1666464484
transform 1 0 98716 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1073
timestamp 1666464484
transform 1 0 99820 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1085
timestamp 1666464484
transform 1 0 100924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1091
timestamp 1666464484
transform 1 0 101476 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1093
timestamp 1666464484
transform 1 0 101660 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1105
timestamp 1666464484
transform 1 0 102764 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1117
timestamp 1666464484
transform 1 0 103868 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1129
timestamp 1666464484
transform 1 0 104972 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1141
timestamp 1666464484
transform 1 0 106076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1147
timestamp 1666464484
transform 1 0 106628 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1149
timestamp 1666464484
transform 1 0 106812 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1161
timestamp 1666464484
transform 1 0 107916 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1173
timestamp 1666464484
transform 1 0 109020 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1185
timestamp 1666464484
transform 1 0 110124 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1197
timestamp 1666464484
transform 1 0 111228 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1203
timestamp 1666464484
transform 1 0 111780 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1205
timestamp 1666464484
transform 1 0 111964 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1217
timestamp 1666464484
transform 1 0 113068 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1229
timestamp 1666464484
transform 1 0 114172 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1241
timestamp 1666464484
transform 1 0 115276 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1253
timestamp 1666464484
transform 1 0 116380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1259
timestamp 1666464484
transform 1 0 116932 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1261
timestamp 1666464484
transform 1 0 117116 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1273
timestamp 1666464484
transform 1 0 118220 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1285
timestamp 1666464484
transform 1 0 119324 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1297
timestamp 1666464484
transform 1 0 120428 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1309
timestamp 1666464484
transform 1 0 121532 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1315
timestamp 1666464484
transform 1 0 122084 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1317
timestamp 1666464484
transform 1 0 122268 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1329
timestamp 1666464484
transform 1 0 123372 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1341
timestamp 1666464484
transform 1 0 124476 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1353
timestamp 1666464484
transform 1 0 125580 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1365
timestamp 1666464484
transform 1 0 126684 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1371
timestamp 1666464484
transform 1 0 127236 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1373
timestamp 1666464484
transform 1 0 127420 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1385
timestamp 1666464484
transform 1 0 128524 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1397
timestamp 1666464484
transform 1 0 129628 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1409
timestamp 1666464484
transform 1 0 130732 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1421
timestamp 1666464484
transform 1 0 131836 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1427
timestamp 1666464484
transform 1 0 132388 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1429
timestamp 1666464484
transform 1 0 132572 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1441
timestamp 1666464484
transform 1 0 133676 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1453
timestamp 1666464484
transform 1 0 134780 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1465
timestamp 1666464484
transform 1 0 135884 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1477
timestamp 1666464484
transform 1 0 136988 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1483
timestamp 1666464484
transform 1 0 137540 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1485
timestamp 1666464484
transform 1 0 137724 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1497
timestamp 1666464484
transform 1 0 138828 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1509
timestamp 1666464484
transform 1 0 139932 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1521
timestamp 1666464484
transform 1 0 141036 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1533
timestamp 1666464484
transform 1 0 142140 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1539
timestamp 1666464484
transform 1 0 142692 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1541
timestamp 1666464484
transform 1 0 142876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1553
timestamp 1666464484
transform 1 0 143980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1565
timestamp 1666464484
transform 1 0 145084 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1577
timestamp 1666464484
transform 1 0 146188 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1589
timestamp 1666464484
transform 1 0 147292 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1595
timestamp 1666464484
transform 1 0 147844 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1597
timestamp 1666464484
transform 1 0 148028 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1666464484
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1666464484
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1666464484
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1666464484
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1666464484
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1666464484
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1666464484
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1666464484
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1666464484
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1666464484
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1666464484
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1666464484
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1666464484
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1666464484
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1666464484
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1666464484
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1666464484
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1666464484
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1666464484
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1666464484
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1666464484
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1666464484
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1666464484
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1666464484
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1666464484
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1666464484
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1666464484
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1666464484
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1666464484
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1666464484
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1666464484
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1666464484
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1666464484
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1666464484
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1666464484
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1666464484
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1666464484
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1666464484
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1666464484
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1666464484
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1666464484
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1666464484
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1666464484
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1666464484
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1666464484
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1666464484
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1666464484
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1666464484
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1666464484
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1666464484
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1666464484
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1666464484
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1666464484
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1666464484
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1666464484
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1666464484
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1666464484
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1666464484
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1666464484
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1666464484
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_597
timestamp 1666464484
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1666464484
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1666464484
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_617
timestamp 1666464484
transform 1 0 57868 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_629
timestamp 1666464484
transform 1 0 58972 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_641
timestamp 1666464484
transform 1 0 60076 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_653
timestamp 1666464484
transform 1 0 61180 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_665
timestamp 1666464484
transform 1 0 62284 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_671
timestamp 1666464484
transform 1 0 62836 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_673
timestamp 1666464484
transform 1 0 63020 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_685
timestamp 1666464484
transform 1 0 64124 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_697
timestamp 1666464484
transform 1 0 65228 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_709
timestamp 1666464484
transform 1 0 66332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_721
timestamp 1666464484
transform 1 0 67436 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_727
timestamp 1666464484
transform 1 0 67988 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_729
timestamp 1666464484
transform 1 0 68172 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_741
timestamp 1666464484
transform 1 0 69276 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_753
timestamp 1666464484
transform 1 0 70380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_765
timestamp 1666464484
transform 1 0 71484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_777
timestamp 1666464484
transform 1 0 72588 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_783
timestamp 1666464484
transform 1 0 73140 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_785
timestamp 1666464484
transform 1 0 73324 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_797
timestamp 1666464484
transform 1 0 74428 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_809
timestamp 1666464484
transform 1 0 75532 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_821
timestamp 1666464484
transform 1 0 76636 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_833
timestamp 1666464484
transform 1 0 77740 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_839
timestamp 1666464484
transform 1 0 78292 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_841
timestamp 1666464484
transform 1 0 78476 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_853
timestamp 1666464484
transform 1 0 79580 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_865
timestamp 1666464484
transform 1 0 80684 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_877
timestamp 1666464484
transform 1 0 81788 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_889
timestamp 1666464484
transform 1 0 82892 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_895
timestamp 1666464484
transform 1 0 83444 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_897
timestamp 1666464484
transform 1 0 83628 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_909
timestamp 1666464484
transform 1 0 84732 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_921
timestamp 1666464484
transform 1 0 85836 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_933
timestamp 1666464484
transform 1 0 86940 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_945
timestamp 1666464484
transform 1 0 88044 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_951
timestamp 1666464484
transform 1 0 88596 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_953
timestamp 1666464484
transform 1 0 88780 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_965
timestamp 1666464484
transform 1 0 89884 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_977
timestamp 1666464484
transform 1 0 90988 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_989
timestamp 1666464484
transform 1 0 92092 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1001
timestamp 1666464484
transform 1 0 93196 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1007
timestamp 1666464484
transform 1 0 93748 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1009
timestamp 1666464484
transform 1 0 93932 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1021
timestamp 1666464484
transform 1 0 95036 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1033
timestamp 1666464484
transform 1 0 96140 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1045
timestamp 1666464484
transform 1 0 97244 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1057
timestamp 1666464484
transform 1 0 98348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1063
timestamp 1666464484
transform 1 0 98900 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1065
timestamp 1666464484
transform 1 0 99084 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1077
timestamp 1666464484
transform 1 0 100188 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1089
timestamp 1666464484
transform 1 0 101292 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1101
timestamp 1666464484
transform 1 0 102396 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1113
timestamp 1666464484
transform 1 0 103500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1119
timestamp 1666464484
transform 1 0 104052 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1121
timestamp 1666464484
transform 1 0 104236 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1133
timestamp 1666464484
transform 1 0 105340 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1145
timestamp 1666464484
transform 1 0 106444 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1157
timestamp 1666464484
transform 1 0 107548 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1169
timestamp 1666464484
transform 1 0 108652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1175
timestamp 1666464484
transform 1 0 109204 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1177
timestamp 1666464484
transform 1 0 109388 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1189
timestamp 1666464484
transform 1 0 110492 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1201
timestamp 1666464484
transform 1 0 111596 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1213
timestamp 1666464484
transform 1 0 112700 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1225
timestamp 1666464484
transform 1 0 113804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1231
timestamp 1666464484
transform 1 0 114356 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1233
timestamp 1666464484
transform 1 0 114540 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1245
timestamp 1666464484
transform 1 0 115644 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1257
timestamp 1666464484
transform 1 0 116748 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1269
timestamp 1666464484
transform 1 0 117852 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1281
timestamp 1666464484
transform 1 0 118956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1287
timestamp 1666464484
transform 1 0 119508 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1289
timestamp 1666464484
transform 1 0 119692 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1301
timestamp 1666464484
transform 1 0 120796 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1313
timestamp 1666464484
transform 1 0 121900 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1325
timestamp 1666464484
transform 1 0 123004 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1337
timestamp 1666464484
transform 1 0 124108 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1343
timestamp 1666464484
transform 1 0 124660 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1345
timestamp 1666464484
transform 1 0 124844 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1357
timestamp 1666464484
transform 1 0 125948 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1369
timestamp 1666464484
transform 1 0 127052 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1381
timestamp 1666464484
transform 1 0 128156 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1393
timestamp 1666464484
transform 1 0 129260 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1399
timestamp 1666464484
transform 1 0 129812 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1401
timestamp 1666464484
transform 1 0 129996 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1413
timestamp 1666464484
transform 1 0 131100 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1425
timestamp 1666464484
transform 1 0 132204 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1437
timestamp 1666464484
transform 1 0 133308 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1449
timestamp 1666464484
transform 1 0 134412 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1455
timestamp 1666464484
transform 1 0 134964 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1457
timestamp 1666464484
transform 1 0 135148 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1469
timestamp 1666464484
transform 1 0 136252 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1481
timestamp 1666464484
transform 1 0 137356 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1493
timestamp 1666464484
transform 1 0 138460 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1505
timestamp 1666464484
transform 1 0 139564 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1511
timestamp 1666464484
transform 1 0 140116 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1513
timestamp 1666464484
transform 1 0 140300 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1525
timestamp 1666464484
transform 1 0 141404 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1537
timestamp 1666464484
transform 1 0 142508 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1549
timestamp 1666464484
transform 1 0 143612 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1561
timestamp 1666464484
transform 1 0 144716 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1567
timestamp 1666464484
transform 1 0 145268 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1569
timestamp 1666464484
transform 1 0 145452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1581
timestamp 1666464484
transform 1 0 146556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1593
timestamp 1666464484
transform 1 0 147660 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1601
timestamp 1666464484
transform 1 0 148396 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1666464484
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1666464484
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1666464484
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1666464484
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1666464484
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1666464484
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1666464484
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1666464484
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1666464484
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1666464484
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1666464484
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1666464484
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1666464484
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1666464484
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1666464484
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1666464484
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1666464484
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1666464484
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1666464484
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1666464484
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1666464484
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1666464484
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1666464484
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1666464484
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1666464484
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1666464484
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1666464484
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1666464484
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1666464484
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1666464484
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1666464484
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1666464484
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1666464484
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1666464484
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1666464484
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1666464484
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1666464484
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1666464484
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1666464484
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1666464484
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1666464484
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1666464484
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1666464484
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1666464484
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1666464484
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1666464484
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1666464484
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1666464484
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1666464484
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1666464484
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1666464484
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1666464484
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1666464484
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1666464484
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1666464484
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1666464484
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1666464484
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1666464484
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1666464484
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1666464484
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_601
timestamp 1666464484
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_613
timestamp 1666464484
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_625
timestamp 1666464484
transform 1 0 58604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_637
timestamp 1666464484
transform 1 0 59708 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_643
timestamp 1666464484
transform 1 0 60260 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_645
timestamp 1666464484
transform 1 0 60444 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_657
timestamp 1666464484
transform 1 0 61548 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_669
timestamp 1666464484
transform 1 0 62652 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_681
timestamp 1666464484
transform 1 0 63756 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_693
timestamp 1666464484
transform 1 0 64860 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_699
timestamp 1666464484
transform 1 0 65412 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_701
timestamp 1666464484
transform 1 0 65596 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_713
timestamp 1666464484
transform 1 0 66700 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_725
timestamp 1666464484
transform 1 0 67804 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_737
timestamp 1666464484
transform 1 0 68908 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_749
timestamp 1666464484
transform 1 0 70012 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_755
timestamp 1666464484
transform 1 0 70564 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_757
timestamp 1666464484
transform 1 0 70748 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_769
timestamp 1666464484
transform 1 0 71852 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_781
timestamp 1666464484
transform 1 0 72956 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_793
timestamp 1666464484
transform 1 0 74060 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_805
timestamp 1666464484
transform 1 0 75164 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_811
timestamp 1666464484
transform 1 0 75716 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_813
timestamp 1666464484
transform 1 0 75900 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_825
timestamp 1666464484
transform 1 0 77004 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_837
timestamp 1666464484
transform 1 0 78108 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_849
timestamp 1666464484
transform 1 0 79212 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_861
timestamp 1666464484
transform 1 0 80316 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_867
timestamp 1666464484
transform 1 0 80868 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_869
timestamp 1666464484
transform 1 0 81052 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_881
timestamp 1666464484
transform 1 0 82156 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_893
timestamp 1666464484
transform 1 0 83260 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_905
timestamp 1666464484
transform 1 0 84364 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_917
timestamp 1666464484
transform 1 0 85468 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_923
timestamp 1666464484
transform 1 0 86020 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_925
timestamp 1666464484
transform 1 0 86204 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_937
timestamp 1666464484
transform 1 0 87308 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_949
timestamp 1666464484
transform 1 0 88412 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_961
timestamp 1666464484
transform 1 0 89516 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_973
timestamp 1666464484
transform 1 0 90620 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_979
timestamp 1666464484
transform 1 0 91172 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_981
timestamp 1666464484
transform 1 0 91356 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_993
timestamp 1666464484
transform 1 0 92460 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1005
timestamp 1666464484
transform 1 0 93564 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1017
timestamp 1666464484
transform 1 0 94668 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1029
timestamp 1666464484
transform 1 0 95772 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1035
timestamp 1666464484
transform 1 0 96324 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1037
timestamp 1666464484
transform 1 0 96508 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1049
timestamp 1666464484
transform 1 0 97612 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1061
timestamp 1666464484
transform 1 0 98716 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1073
timestamp 1666464484
transform 1 0 99820 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1085
timestamp 1666464484
transform 1 0 100924 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1091
timestamp 1666464484
transform 1 0 101476 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1093
timestamp 1666464484
transform 1 0 101660 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1105
timestamp 1666464484
transform 1 0 102764 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1117
timestamp 1666464484
transform 1 0 103868 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1129
timestamp 1666464484
transform 1 0 104972 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1141
timestamp 1666464484
transform 1 0 106076 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1147
timestamp 1666464484
transform 1 0 106628 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1149
timestamp 1666464484
transform 1 0 106812 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1161
timestamp 1666464484
transform 1 0 107916 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1173
timestamp 1666464484
transform 1 0 109020 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1185
timestamp 1666464484
transform 1 0 110124 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1197
timestamp 1666464484
transform 1 0 111228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1203
timestamp 1666464484
transform 1 0 111780 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1205
timestamp 1666464484
transform 1 0 111964 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1217
timestamp 1666464484
transform 1 0 113068 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1229
timestamp 1666464484
transform 1 0 114172 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1241
timestamp 1666464484
transform 1 0 115276 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1253
timestamp 1666464484
transform 1 0 116380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1259
timestamp 1666464484
transform 1 0 116932 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1261
timestamp 1666464484
transform 1 0 117116 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1273
timestamp 1666464484
transform 1 0 118220 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1285
timestamp 1666464484
transform 1 0 119324 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1297
timestamp 1666464484
transform 1 0 120428 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1309
timestamp 1666464484
transform 1 0 121532 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1315
timestamp 1666464484
transform 1 0 122084 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1317
timestamp 1666464484
transform 1 0 122268 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1329
timestamp 1666464484
transform 1 0 123372 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1341
timestamp 1666464484
transform 1 0 124476 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1353
timestamp 1666464484
transform 1 0 125580 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1365
timestamp 1666464484
transform 1 0 126684 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1371
timestamp 1666464484
transform 1 0 127236 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1373
timestamp 1666464484
transform 1 0 127420 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1385
timestamp 1666464484
transform 1 0 128524 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1397
timestamp 1666464484
transform 1 0 129628 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1409
timestamp 1666464484
transform 1 0 130732 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1421
timestamp 1666464484
transform 1 0 131836 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1427
timestamp 1666464484
transform 1 0 132388 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1429
timestamp 1666464484
transform 1 0 132572 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1441
timestamp 1666464484
transform 1 0 133676 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1453
timestamp 1666464484
transform 1 0 134780 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1465
timestamp 1666464484
transform 1 0 135884 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1477
timestamp 1666464484
transform 1 0 136988 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1483
timestamp 1666464484
transform 1 0 137540 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1485
timestamp 1666464484
transform 1 0 137724 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1497
timestamp 1666464484
transform 1 0 138828 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1509
timestamp 1666464484
transform 1 0 139932 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1521
timestamp 1666464484
transform 1 0 141036 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1533
timestamp 1666464484
transform 1 0 142140 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1539
timestamp 1666464484
transform 1 0 142692 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1541
timestamp 1666464484
transform 1 0 142876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1553
timestamp 1666464484
transform 1 0 143980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1565
timestamp 1666464484
transform 1 0 145084 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1577
timestamp 1666464484
transform 1 0 146188 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1589
timestamp 1666464484
transform 1 0 147292 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1595
timestamp 1666464484
transform 1 0 147844 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1597
timestamp 1666464484
transform 1 0 148028 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1666464484
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1666464484
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1666464484
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1666464484
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1666464484
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1666464484
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1666464484
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1666464484
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1666464484
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1666464484
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1666464484
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1666464484
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1666464484
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1666464484
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1666464484
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1666464484
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1666464484
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1666464484
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1666464484
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1666464484
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1666464484
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1666464484
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1666464484
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1666464484
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1666464484
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1666464484
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1666464484
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1666464484
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1666464484
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1666464484
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1666464484
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1666464484
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1666464484
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1666464484
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1666464484
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1666464484
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1666464484
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1666464484
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1666464484
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1666464484
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1666464484
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1666464484
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1666464484
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1666464484
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1666464484
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1666464484
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1666464484
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1666464484
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1666464484
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1666464484
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1666464484
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1666464484
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1666464484
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1666464484
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1666464484
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1666464484
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1666464484
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1666464484
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1666464484
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1666464484
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_597
timestamp 1666464484
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1666464484
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1666464484
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_617
timestamp 1666464484
transform 1 0 57868 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_629
timestamp 1666464484
transform 1 0 58972 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_641
timestamp 1666464484
transform 1 0 60076 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_653
timestamp 1666464484
transform 1 0 61180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_665
timestamp 1666464484
transform 1 0 62284 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_671
timestamp 1666464484
transform 1 0 62836 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_673
timestamp 1666464484
transform 1 0 63020 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_685
timestamp 1666464484
transform 1 0 64124 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_697
timestamp 1666464484
transform 1 0 65228 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_709
timestamp 1666464484
transform 1 0 66332 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_721
timestamp 1666464484
transform 1 0 67436 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_727
timestamp 1666464484
transform 1 0 67988 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_729
timestamp 1666464484
transform 1 0 68172 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_741
timestamp 1666464484
transform 1 0 69276 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_753
timestamp 1666464484
transform 1 0 70380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_765
timestamp 1666464484
transform 1 0 71484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_777
timestamp 1666464484
transform 1 0 72588 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_783
timestamp 1666464484
transform 1 0 73140 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_785
timestamp 1666464484
transform 1 0 73324 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_797
timestamp 1666464484
transform 1 0 74428 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_809
timestamp 1666464484
transform 1 0 75532 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_821
timestamp 1666464484
transform 1 0 76636 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_833
timestamp 1666464484
transform 1 0 77740 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_839
timestamp 1666464484
transform 1 0 78292 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_841
timestamp 1666464484
transform 1 0 78476 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_853
timestamp 1666464484
transform 1 0 79580 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_865
timestamp 1666464484
transform 1 0 80684 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_877
timestamp 1666464484
transform 1 0 81788 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_889
timestamp 1666464484
transform 1 0 82892 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_895
timestamp 1666464484
transform 1 0 83444 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_897
timestamp 1666464484
transform 1 0 83628 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_909
timestamp 1666464484
transform 1 0 84732 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_921
timestamp 1666464484
transform 1 0 85836 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_933
timestamp 1666464484
transform 1 0 86940 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_945
timestamp 1666464484
transform 1 0 88044 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_951
timestamp 1666464484
transform 1 0 88596 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_953
timestamp 1666464484
transform 1 0 88780 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_965
timestamp 1666464484
transform 1 0 89884 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_977
timestamp 1666464484
transform 1 0 90988 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_989
timestamp 1666464484
transform 1 0 92092 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1001
timestamp 1666464484
transform 1 0 93196 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1007
timestamp 1666464484
transform 1 0 93748 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1009
timestamp 1666464484
transform 1 0 93932 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1021
timestamp 1666464484
transform 1 0 95036 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1033
timestamp 1666464484
transform 1 0 96140 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1045
timestamp 1666464484
transform 1 0 97244 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1057
timestamp 1666464484
transform 1 0 98348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1063
timestamp 1666464484
transform 1 0 98900 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1065
timestamp 1666464484
transform 1 0 99084 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1077
timestamp 1666464484
transform 1 0 100188 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1089
timestamp 1666464484
transform 1 0 101292 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1101
timestamp 1666464484
transform 1 0 102396 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1113
timestamp 1666464484
transform 1 0 103500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1119
timestamp 1666464484
transform 1 0 104052 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1121
timestamp 1666464484
transform 1 0 104236 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1133
timestamp 1666464484
transform 1 0 105340 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1145
timestamp 1666464484
transform 1 0 106444 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1157
timestamp 1666464484
transform 1 0 107548 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1169
timestamp 1666464484
transform 1 0 108652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1175
timestamp 1666464484
transform 1 0 109204 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1177
timestamp 1666464484
transform 1 0 109388 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1189
timestamp 1666464484
transform 1 0 110492 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1201
timestamp 1666464484
transform 1 0 111596 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1213
timestamp 1666464484
transform 1 0 112700 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1225
timestamp 1666464484
transform 1 0 113804 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1231
timestamp 1666464484
transform 1 0 114356 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1233
timestamp 1666464484
transform 1 0 114540 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1245
timestamp 1666464484
transform 1 0 115644 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1257
timestamp 1666464484
transform 1 0 116748 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1269
timestamp 1666464484
transform 1 0 117852 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1281
timestamp 1666464484
transform 1 0 118956 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1287
timestamp 1666464484
transform 1 0 119508 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1289
timestamp 1666464484
transform 1 0 119692 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1301
timestamp 1666464484
transform 1 0 120796 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1313
timestamp 1666464484
transform 1 0 121900 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1325
timestamp 1666464484
transform 1 0 123004 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1337
timestamp 1666464484
transform 1 0 124108 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1343
timestamp 1666464484
transform 1 0 124660 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1345
timestamp 1666464484
transform 1 0 124844 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1357
timestamp 1666464484
transform 1 0 125948 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1369
timestamp 1666464484
transform 1 0 127052 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1381
timestamp 1666464484
transform 1 0 128156 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1393
timestamp 1666464484
transform 1 0 129260 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1399
timestamp 1666464484
transform 1 0 129812 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1401
timestamp 1666464484
transform 1 0 129996 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1413
timestamp 1666464484
transform 1 0 131100 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1425
timestamp 1666464484
transform 1 0 132204 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1437
timestamp 1666464484
transform 1 0 133308 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1449
timestamp 1666464484
transform 1 0 134412 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1455
timestamp 1666464484
transform 1 0 134964 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1457
timestamp 1666464484
transform 1 0 135148 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1469
timestamp 1666464484
transform 1 0 136252 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1481
timestamp 1666464484
transform 1 0 137356 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1493
timestamp 1666464484
transform 1 0 138460 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1505
timestamp 1666464484
transform 1 0 139564 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1511
timestamp 1666464484
transform 1 0 140116 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1513
timestamp 1666464484
transform 1 0 140300 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1525
timestamp 1666464484
transform 1 0 141404 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1537
timestamp 1666464484
transform 1 0 142508 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1549
timestamp 1666464484
transform 1 0 143612 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1561
timestamp 1666464484
transform 1 0 144716 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1567
timestamp 1666464484
transform 1 0 145268 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1569
timestamp 1666464484
transform 1 0 145452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1581
timestamp 1666464484
transform 1 0 146556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1593
timestamp 1666464484
transform 1 0 147660 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1601
timestamp 1666464484
transform 1 0 148396 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1666464484
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1666464484
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1666464484
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1666464484
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1666464484
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1666464484
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1666464484
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1666464484
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1666464484
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1666464484
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1666464484
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1666464484
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1666464484
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1666464484
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1666464484
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1666464484
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1666464484
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1666464484
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1666464484
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1666464484
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1666464484
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1666464484
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1666464484
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1666464484
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1666464484
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1666464484
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1666464484
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1666464484
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1666464484
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1666464484
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1666464484
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1666464484
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1666464484
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1666464484
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1666464484
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1666464484
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1666464484
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1666464484
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1666464484
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1666464484
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1666464484
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1666464484
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1666464484
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1666464484
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1666464484
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1666464484
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1666464484
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1666464484
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1666464484
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1666464484
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1666464484
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1666464484
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1666464484
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1666464484
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1666464484
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1666464484
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1666464484
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1666464484
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1666464484
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1666464484
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_601
timestamp 1666464484
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_613
timestamp 1666464484
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_625
timestamp 1666464484
transform 1 0 58604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_637
timestamp 1666464484
transform 1 0 59708 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_643
timestamp 1666464484
transform 1 0 60260 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_645
timestamp 1666464484
transform 1 0 60444 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_657
timestamp 1666464484
transform 1 0 61548 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_669
timestamp 1666464484
transform 1 0 62652 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_681
timestamp 1666464484
transform 1 0 63756 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_693
timestamp 1666464484
transform 1 0 64860 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_699
timestamp 1666464484
transform 1 0 65412 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_701
timestamp 1666464484
transform 1 0 65596 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_713
timestamp 1666464484
transform 1 0 66700 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_725
timestamp 1666464484
transform 1 0 67804 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_737
timestamp 1666464484
transform 1 0 68908 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_749
timestamp 1666464484
transform 1 0 70012 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_755
timestamp 1666464484
transform 1 0 70564 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_757
timestamp 1666464484
transform 1 0 70748 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_769
timestamp 1666464484
transform 1 0 71852 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_781
timestamp 1666464484
transform 1 0 72956 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_793
timestamp 1666464484
transform 1 0 74060 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_805
timestamp 1666464484
transform 1 0 75164 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_811
timestamp 1666464484
transform 1 0 75716 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_813
timestamp 1666464484
transform 1 0 75900 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_825
timestamp 1666464484
transform 1 0 77004 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_837
timestamp 1666464484
transform 1 0 78108 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_849
timestamp 1666464484
transform 1 0 79212 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_861
timestamp 1666464484
transform 1 0 80316 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_867
timestamp 1666464484
transform 1 0 80868 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_869
timestamp 1666464484
transform 1 0 81052 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_881
timestamp 1666464484
transform 1 0 82156 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_893
timestamp 1666464484
transform 1 0 83260 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_905
timestamp 1666464484
transform 1 0 84364 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_917
timestamp 1666464484
transform 1 0 85468 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_923
timestamp 1666464484
transform 1 0 86020 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_925
timestamp 1666464484
transform 1 0 86204 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_937
timestamp 1666464484
transform 1 0 87308 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_949
timestamp 1666464484
transform 1 0 88412 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_961
timestamp 1666464484
transform 1 0 89516 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_973
timestamp 1666464484
transform 1 0 90620 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_979
timestamp 1666464484
transform 1 0 91172 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_981
timestamp 1666464484
transform 1 0 91356 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_993
timestamp 1666464484
transform 1 0 92460 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1005
timestamp 1666464484
transform 1 0 93564 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1017
timestamp 1666464484
transform 1 0 94668 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1029
timestamp 1666464484
transform 1 0 95772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1035
timestamp 1666464484
transform 1 0 96324 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1037
timestamp 1666464484
transform 1 0 96508 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1049
timestamp 1666464484
transform 1 0 97612 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1061
timestamp 1666464484
transform 1 0 98716 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1073
timestamp 1666464484
transform 1 0 99820 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1085
timestamp 1666464484
transform 1 0 100924 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1091
timestamp 1666464484
transform 1 0 101476 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1093
timestamp 1666464484
transform 1 0 101660 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1105
timestamp 1666464484
transform 1 0 102764 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1117
timestamp 1666464484
transform 1 0 103868 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1129
timestamp 1666464484
transform 1 0 104972 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1141
timestamp 1666464484
transform 1 0 106076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1147
timestamp 1666464484
transform 1 0 106628 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1149
timestamp 1666464484
transform 1 0 106812 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1161
timestamp 1666464484
transform 1 0 107916 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1173
timestamp 1666464484
transform 1 0 109020 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1185
timestamp 1666464484
transform 1 0 110124 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1197
timestamp 1666464484
transform 1 0 111228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1203
timestamp 1666464484
transform 1 0 111780 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1205
timestamp 1666464484
transform 1 0 111964 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1217
timestamp 1666464484
transform 1 0 113068 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1229
timestamp 1666464484
transform 1 0 114172 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1241
timestamp 1666464484
transform 1 0 115276 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1253
timestamp 1666464484
transform 1 0 116380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1259
timestamp 1666464484
transform 1 0 116932 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1261
timestamp 1666464484
transform 1 0 117116 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1273
timestamp 1666464484
transform 1 0 118220 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1285
timestamp 1666464484
transform 1 0 119324 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1297
timestamp 1666464484
transform 1 0 120428 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1309
timestamp 1666464484
transform 1 0 121532 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1315
timestamp 1666464484
transform 1 0 122084 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1317
timestamp 1666464484
transform 1 0 122268 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1329
timestamp 1666464484
transform 1 0 123372 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1341
timestamp 1666464484
transform 1 0 124476 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1353
timestamp 1666464484
transform 1 0 125580 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1365
timestamp 1666464484
transform 1 0 126684 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1371
timestamp 1666464484
transform 1 0 127236 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1373
timestamp 1666464484
transform 1 0 127420 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1385
timestamp 1666464484
transform 1 0 128524 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1397
timestamp 1666464484
transform 1 0 129628 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1409
timestamp 1666464484
transform 1 0 130732 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1421
timestamp 1666464484
transform 1 0 131836 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1427
timestamp 1666464484
transform 1 0 132388 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1429
timestamp 1666464484
transform 1 0 132572 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1441
timestamp 1666464484
transform 1 0 133676 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1453
timestamp 1666464484
transform 1 0 134780 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1465
timestamp 1666464484
transform 1 0 135884 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1477
timestamp 1666464484
transform 1 0 136988 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1483
timestamp 1666464484
transform 1 0 137540 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1485
timestamp 1666464484
transform 1 0 137724 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1497
timestamp 1666464484
transform 1 0 138828 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1509
timestamp 1666464484
transform 1 0 139932 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1521
timestamp 1666464484
transform 1 0 141036 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1533
timestamp 1666464484
transform 1 0 142140 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1539
timestamp 1666464484
transform 1 0 142692 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1541
timestamp 1666464484
transform 1 0 142876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1553
timestamp 1666464484
transform 1 0 143980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1565
timestamp 1666464484
transform 1 0 145084 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1577
timestamp 1666464484
transform 1 0 146188 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1589
timestamp 1666464484
transform 1 0 147292 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1595
timestamp 1666464484
transform 1 0 147844 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1597
timestamp 1666464484
transform 1 0 148028 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1666464484
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1666464484
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1666464484
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1666464484
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1666464484
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1666464484
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1666464484
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1666464484
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1666464484
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1666464484
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1666464484
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1666464484
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1666464484
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1666464484
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1666464484
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1666464484
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1666464484
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1666464484
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1666464484
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1666464484
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1666464484
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1666464484
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1666464484
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1666464484
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1666464484
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1666464484
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1666464484
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1666464484
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1666464484
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1666464484
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1666464484
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1666464484
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1666464484
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1666464484
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1666464484
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1666464484
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1666464484
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1666464484
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1666464484
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1666464484
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1666464484
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1666464484
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1666464484
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1666464484
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1666464484
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1666464484
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1666464484
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1666464484
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1666464484
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1666464484
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1666464484
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1666464484
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1666464484
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1666464484
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1666464484
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1666464484
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1666464484
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1666464484
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1666464484
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1666464484
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_597
timestamp 1666464484
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1666464484
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1666464484
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_617
timestamp 1666464484
transform 1 0 57868 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_629
timestamp 1666464484
transform 1 0 58972 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_641
timestamp 1666464484
transform 1 0 60076 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_653
timestamp 1666464484
transform 1 0 61180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_665
timestamp 1666464484
transform 1 0 62284 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_671
timestamp 1666464484
transform 1 0 62836 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_673
timestamp 1666464484
transform 1 0 63020 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_685
timestamp 1666464484
transform 1 0 64124 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_697
timestamp 1666464484
transform 1 0 65228 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_709
timestamp 1666464484
transform 1 0 66332 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_721
timestamp 1666464484
transform 1 0 67436 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_727
timestamp 1666464484
transform 1 0 67988 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_729
timestamp 1666464484
transform 1 0 68172 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_741
timestamp 1666464484
transform 1 0 69276 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_753
timestamp 1666464484
transform 1 0 70380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_765
timestamp 1666464484
transform 1 0 71484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_777
timestamp 1666464484
transform 1 0 72588 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_783
timestamp 1666464484
transform 1 0 73140 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_785
timestamp 1666464484
transform 1 0 73324 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_797
timestamp 1666464484
transform 1 0 74428 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_809
timestamp 1666464484
transform 1 0 75532 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_821
timestamp 1666464484
transform 1 0 76636 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_833
timestamp 1666464484
transform 1 0 77740 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_839
timestamp 1666464484
transform 1 0 78292 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_841
timestamp 1666464484
transform 1 0 78476 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_853
timestamp 1666464484
transform 1 0 79580 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_865
timestamp 1666464484
transform 1 0 80684 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_877
timestamp 1666464484
transform 1 0 81788 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_889
timestamp 1666464484
transform 1 0 82892 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_895
timestamp 1666464484
transform 1 0 83444 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_897
timestamp 1666464484
transform 1 0 83628 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_909
timestamp 1666464484
transform 1 0 84732 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_921
timestamp 1666464484
transform 1 0 85836 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_933
timestamp 1666464484
transform 1 0 86940 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_945
timestamp 1666464484
transform 1 0 88044 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_951
timestamp 1666464484
transform 1 0 88596 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_953
timestamp 1666464484
transform 1 0 88780 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_965
timestamp 1666464484
transform 1 0 89884 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_977
timestamp 1666464484
transform 1 0 90988 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_989
timestamp 1666464484
transform 1 0 92092 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1001
timestamp 1666464484
transform 1 0 93196 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1007
timestamp 1666464484
transform 1 0 93748 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1009
timestamp 1666464484
transform 1 0 93932 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1021
timestamp 1666464484
transform 1 0 95036 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1033
timestamp 1666464484
transform 1 0 96140 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1045
timestamp 1666464484
transform 1 0 97244 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1057
timestamp 1666464484
transform 1 0 98348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1063
timestamp 1666464484
transform 1 0 98900 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1065
timestamp 1666464484
transform 1 0 99084 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1077
timestamp 1666464484
transform 1 0 100188 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1089
timestamp 1666464484
transform 1 0 101292 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1101
timestamp 1666464484
transform 1 0 102396 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1113
timestamp 1666464484
transform 1 0 103500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1119
timestamp 1666464484
transform 1 0 104052 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1121
timestamp 1666464484
transform 1 0 104236 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1133
timestamp 1666464484
transform 1 0 105340 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1145
timestamp 1666464484
transform 1 0 106444 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1157
timestamp 1666464484
transform 1 0 107548 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1169
timestamp 1666464484
transform 1 0 108652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1175
timestamp 1666464484
transform 1 0 109204 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1177
timestamp 1666464484
transform 1 0 109388 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1189
timestamp 1666464484
transform 1 0 110492 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1201
timestamp 1666464484
transform 1 0 111596 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1213
timestamp 1666464484
transform 1 0 112700 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1225
timestamp 1666464484
transform 1 0 113804 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1231
timestamp 1666464484
transform 1 0 114356 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1233
timestamp 1666464484
transform 1 0 114540 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1245
timestamp 1666464484
transform 1 0 115644 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1257
timestamp 1666464484
transform 1 0 116748 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1269
timestamp 1666464484
transform 1 0 117852 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1281
timestamp 1666464484
transform 1 0 118956 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1287
timestamp 1666464484
transform 1 0 119508 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1289
timestamp 1666464484
transform 1 0 119692 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1301
timestamp 1666464484
transform 1 0 120796 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1313
timestamp 1666464484
transform 1 0 121900 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1325
timestamp 1666464484
transform 1 0 123004 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1337
timestamp 1666464484
transform 1 0 124108 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1343
timestamp 1666464484
transform 1 0 124660 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1345
timestamp 1666464484
transform 1 0 124844 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1357
timestamp 1666464484
transform 1 0 125948 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1369
timestamp 1666464484
transform 1 0 127052 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1381
timestamp 1666464484
transform 1 0 128156 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1393
timestamp 1666464484
transform 1 0 129260 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1399
timestamp 1666464484
transform 1 0 129812 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1401
timestamp 1666464484
transform 1 0 129996 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1413
timestamp 1666464484
transform 1 0 131100 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1425
timestamp 1666464484
transform 1 0 132204 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1437
timestamp 1666464484
transform 1 0 133308 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1449
timestamp 1666464484
transform 1 0 134412 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1455
timestamp 1666464484
transform 1 0 134964 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1457
timestamp 1666464484
transform 1 0 135148 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1469
timestamp 1666464484
transform 1 0 136252 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1481
timestamp 1666464484
transform 1 0 137356 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1493
timestamp 1666464484
transform 1 0 138460 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1505
timestamp 1666464484
transform 1 0 139564 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1511
timestamp 1666464484
transform 1 0 140116 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1513
timestamp 1666464484
transform 1 0 140300 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1525
timestamp 1666464484
transform 1 0 141404 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1537
timestamp 1666464484
transform 1 0 142508 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1549
timestamp 1666464484
transform 1 0 143612 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1561
timestamp 1666464484
transform 1 0 144716 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1567
timestamp 1666464484
transform 1 0 145268 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1569
timestamp 1666464484
transform 1 0 145452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1581
timestamp 1666464484
transform 1 0 146556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1593
timestamp 1666464484
transform 1 0 147660 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1601
timestamp 1666464484
transform 1 0 148396 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1666464484
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1666464484
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1666464484
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1666464484
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1666464484
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1666464484
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1666464484
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1666464484
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1666464484
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1666464484
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1666464484
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1666464484
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1666464484
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1666464484
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1666464484
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1666464484
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1666464484
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1666464484
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1666464484
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1666464484
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1666464484
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1666464484
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1666464484
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1666464484
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1666464484
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1666464484
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1666464484
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1666464484
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1666464484
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1666464484
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1666464484
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1666464484
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1666464484
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1666464484
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1666464484
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1666464484
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1666464484
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1666464484
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1666464484
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1666464484
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1666464484
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1666464484
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1666464484
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1666464484
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1666464484
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1666464484
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1666464484
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1666464484
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1666464484
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1666464484
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1666464484
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1666464484
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1666464484
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1666464484
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1666464484
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1666464484
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1666464484
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1666464484
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1666464484
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1666464484
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_601
timestamp 1666464484
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_613
timestamp 1666464484
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_625
timestamp 1666464484
transform 1 0 58604 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_637
timestamp 1666464484
transform 1 0 59708 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_643
timestamp 1666464484
transform 1 0 60260 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_645
timestamp 1666464484
transform 1 0 60444 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_657
timestamp 1666464484
transform 1 0 61548 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_669
timestamp 1666464484
transform 1 0 62652 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_681
timestamp 1666464484
transform 1 0 63756 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_693
timestamp 1666464484
transform 1 0 64860 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_699
timestamp 1666464484
transform 1 0 65412 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_701
timestamp 1666464484
transform 1 0 65596 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_713
timestamp 1666464484
transform 1 0 66700 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_725
timestamp 1666464484
transform 1 0 67804 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_737
timestamp 1666464484
transform 1 0 68908 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_749
timestamp 1666464484
transform 1 0 70012 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_755
timestamp 1666464484
transform 1 0 70564 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_757
timestamp 1666464484
transform 1 0 70748 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_769
timestamp 1666464484
transform 1 0 71852 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_781
timestamp 1666464484
transform 1 0 72956 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_793
timestamp 1666464484
transform 1 0 74060 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_805
timestamp 1666464484
transform 1 0 75164 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_811
timestamp 1666464484
transform 1 0 75716 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_813
timestamp 1666464484
transform 1 0 75900 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_825
timestamp 1666464484
transform 1 0 77004 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_837
timestamp 1666464484
transform 1 0 78108 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_849
timestamp 1666464484
transform 1 0 79212 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_861
timestamp 1666464484
transform 1 0 80316 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_867
timestamp 1666464484
transform 1 0 80868 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_869
timestamp 1666464484
transform 1 0 81052 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_881
timestamp 1666464484
transform 1 0 82156 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_893
timestamp 1666464484
transform 1 0 83260 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_905
timestamp 1666464484
transform 1 0 84364 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_917
timestamp 1666464484
transform 1 0 85468 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_923
timestamp 1666464484
transform 1 0 86020 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_925
timestamp 1666464484
transform 1 0 86204 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_937
timestamp 1666464484
transform 1 0 87308 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_949
timestamp 1666464484
transform 1 0 88412 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_961
timestamp 1666464484
transform 1 0 89516 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_973
timestamp 1666464484
transform 1 0 90620 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_979
timestamp 1666464484
transform 1 0 91172 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_981
timestamp 1666464484
transform 1 0 91356 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_993
timestamp 1666464484
transform 1 0 92460 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1005
timestamp 1666464484
transform 1 0 93564 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1017
timestamp 1666464484
transform 1 0 94668 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1029
timestamp 1666464484
transform 1 0 95772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1035
timestamp 1666464484
transform 1 0 96324 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1037
timestamp 1666464484
transform 1 0 96508 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1049
timestamp 1666464484
transform 1 0 97612 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1061
timestamp 1666464484
transform 1 0 98716 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1073
timestamp 1666464484
transform 1 0 99820 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1085
timestamp 1666464484
transform 1 0 100924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1091
timestamp 1666464484
transform 1 0 101476 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1093
timestamp 1666464484
transform 1 0 101660 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1105
timestamp 1666464484
transform 1 0 102764 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1117
timestamp 1666464484
transform 1 0 103868 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1129
timestamp 1666464484
transform 1 0 104972 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1141
timestamp 1666464484
transform 1 0 106076 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1147
timestamp 1666464484
transform 1 0 106628 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1149
timestamp 1666464484
transform 1 0 106812 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1161
timestamp 1666464484
transform 1 0 107916 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1173
timestamp 1666464484
transform 1 0 109020 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1185
timestamp 1666464484
transform 1 0 110124 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1197
timestamp 1666464484
transform 1 0 111228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1203
timestamp 1666464484
transform 1 0 111780 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1205
timestamp 1666464484
transform 1 0 111964 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1217
timestamp 1666464484
transform 1 0 113068 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1229
timestamp 1666464484
transform 1 0 114172 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1241
timestamp 1666464484
transform 1 0 115276 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1253
timestamp 1666464484
transform 1 0 116380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1259
timestamp 1666464484
transform 1 0 116932 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1261
timestamp 1666464484
transform 1 0 117116 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1273
timestamp 1666464484
transform 1 0 118220 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1285
timestamp 1666464484
transform 1 0 119324 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1297
timestamp 1666464484
transform 1 0 120428 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1309
timestamp 1666464484
transform 1 0 121532 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1315
timestamp 1666464484
transform 1 0 122084 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1317
timestamp 1666464484
transform 1 0 122268 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1329
timestamp 1666464484
transform 1 0 123372 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1341
timestamp 1666464484
transform 1 0 124476 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1353
timestamp 1666464484
transform 1 0 125580 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1365
timestamp 1666464484
transform 1 0 126684 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1371
timestamp 1666464484
transform 1 0 127236 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1373
timestamp 1666464484
transform 1 0 127420 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1385
timestamp 1666464484
transform 1 0 128524 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1397
timestamp 1666464484
transform 1 0 129628 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1409
timestamp 1666464484
transform 1 0 130732 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1421
timestamp 1666464484
transform 1 0 131836 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1427
timestamp 1666464484
transform 1 0 132388 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1429
timestamp 1666464484
transform 1 0 132572 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1441
timestamp 1666464484
transform 1 0 133676 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1453
timestamp 1666464484
transform 1 0 134780 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1465
timestamp 1666464484
transform 1 0 135884 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1477
timestamp 1666464484
transform 1 0 136988 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1483
timestamp 1666464484
transform 1 0 137540 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1485
timestamp 1666464484
transform 1 0 137724 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1497
timestamp 1666464484
transform 1 0 138828 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1509
timestamp 1666464484
transform 1 0 139932 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1521
timestamp 1666464484
transform 1 0 141036 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1533
timestamp 1666464484
transform 1 0 142140 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1539
timestamp 1666464484
transform 1 0 142692 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1541
timestamp 1666464484
transform 1 0 142876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1553
timestamp 1666464484
transform 1 0 143980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1565
timestamp 1666464484
transform 1 0 145084 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1577
timestamp 1666464484
transform 1 0 146188 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1589
timestamp 1666464484
transform 1 0 147292 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1595
timestamp 1666464484
transform 1 0 147844 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1597
timestamp 1666464484
transform 1 0 148028 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1666464484
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1666464484
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1666464484
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1666464484
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1666464484
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1666464484
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1666464484
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1666464484
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1666464484
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1666464484
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1666464484
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1666464484
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1666464484
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1666464484
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1666464484
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1666464484
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1666464484
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1666464484
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1666464484
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1666464484
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1666464484
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1666464484
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1666464484
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1666464484
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1666464484
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1666464484
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1666464484
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1666464484
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1666464484
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1666464484
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1666464484
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1666464484
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1666464484
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1666464484
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1666464484
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1666464484
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1666464484
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1666464484
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1666464484
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1666464484
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1666464484
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1666464484
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1666464484
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1666464484
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1666464484
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1666464484
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1666464484
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1666464484
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1666464484
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1666464484
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1666464484
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1666464484
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1666464484
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1666464484
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1666464484
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1666464484
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1666464484
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1666464484
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1666464484
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1666464484
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_597
timestamp 1666464484
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1666464484
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1666464484
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_617
timestamp 1666464484
transform 1 0 57868 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_629
timestamp 1666464484
transform 1 0 58972 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_641
timestamp 1666464484
transform 1 0 60076 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_653
timestamp 1666464484
transform 1 0 61180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_665
timestamp 1666464484
transform 1 0 62284 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_671
timestamp 1666464484
transform 1 0 62836 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_673
timestamp 1666464484
transform 1 0 63020 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_685
timestamp 1666464484
transform 1 0 64124 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_697
timestamp 1666464484
transform 1 0 65228 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_709
timestamp 1666464484
transform 1 0 66332 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_721
timestamp 1666464484
transform 1 0 67436 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_727
timestamp 1666464484
transform 1 0 67988 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_729
timestamp 1666464484
transform 1 0 68172 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_741
timestamp 1666464484
transform 1 0 69276 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_753
timestamp 1666464484
transform 1 0 70380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_765
timestamp 1666464484
transform 1 0 71484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_777
timestamp 1666464484
transform 1 0 72588 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_783
timestamp 1666464484
transform 1 0 73140 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_785
timestamp 1666464484
transform 1 0 73324 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_797
timestamp 1666464484
transform 1 0 74428 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_809
timestamp 1666464484
transform 1 0 75532 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_821
timestamp 1666464484
transform 1 0 76636 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_833
timestamp 1666464484
transform 1 0 77740 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_839
timestamp 1666464484
transform 1 0 78292 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_841
timestamp 1666464484
transform 1 0 78476 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_853
timestamp 1666464484
transform 1 0 79580 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_865
timestamp 1666464484
transform 1 0 80684 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_877
timestamp 1666464484
transform 1 0 81788 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_889
timestamp 1666464484
transform 1 0 82892 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_895
timestamp 1666464484
transform 1 0 83444 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_897
timestamp 1666464484
transform 1 0 83628 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_909
timestamp 1666464484
transform 1 0 84732 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_921
timestamp 1666464484
transform 1 0 85836 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_933
timestamp 1666464484
transform 1 0 86940 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_945
timestamp 1666464484
transform 1 0 88044 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_951
timestamp 1666464484
transform 1 0 88596 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_953
timestamp 1666464484
transform 1 0 88780 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_965
timestamp 1666464484
transform 1 0 89884 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_977
timestamp 1666464484
transform 1 0 90988 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_989
timestamp 1666464484
transform 1 0 92092 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1001
timestamp 1666464484
transform 1 0 93196 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1007
timestamp 1666464484
transform 1 0 93748 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1009
timestamp 1666464484
transform 1 0 93932 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1021
timestamp 1666464484
transform 1 0 95036 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1033
timestamp 1666464484
transform 1 0 96140 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1045
timestamp 1666464484
transform 1 0 97244 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1057
timestamp 1666464484
transform 1 0 98348 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1063
timestamp 1666464484
transform 1 0 98900 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1065
timestamp 1666464484
transform 1 0 99084 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1077
timestamp 1666464484
transform 1 0 100188 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1089
timestamp 1666464484
transform 1 0 101292 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1101
timestamp 1666464484
transform 1 0 102396 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1113
timestamp 1666464484
transform 1 0 103500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1119
timestamp 1666464484
transform 1 0 104052 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1121
timestamp 1666464484
transform 1 0 104236 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1133
timestamp 1666464484
transform 1 0 105340 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1145
timestamp 1666464484
transform 1 0 106444 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1157
timestamp 1666464484
transform 1 0 107548 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1169
timestamp 1666464484
transform 1 0 108652 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1175
timestamp 1666464484
transform 1 0 109204 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1177
timestamp 1666464484
transform 1 0 109388 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1189
timestamp 1666464484
transform 1 0 110492 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1201
timestamp 1666464484
transform 1 0 111596 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1213
timestamp 1666464484
transform 1 0 112700 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1225
timestamp 1666464484
transform 1 0 113804 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1231
timestamp 1666464484
transform 1 0 114356 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1233
timestamp 1666464484
transform 1 0 114540 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1245
timestamp 1666464484
transform 1 0 115644 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1257
timestamp 1666464484
transform 1 0 116748 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1269
timestamp 1666464484
transform 1 0 117852 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1281
timestamp 1666464484
transform 1 0 118956 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1287
timestamp 1666464484
transform 1 0 119508 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1289
timestamp 1666464484
transform 1 0 119692 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1301
timestamp 1666464484
transform 1 0 120796 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1313
timestamp 1666464484
transform 1 0 121900 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1325
timestamp 1666464484
transform 1 0 123004 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1337
timestamp 1666464484
transform 1 0 124108 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1343
timestamp 1666464484
transform 1 0 124660 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1345
timestamp 1666464484
transform 1 0 124844 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1357
timestamp 1666464484
transform 1 0 125948 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1369
timestamp 1666464484
transform 1 0 127052 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1381
timestamp 1666464484
transform 1 0 128156 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1393
timestamp 1666464484
transform 1 0 129260 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1399
timestamp 1666464484
transform 1 0 129812 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1401
timestamp 1666464484
transform 1 0 129996 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1413
timestamp 1666464484
transform 1 0 131100 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1425
timestamp 1666464484
transform 1 0 132204 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1437
timestamp 1666464484
transform 1 0 133308 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1449
timestamp 1666464484
transform 1 0 134412 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1455
timestamp 1666464484
transform 1 0 134964 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1457
timestamp 1666464484
transform 1 0 135148 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1469
timestamp 1666464484
transform 1 0 136252 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1481
timestamp 1666464484
transform 1 0 137356 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1493
timestamp 1666464484
transform 1 0 138460 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1505
timestamp 1666464484
transform 1 0 139564 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1511
timestamp 1666464484
transform 1 0 140116 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1513
timestamp 1666464484
transform 1 0 140300 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1525
timestamp 1666464484
transform 1 0 141404 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1537
timestamp 1666464484
transform 1 0 142508 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1549
timestamp 1666464484
transform 1 0 143612 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1561
timestamp 1666464484
transform 1 0 144716 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1567
timestamp 1666464484
transform 1 0 145268 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1569
timestamp 1666464484
transform 1 0 145452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1581
timestamp 1666464484
transform 1 0 146556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1593
timestamp 1666464484
transform 1 0 147660 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1601
timestamp 1666464484
transform 1 0 148396 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1666464484
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1666464484
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1666464484
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1666464484
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1666464484
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1666464484
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1666464484
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1666464484
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1666464484
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1666464484
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1666464484
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1666464484
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1666464484
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1666464484
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1666464484
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1666464484
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1666464484
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1666464484
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1666464484
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1666464484
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1666464484
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1666464484
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1666464484
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1666464484
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1666464484
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1666464484
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1666464484
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1666464484
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1666464484
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1666464484
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1666464484
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1666464484
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1666464484
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1666464484
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1666464484
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1666464484
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1666464484
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1666464484
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1666464484
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1666464484
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1666464484
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1666464484
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1666464484
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1666464484
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1666464484
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1666464484
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1666464484
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1666464484
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1666464484
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1666464484
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1666464484
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1666464484
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1666464484
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1666464484
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1666464484
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1666464484
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1666464484
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1666464484
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1666464484
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1666464484
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_601
timestamp 1666464484
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_613
timestamp 1666464484
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_625
timestamp 1666464484
transform 1 0 58604 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_637
timestamp 1666464484
transform 1 0 59708 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_643
timestamp 1666464484
transform 1 0 60260 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_645
timestamp 1666464484
transform 1 0 60444 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_657
timestamp 1666464484
transform 1 0 61548 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_669
timestamp 1666464484
transform 1 0 62652 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_681
timestamp 1666464484
transform 1 0 63756 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_693
timestamp 1666464484
transform 1 0 64860 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_699
timestamp 1666464484
transform 1 0 65412 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_701
timestamp 1666464484
transform 1 0 65596 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_713
timestamp 1666464484
transform 1 0 66700 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_725
timestamp 1666464484
transform 1 0 67804 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_737
timestamp 1666464484
transform 1 0 68908 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_749
timestamp 1666464484
transform 1 0 70012 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_755
timestamp 1666464484
transform 1 0 70564 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_757
timestamp 1666464484
transform 1 0 70748 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_769
timestamp 1666464484
transform 1 0 71852 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_781
timestamp 1666464484
transform 1 0 72956 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_793
timestamp 1666464484
transform 1 0 74060 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_805
timestamp 1666464484
transform 1 0 75164 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_811
timestamp 1666464484
transform 1 0 75716 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_813
timestamp 1666464484
transform 1 0 75900 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_825
timestamp 1666464484
transform 1 0 77004 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_837
timestamp 1666464484
transform 1 0 78108 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_849
timestamp 1666464484
transform 1 0 79212 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_861
timestamp 1666464484
transform 1 0 80316 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_867
timestamp 1666464484
transform 1 0 80868 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_869
timestamp 1666464484
transform 1 0 81052 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_881
timestamp 1666464484
transform 1 0 82156 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_893
timestamp 1666464484
transform 1 0 83260 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_905
timestamp 1666464484
transform 1 0 84364 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_917
timestamp 1666464484
transform 1 0 85468 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_923
timestamp 1666464484
transform 1 0 86020 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_925
timestamp 1666464484
transform 1 0 86204 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_937
timestamp 1666464484
transform 1 0 87308 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_949
timestamp 1666464484
transform 1 0 88412 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_961
timestamp 1666464484
transform 1 0 89516 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_973
timestamp 1666464484
transform 1 0 90620 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_979
timestamp 1666464484
transform 1 0 91172 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_981
timestamp 1666464484
transform 1 0 91356 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_993
timestamp 1666464484
transform 1 0 92460 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1005
timestamp 1666464484
transform 1 0 93564 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1017
timestamp 1666464484
transform 1 0 94668 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1029
timestamp 1666464484
transform 1 0 95772 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1035
timestamp 1666464484
transform 1 0 96324 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1037
timestamp 1666464484
transform 1 0 96508 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1049
timestamp 1666464484
transform 1 0 97612 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1061
timestamp 1666464484
transform 1 0 98716 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1073
timestamp 1666464484
transform 1 0 99820 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1085
timestamp 1666464484
transform 1 0 100924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1091
timestamp 1666464484
transform 1 0 101476 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1093
timestamp 1666464484
transform 1 0 101660 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1105
timestamp 1666464484
transform 1 0 102764 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1117
timestamp 1666464484
transform 1 0 103868 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1129
timestamp 1666464484
transform 1 0 104972 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1141
timestamp 1666464484
transform 1 0 106076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1147
timestamp 1666464484
transform 1 0 106628 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1149
timestamp 1666464484
transform 1 0 106812 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1161
timestamp 1666464484
transform 1 0 107916 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1173
timestamp 1666464484
transform 1 0 109020 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1185
timestamp 1666464484
transform 1 0 110124 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1197
timestamp 1666464484
transform 1 0 111228 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1203
timestamp 1666464484
transform 1 0 111780 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1205
timestamp 1666464484
transform 1 0 111964 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1217
timestamp 1666464484
transform 1 0 113068 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1229
timestamp 1666464484
transform 1 0 114172 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1241
timestamp 1666464484
transform 1 0 115276 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1253
timestamp 1666464484
transform 1 0 116380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1259
timestamp 1666464484
transform 1 0 116932 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1261
timestamp 1666464484
transform 1 0 117116 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1273
timestamp 1666464484
transform 1 0 118220 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1285
timestamp 1666464484
transform 1 0 119324 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1297
timestamp 1666464484
transform 1 0 120428 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1309
timestamp 1666464484
transform 1 0 121532 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1315
timestamp 1666464484
transform 1 0 122084 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1317
timestamp 1666464484
transform 1 0 122268 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1329
timestamp 1666464484
transform 1 0 123372 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1341
timestamp 1666464484
transform 1 0 124476 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1353
timestamp 1666464484
transform 1 0 125580 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1365
timestamp 1666464484
transform 1 0 126684 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1371
timestamp 1666464484
transform 1 0 127236 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1373
timestamp 1666464484
transform 1 0 127420 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1385
timestamp 1666464484
transform 1 0 128524 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1397
timestamp 1666464484
transform 1 0 129628 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1409
timestamp 1666464484
transform 1 0 130732 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1421
timestamp 1666464484
transform 1 0 131836 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1427
timestamp 1666464484
transform 1 0 132388 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1429
timestamp 1666464484
transform 1 0 132572 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1441
timestamp 1666464484
transform 1 0 133676 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1453
timestamp 1666464484
transform 1 0 134780 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1465
timestamp 1666464484
transform 1 0 135884 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1477
timestamp 1666464484
transform 1 0 136988 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1483
timestamp 1666464484
transform 1 0 137540 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1485
timestamp 1666464484
transform 1 0 137724 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1497
timestamp 1666464484
transform 1 0 138828 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1509
timestamp 1666464484
transform 1 0 139932 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1521
timestamp 1666464484
transform 1 0 141036 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1533
timestamp 1666464484
transform 1 0 142140 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1539
timestamp 1666464484
transform 1 0 142692 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1541
timestamp 1666464484
transform 1 0 142876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1553
timestamp 1666464484
transform 1 0 143980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1565
timestamp 1666464484
transform 1 0 145084 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1577
timestamp 1666464484
transform 1 0 146188 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1589
timestamp 1666464484
transform 1 0 147292 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1595
timestamp 1666464484
transform 1 0 147844 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1597
timestamp 1666464484
transform 1 0 148028 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1666464484
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1666464484
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1666464484
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1666464484
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1666464484
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1666464484
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1666464484
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1666464484
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1666464484
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1666464484
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1666464484
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1666464484
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1666464484
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1666464484
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1666464484
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1666464484
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1666464484
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1666464484
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1666464484
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1666464484
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1666464484
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1666464484
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1666464484
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1666464484
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1666464484
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1666464484
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1666464484
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1666464484
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1666464484
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1666464484
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1666464484
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1666464484
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1666464484
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1666464484
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1666464484
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1666464484
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1666464484
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1666464484
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1666464484
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1666464484
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1666464484
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1666464484
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1666464484
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1666464484
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1666464484
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1666464484
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1666464484
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1666464484
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1666464484
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1666464484
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1666464484
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1666464484
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1666464484
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1666464484
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1666464484
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1666464484
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1666464484
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1666464484
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1666464484
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1666464484
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_597
timestamp 1666464484
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1666464484
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1666464484
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_617
timestamp 1666464484
transform 1 0 57868 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_629
timestamp 1666464484
transform 1 0 58972 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_641
timestamp 1666464484
transform 1 0 60076 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_653
timestamp 1666464484
transform 1 0 61180 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_665
timestamp 1666464484
transform 1 0 62284 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_671
timestamp 1666464484
transform 1 0 62836 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_673
timestamp 1666464484
transform 1 0 63020 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_685
timestamp 1666464484
transform 1 0 64124 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_697
timestamp 1666464484
transform 1 0 65228 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_709
timestamp 1666464484
transform 1 0 66332 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_721
timestamp 1666464484
transform 1 0 67436 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_727
timestamp 1666464484
transform 1 0 67988 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_729
timestamp 1666464484
transform 1 0 68172 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_741
timestamp 1666464484
transform 1 0 69276 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_753
timestamp 1666464484
transform 1 0 70380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_765
timestamp 1666464484
transform 1 0 71484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_777
timestamp 1666464484
transform 1 0 72588 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_783
timestamp 1666464484
transform 1 0 73140 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_785
timestamp 1666464484
transform 1 0 73324 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_797
timestamp 1666464484
transform 1 0 74428 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_809
timestamp 1666464484
transform 1 0 75532 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_821
timestamp 1666464484
transform 1 0 76636 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_833
timestamp 1666464484
transform 1 0 77740 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_839
timestamp 1666464484
transform 1 0 78292 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_841
timestamp 1666464484
transform 1 0 78476 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_853
timestamp 1666464484
transform 1 0 79580 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_865
timestamp 1666464484
transform 1 0 80684 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_877
timestamp 1666464484
transform 1 0 81788 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_889
timestamp 1666464484
transform 1 0 82892 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_895
timestamp 1666464484
transform 1 0 83444 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_897
timestamp 1666464484
transform 1 0 83628 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_909
timestamp 1666464484
transform 1 0 84732 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_921
timestamp 1666464484
transform 1 0 85836 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_933
timestamp 1666464484
transform 1 0 86940 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_945
timestamp 1666464484
transform 1 0 88044 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_951
timestamp 1666464484
transform 1 0 88596 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_953
timestamp 1666464484
transform 1 0 88780 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_965
timestamp 1666464484
transform 1 0 89884 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_977
timestamp 1666464484
transform 1 0 90988 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_989
timestamp 1666464484
transform 1 0 92092 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1001
timestamp 1666464484
transform 1 0 93196 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1007
timestamp 1666464484
transform 1 0 93748 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1009
timestamp 1666464484
transform 1 0 93932 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1021
timestamp 1666464484
transform 1 0 95036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1033
timestamp 1666464484
transform 1 0 96140 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1045
timestamp 1666464484
transform 1 0 97244 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1057
timestamp 1666464484
transform 1 0 98348 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1063
timestamp 1666464484
transform 1 0 98900 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1065
timestamp 1666464484
transform 1 0 99084 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1077
timestamp 1666464484
transform 1 0 100188 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1089
timestamp 1666464484
transform 1 0 101292 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1101
timestamp 1666464484
transform 1 0 102396 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1113
timestamp 1666464484
transform 1 0 103500 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1119
timestamp 1666464484
transform 1 0 104052 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1121
timestamp 1666464484
transform 1 0 104236 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1133
timestamp 1666464484
transform 1 0 105340 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1145
timestamp 1666464484
transform 1 0 106444 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1157
timestamp 1666464484
transform 1 0 107548 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1169
timestamp 1666464484
transform 1 0 108652 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1175
timestamp 1666464484
transform 1 0 109204 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1177
timestamp 1666464484
transform 1 0 109388 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1189
timestamp 1666464484
transform 1 0 110492 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1201
timestamp 1666464484
transform 1 0 111596 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1213
timestamp 1666464484
transform 1 0 112700 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1225
timestamp 1666464484
transform 1 0 113804 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1231
timestamp 1666464484
transform 1 0 114356 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1233
timestamp 1666464484
transform 1 0 114540 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1245
timestamp 1666464484
transform 1 0 115644 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1257
timestamp 1666464484
transform 1 0 116748 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1269
timestamp 1666464484
transform 1 0 117852 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1281
timestamp 1666464484
transform 1 0 118956 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1287
timestamp 1666464484
transform 1 0 119508 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1289
timestamp 1666464484
transform 1 0 119692 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1301
timestamp 1666464484
transform 1 0 120796 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1313
timestamp 1666464484
transform 1 0 121900 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1325
timestamp 1666464484
transform 1 0 123004 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1337
timestamp 1666464484
transform 1 0 124108 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1343
timestamp 1666464484
transform 1 0 124660 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1345
timestamp 1666464484
transform 1 0 124844 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1357
timestamp 1666464484
transform 1 0 125948 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1369
timestamp 1666464484
transform 1 0 127052 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1381
timestamp 1666464484
transform 1 0 128156 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1393
timestamp 1666464484
transform 1 0 129260 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1399
timestamp 1666464484
transform 1 0 129812 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1401
timestamp 1666464484
transform 1 0 129996 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1413
timestamp 1666464484
transform 1 0 131100 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1425
timestamp 1666464484
transform 1 0 132204 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1437
timestamp 1666464484
transform 1 0 133308 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1449
timestamp 1666464484
transform 1 0 134412 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1455
timestamp 1666464484
transform 1 0 134964 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1457
timestamp 1666464484
transform 1 0 135148 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1469
timestamp 1666464484
transform 1 0 136252 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1481
timestamp 1666464484
transform 1 0 137356 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1493
timestamp 1666464484
transform 1 0 138460 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1505
timestamp 1666464484
transform 1 0 139564 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1511
timestamp 1666464484
transform 1 0 140116 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1513
timestamp 1666464484
transform 1 0 140300 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1525
timestamp 1666464484
transform 1 0 141404 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1537
timestamp 1666464484
transform 1 0 142508 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1549
timestamp 1666464484
transform 1 0 143612 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1561
timestamp 1666464484
transform 1 0 144716 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1567
timestamp 1666464484
transform 1 0 145268 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1569
timestamp 1666464484
transform 1 0 145452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1581
timestamp 1666464484
transform 1 0 146556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_1593
timestamp 1666464484
transform 1 0 147660 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_1601
timestamp 1666464484
transform 1 0 148396 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1666464484
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1666464484
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1666464484
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1666464484
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1666464484
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1666464484
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1666464484
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1666464484
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1666464484
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1666464484
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1666464484
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1666464484
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1666464484
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1666464484
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1666464484
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1666464484
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1666464484
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1666464484
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1666464484
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1666464484
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1666464484
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1666464484
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1666464484
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1666464484
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1666464484
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1666464484
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1666464484
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1666464484
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1666464484
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1666464484
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1666464484
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1666464484
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1666464484
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1666464484
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1666464484
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1666464484
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1666464484
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1666464484
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1666464484
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1666464484
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1666464484
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1666464484
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1666464484
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1666464484
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1666464484
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1666464484
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1666464484
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1666464484
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1666464484
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1666464484
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1666464484
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1666464484
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1666464484
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1666464484
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1666464484
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1666464484
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1666464484
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1666464484
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1666464484
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1666464484
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1666464484
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_613
timestamp 1666464484
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_625
timestamp 1666464484
transform 1 0 58604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_637
timestamp 1666464484
transform 1 0 59708 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_643
timestamp 1666464484
transform 1 0 60260 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_645
timestamp 1666464484
transform 1 0 60444 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_657
timestamp 1666464484
transform 1 0 61548 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_669
timestamp 1666464484
transform 1 0 62652 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_681
timestamp 1666464484
transform 1 0 63756 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_693
timestamp 1666464484
transform 1 0 64860 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_699
timestamp 1666464484
transform 1 0 65412 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_701
timestamp 1666464484
transform 1 0 65596 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_713
timestamp 1666464484
transform 1 0 66700 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_725
timestamp 1666464484
transform 1 0 67804 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_737
timestamp 1666464484
transform 1 0 68908 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_749
timestamp 1666464484
transform 1 0 70012 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_755
timestamp 1666464484
transform 1 0 70564 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_757
timestamp 1666464484
transform 1 0 70748 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_769
timestamp 1666464484
transform 1 0 71852 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_781
timestamp 1666464484
transform 1 0 72956 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_793
timestamp 1666464484
transform 1 0 74060 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_805
timestamp 1666464484
transform 1 0 75164 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_811
timestamp 1666464484
transform 1 0 75716 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_813
timestamp 1666464484
transform 1 0 75900 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_825
timestamp 1666464484
transform 1 0 77004 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_837
timestamp 1666464484
transform 1 0 78108 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_849
timestamp 1666464484
transform 1 0 79212 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_861
timestamp 1666464484
transform 1 0 80316 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_867
timestamp 1666464484
transform 1 0 80868 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_869
timestamp 1666464484
transform 1 0 81052 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_881
timestamp 1666464484
transform 1 0 82156 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_893
timestamp 1666464484
transform 1 0 83260 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_905
timestamp 1666464484
transform 1 0 84364 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_917
timestamp 1666464484
transform 1 0 85468 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_923
timestamp 1666464484
transform 1 0 86020 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_925
timestamp 1666464484
transform 1 0 86204 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_937
timestamp 1666464484
transform 1 0 87308 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_949
timestamp 1666464484
transform 1 0 88412 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_961
timestamp 1666464484
transform 1 0 89516 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_973
timestamp 1666464484
transform 1 0 90620 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_979
timestamp 1666464484
transform 1 0 91172 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_981
timestamp 1666464484
transform 1 0 91356 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_993
timestamp 1666464484
transform 1 0 92460 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1005
timestamp 1666464484
transform 1 0 93564 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1017
timestamp 1666464484
transform 1 0 94668 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1029
timestamp 1666464484
transform 1 0 95772 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1035
timestamp 1666464484
transform 1 0 96324 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1037
timestamp 1666464484
transform 1 0 96508 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1049
timestamp 1666464484
transform 1 0 97612 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1061
timestamp 1666464484
transform 1 0 98716 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1073
timestamp 1666464484
transform 1 0 99820 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1085
timestamp 1666464484
transform 1 0 100924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1091
timestamp 1666464484
transform 1 0 101476 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1093
timestamp 1666464484
transform 1 0 101660 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1105
timestamp 1666464484
transform 1 0 102764 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1117
timestamp 1666464484
transform 1 0 103868 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1129
timestamp 1666464484
transform 1 0 104972 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1141
timestamp 1666464484
transform 1 0 106076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1147
timestamp 1666464484
transform 1 0 106628 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1149
timestamp 1666464484
transform 1 0 106812 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1161
timestamp 1666464484
transform 1 0 107916 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1173
timestamp 1666464484
transform 1 0 109020 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1185
timestamp 1666464484
transform 1 0 110124 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1197
timestamp 1666464484
transform 1 0 111228 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1203
timestamp 1666464484
transform 1 0 111780 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1205
timestamp 1666464484
transform 1 0 111964 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1217
timestamp 1666464484
transform 1 0 113068 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1229
timestamp 1666464484
transform 1 0 114172 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1241
timestamp 1666464484
transform 1 0 115276 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1253
timestamp 1666464484
transform 1 0 116380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1259
timestamp 1666464484
transform 1 0 116932 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1261
timestamp 1666464484
transform 1 0 117116 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1273
timestamp 1666464484
transform 1 0 118220 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1285
timestamp 1666464484
transform 1 0 119324 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1297
timestamp 1666464484
transform 1 0 120428 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1309
timestamp 1666464484
transform 1 0 121532 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1315
timestamp 1666464484
transform 1 0 122084 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1317
timestamp 1666464484
transform 1 0 122268 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1329
timestamp 1666464484
transform 1 0 123372 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1341
timestamp 1666464484
transform 1 0 124476 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1353
timestamp 1666464484
transform 1 0 125580 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1365
timestamp 1666464484
transform 1 0 126684 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1371
timestamp 1666464484
transform 1 0 127236 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1373
timestamp 1666464484
transform 1 0 127420 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1385
timestamp 1666464484
transform 1 0 128524 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1397
timestamp 1666464484
transform 1 0 129628 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1409
timestamp 1666464484
transform 1 0 130732 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1421
timestamp 1666464484
transform 1 0 131836 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1427
timestamp 1666464484
transform 1 0 132388 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1429
timestamp 1666464484
transform 1 0 132572 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1441
timestamp 1666464484
transform 1 0 133676 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1453
timestamp 1666464484
transform 1 0 134780 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1465
timestamp 1666464484
transform 1 0 135884 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1477
timestamp 1666464484
transform 1 0 136988 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1483
timestamp 1666464484
transform 1 0 137540 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1485
timestamp 1666464484
transform 1 0 137724 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1497
timestamp 1666464484
transform 1 0 138828 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1509
timestamp 1666464484
transform 1 0 139932 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1521
timestamp 1666464484
transform 1 0 141036 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1533
timestamp 1666464484
transform 1 0 142140 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1539
timestamp 1666464484
transform 1 0 142692 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1541
timestamp 1666464484
transform 1 0 142876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1553
timestamp 1666464484
transform 1 0 143980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1565
timestamp 1666464484
transform 1 0 145084 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1577
timestamp 1666464484
transform 1 0 146188 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1589
timestamp 1666464484
transform 1 0 147292 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1595
timestamp 1666464484
transform 1 0 147844 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1597
timestamp 1666464484
transform 1 0 148028 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1666464484
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1666464484
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1666464484
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1666464484
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1666464484
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1666464484
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1666464484
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1666464484
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1666464484
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1666464484
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1666464484
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1666464484
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1666464484
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1666464484
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1666464484
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1666464484
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1666464484
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1666464484
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1666464484
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1666464484
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1666464484
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1666464484
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1666464484
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1666464484
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1666464484
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1666464484
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1666464484
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1666464484
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1666464484
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1666464484
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1666464484
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1666464484
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1666464484
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1666464484
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1666464484
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1666464484
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1666464484
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1666464484
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1666464484
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1666464484
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1666464484
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1666464484
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1666464484
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1666464484
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1666464484
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1666464484
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1666464484
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1666464484
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1666464484
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1666464484
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1666464484
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1666464484
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1666464484
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1666464484
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1666464484
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1666464484
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1666464484
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1666464484
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1666464484
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1666464484
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1666464484
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1666464484
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1666464484
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_617
timestamp 1666464484
transform 1 0 57868 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_629
timestamp 1666464484
transform 1 0 58972 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_641
timestamp 1666464484
transform 1 0 60076 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_653
timestamp 1666464484
transform 1 0 61180 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_665
timestamp 1666464484
transform 1 0 62284 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_671
timestamp 1666464484
transform 1 0 62836 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_673
timestamp 1666464484
transform 1 0 63020 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_685
timestamp 1666464484
transform 1 0 64124 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_697
timestamp 1666464484
transform 1 0 65228 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_709
timestamp 1666464484
transform 1 0 66332 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_721
timestamp 1666464484
transform 1 0 67436 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_727
timestamp 1666464484
transform 1 0 67988 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_729
timestamp 1666464484
transform 1 0 68172 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_741
timestamp 1666464484
transform 1 0 69276 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_753
timestamp 1666464484
transform 1 0 70380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_765
timestamp 1666464484
transform 1 0 71484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_777
timestamp 1666464484
transform 1 0 72588 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_783
timestamp 1666464484
transform 1 0 73140 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_785
timestamp 1666464484
transform 1 0 73324 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_797
timestamp 1666464484
transform 1 0 74428 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_809
timestamp 1666464484
transform 1 0 75532 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_821
timestamp 1666464484
transform 1 0 76636 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_833
timestamp 1666464484
transform 1 0 77740 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_839
timestamp 1666464484
transform 1 0 78292 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_841
timestamp 1666464484
transform 1 0 78476 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_853
timestamp 1666464484
transform 1 0 79580 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_865
timestamp 1666464484
transform 1 0 80684 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_877
timestamp 1666464484
transform 1 0 81788 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_889
timestamp 1666464484
transform 1 0 82892 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_895
timestamp 1666464484
transform 1 0 83444 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_897
timestamp 1666464484
transform 1 0 83628 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_909
timestamp 1666464484
transform 1 0 84732 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_921
timestamp 1666464484
transform 1 0 85836 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_933
timestamp 1666464484
transform 1 0 86940 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_945
timestamp 1666464484
transform 1 0 88044 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_951
timestamp 1666464484
transform 1 0 88596 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_953
timestamp 1666464484
transform 1 0 88780 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_965
timestamp 1666464484
transform 1 0 89884 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_977
timestamp 1666464484
transform 1 0 90988 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_989
timestamp 1666464484
transform 1 0 92092 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1001
timestamp 1666464484
transform 1 0 93196 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1007
timestamp 1666464484
transform 1 0 93748 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1009
timestamp 1666464484
transform 1 0 93932 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1021
timestamp 1666464484
transform 1 0 95036 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1033
timestamp 1666464484
transform 1 0 96140 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1045
timestamp 1666464484
transform 1 0 97244 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1057
timestamp 1666464484
transform 1 0 98348 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1063
timestamp 1666464484
transform 1 0 98900 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1065
timestamp 1666464484
transform 1 0 99084 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1077
timestamp 1666464484
transform 1 0 100188 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1089
timestamp 1666464484
transform 1 0 101292 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1101
timestamp 1666464484
transform 1 0 102396 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1113
timestamp 1666464484
transform 1 0 103500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1119
timestamp 1666464484
transform 1 0 104052 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1121
timestamp 1666464484
transform 1 0 104236 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1133
timestamp 1666464484
transform 1 0 105340 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1145
timestamp 1666464484
transform 1 0 106444 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1157
timestamp 1666464484
transform 1 0 107548 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1169
timestamp 1666464484
transform 1 0 108652 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1175
timestamp 1666464484
transform 1 0 109204 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1177
timestamp 1666464484
transform 1 0 109388 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1189
timestamp 1666464484
transform 1 0 110492 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1201
timestamp 1666464484
transform 1 0 111596 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1213
timestamp 1666464484
transform 1 0 112700 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1225
timestamp 1666464484
transform 1 0 113804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1231
timestamp 1666464484
transform 1 0 114356 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1233
timestamp 1666464484
transform 1 0 114540 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1245
timestamp 1666464484
transform 1 0 115644 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1257
timestamp 1666464484
transform 1 0 116748 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1269
timestamp 1666464484
transform 1 0 117852 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1281
timestamp 1666464484
transform 1 0 118956 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1287
timestamp 1666464484
transform 1 0 119508 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1289
timestamp 1666464484
transform 1 0 119692 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1301
timestamp 1666464484
transform 1 0 120796 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1313
timestamp 1666464484
transform 1 0 121900 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1325
timestamp 1666464484
transform 1 0 123004 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1337
timestamp 1666464484
transform 1 0 124108 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1343
timestamp 1666464484
transform 1 0 124660 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1345
timestamp 1666464484
transform 1 0 124844 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1357
timestamp 1666464484
transform 1 0 125948 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1369
timestamp 1666464484
transform 1 0 127052 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1381
timestamp 1666464484
transform 1 0 128156 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1393
timestamp 1666464484
transform 1 0 129260 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1399
timestamp 1666464484
transform 1 0 129812 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1401
timestamp 1666464484
transform 1 0 129996 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1413
timestamp 1666464484
transform 1 0 131100 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1425
timestamp 1666464484
transform 1 0 132204 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1437
timestamp 1666464484
transform 1 0 133308 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1449
timestamp 1666464484
transform 1 0 134412 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1455
timestamp 1666464484
transform 1 0 134964 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1457
timestamp 1666464484
transform 1 0 135148 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1469
timestamp 1666464484
transform 1 0 136252 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1481
timestamp 1666464484
transform 1 0 137356 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1493
timestamp 1666464484
transform 1 0 138460 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1505
timestamp 1666464484
transform 1 0 139564 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1511
timestamp 1666464484
transform 1 0 140116 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1513
timestamp 1666464484
transform 1 0 140300 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1525
timestamp 1666464484
transform 1 0 141404 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1537
timestamp 1666464484
transform 1 0 142508 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1549
timestamp 1666464484
transform 1 0 143612 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1561
timestamp 1666464484
transform 1 0 144716 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1567
timestamp 1666464484
transform 1 0 145268 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1569
timestamp 1666464484
transform 1 0 145452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1581
timestamp 1666464484
transform 1 0 146556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_1593
timestamp 1666464484
transform 1 0 147660 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_1601
timestamp 1666464484
transform 1 0 148396 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1666464484
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1666464484
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1666464484
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1666464484
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1666464484
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1666464484
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1666464484
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1666464484
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1666464484
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1666464484
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1666464484
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1666464484
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1666464484
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1666464484
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1666464484
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1666464484
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1666464484
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1666464484
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1666464484
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1666464484
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1666464484
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1666464484
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1666464484
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1666464484
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1666464484
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1666464484
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1666464484
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1666464484
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1666464484
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1666464484
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1666464484
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1666464484
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1666464484
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1666464484
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1666464484
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1666464484
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1666464484
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1666464484
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1666464484
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1666464484
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1666464484
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1666464484
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1666464484
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1666464484
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1666464484
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1666464484
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1666464484
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1666464484
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1666464484
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1666464484
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1666464484
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1666464484
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1666464484
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1666464484
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1666464484
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_557
timestamp 1666464484
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_569
timestamp 1666464484
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1666464484
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1666464484
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1666464484
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1666464484
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_613
timestamp 1666464484
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_625
timestamp 1666464484
transform 1 0 58604 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_637
timestamp 1666464484
transform 1 0 59708 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_643
timestamp 1666464484
transform 1 0 60260 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_645
timestamp 1666464484
transform 1 0 60444 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_657
timestamp 1666464484
transform 1 0 61548 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_669
timestamp 1666464484
transform 1 0 62652 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_681
timestamp 1666464484
transform 1 0 63756 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_693
timestamp 1666464484
transform 1 0 64860 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_699
timestamp 1666464484
transform 1 0 65412 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_701
timestamp 1666464484
transform 1 0 65596 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_713
timestamp 1666464484
transform 1 0 66700 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_725
timestamp 1666464484
transform 1 0 67804 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_737
timestamp 1666464484
transform 1 0 68908 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_749
timestamp 1666464484
transform 1 0 70012 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_755
timestamp 1666464484
transform 1 0 70564 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_757
timestamp 1666464484
transform 1 0 70748 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_769
timestamp 1666464484
transform 1 0 71852 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_781
timestamp 1666464484
transform 1 0 72956 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_793
timestamp 1666464484
transform 1 0 74060 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_805
timestamp 1666464484
transform 1 0 75164 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_811
timestamp 1666464484
transform 1 0 75716 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_813
timestamp 1666464484
transform 1 0 75900 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_825
timestamp 1666464484
transform 1 0 77004 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_837
timestamp 1666464484
transform 1 0 78108 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_849
timestamp 1666464484
transform 1 0 79212 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_861
timestamp 1666464484
transform 1 0 80316 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_867
timestamp 1666464484
transform 1 0 80868 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_869
timestamp 1666464484
transform 1 0 81052 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_881
timestamp 1666464484
transform 1 0 82156 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_893
timestamp 1666464484
transform 1 0 83260 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_905
timestamp 1666464484
transform 1 0 84364 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_917
timestamp 1666464484
transform 1 0 85468 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_923
timestamp 1666464484
transform 1 0 86020 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_925
timestamp 1666464484
transform 1 0 86204 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_937
timestamp 1666464484
transform 1 0 87308 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_949
timestamp 1666464484
transform 1 0 88412 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_961
timestamp 1666464484
transform 1 0 89516 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_973
timestamp 1666464484
transform 1 0 90620 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_979
timestamp 1666464484
transform 1 0 91172 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_981
timestamp 1666464484
transform 1 0 91356 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_993
timestamp 1666464484
transform 1 0 92460 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1005
timestamp 1666464484
transform 1 0 93564 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1017
timestamp 1666464484
transform 1 0 94668 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1029
timestamp 1666464484
transform 1 0 95772 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1035
timestamp 1666464484
transform 1 0 96324 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1037
timestamp 1666464484
transform 1 0 96508 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1049
timestamp 1666464484
transform 1 0 97612 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1061
timestamp 1666464484
transform 1 0 98716 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1073
timestamp 1666464484
transform 1 0 99820 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1085
timestamp 1666464484
transform 1 0 100924 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1091
timestamp 1666464484
transform 1 0 101476 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1093
timestamp 1666464484
transform 1 0 101660 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1105
timestamp 1666464484
transform 1 0 102764 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1117
timestamp 1666464484
transform 1 0 103868 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1129
timestamp 1666464484
transform 1 0 104972 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1141
timestamp 1666464484
transform 1 0 106076 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1147
timestamp 1666464484
transform 1 0 106628 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1149
timestamp 1666464484
transform 1 0 106812 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1161
timestamp 1666464484
transform 1 0 107916 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1173
timestamp 1666464484
transform 1 0 109020 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1185
timestamp 1666464484
transform 1 0 110124 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1197
timestamp 1666464484
transform 1 0 111228 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1203
timestamp 1666464484
transform 1 0 111780 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1205
timestamp 1666464484
transform 1 0 111964 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1217
timestamp 1666464484
transform 1 0 113068 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1229
timestamp 1666464484
transform 1 0 114172 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1241
timestamp 1666464484
transform 1 0 115276 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1253
timestamp 1666464484
transform 1 0 116380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1259
timestamp 1666464484
transform 1 0 116932 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1261
timestamp 1666464484
transform 1 0 117116 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1273
timestamp 1666464484
transform 1 0 118220 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1285
timestamp 1666464484
transform 1 0 119324 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1297
timestamp 1666464484
transform 1 0 120428 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1309
timestamp 1666464484
transform 1 0 121532 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1315
timestamp 1666464484
transform 1 0 122084 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1317
timestamp 1666464484
transform 1 0 122268 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1329
timestamp 1666464484
transform 1 0 123372 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1341
timestamp 1666464484
transform 1 0 124476 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1353
timestamp 1666464484
transform 1 0 125580 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1365
timestamp 1666464484
transform 1 0 126684 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1371
timestamp 1666464484
transform 1 0 127236 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1373
timestamp 1666464484
transform 1 0 127420 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1385
timestamp 1666464484
transform 1 0 128524 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1397
timestamp 1666464484
transform 1 0 129628 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1409
timestamp 1666464484
transform 1 0 130732 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1421
timestamp 1666464484
transform 1 0 131836 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1427
timestamp 1666464484
transform 1 0 132388 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1429
timestamp 1666464484
transform 1 0 132572 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1441
timestamp 1666464484
transform 1 0 133676 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1453
timestamp 1666464484
transform 1 0 134780 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1465
timestamp 1666464484
transform 1 0 135884 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1477
timestamp 1666464484
transform 1 0 136988 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1483
timestamp 1666464484
transform 1 0 137540 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1485
timestamp 1666464484
transform 1 0 137724 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1497
timestamp 1666464484
transform 1 0 138828 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1509
timestamp 1666464484
transform 1 0 139932 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1521
timestamp 1666464484
transform 1 0 141036 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1533
timestamp 1666464484
transform 1 0 142140 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1539
timestamp 1666464484
transform 1 0 142692 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1541
timestamp 1666464484
transform 1 0 142876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1553
timestamp 1666464484
transform 1 0 143980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1565
timestamp 1666464484
transform 1 0 145084 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1577
timestamp 1666464484
transform 1 0 146188 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1589
timestamp 1666464484
transform 1 0 147292 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1595
timestamp 1666464484
transform 1 0 147844 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1597
timestamp 1666464484
transform 1 0 148028 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1666464484
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1666464484
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1666464484
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1666464484
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1666464484
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1666464484
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1666464484
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1666464484
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1666464484
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1666464484
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1666464484
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1666464484
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1666464484
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1666464484
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1666464484
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1666464484
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1666464484
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1666464484
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1666464484
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1666464484
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1666464484
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1666464484
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1666464484
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1666464484
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1666464484
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1666464484
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1666464484
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1666464484
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1666464484
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1666464484
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1666464484
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1666464484
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1666464484
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1666464484
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1666464484
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1666464484
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1666464484
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1666464484
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1666464484
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1666464484
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1666464484
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1666464484
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1666464484
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1666464484
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1666464484
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1666464484
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1666464484
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1666464484
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1666464484
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1666464484
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1666464484
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1666464484
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1666464484
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1666464484
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1666464484
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1666464484
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1666464484
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1666464484
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1666464484
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1666464484
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_573
timestamp 1666464484
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1666464484
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_597
timestamp 1666464484
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1666464484
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1666464484
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_617
timestamp 1666464484
transform 1 0 57868 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_629
timestamp 1666464484
transform 1 0 58972 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_641
timestamp 1666464484
transform 1 0 60076 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_653
timestamp 1666464484
transform 1 0 61180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_665
timestamp 1666464484
transform 1 0 62284 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_671
timestamp 1666464484
transform 1 0 62836 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_673
timestamp 1666464484
transform 1 0 63020 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_685
timestamp 1666464484
transform 1 0 64124 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_697
timestamp 1666464484
transform 1 0 65228 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_709
timestamp 1666464484
transform 1 0 66332 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_721
timestamp 1666464484
transform 1 0 67436 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_727
timestamp 1666464484
transform 1 0 67988 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_729
timestamp 1666464484
transform 1 0 68172 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_741
timestamp 1666464484
transform 1 0 69276 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_753
timestamp 1666464484
transform 1 0 70380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_765
timestamp 1666464484
transform 1 0 71484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_777
timestamp 1666464484
transform 1 0 72588 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_783
timestamp 1666464484
transform 1 0 73140 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_785
timestamp 1666464484
transform 1 0 73324 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_797
timestamp 1666464484
transform 1 0 74428 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_809
timestamp 1666464484
transform 1 0 75532 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_821
timestamp 1666464484
transform 1 0 76636 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_833
timestamp 1666464484
transform 1 0 77740 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_839
timestamp 1666464484
transform 1 0 78292 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_841
timestamp 1666464484
transform 1 0 78476 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_853
timestamp 1666464484
transform 1 0 79580 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_865
timestamp 1666464484
transform 1 0 80684 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_877
timestamp 1666464484
transform 1 0 81788 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_889
timestamp 1666464484
transform 1 0 82892 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_895
timestamp 1666464484
transform 1 0 83444 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_897
timestamp 1666464484
transform 1 0 83628 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_909
timestamp 1666464484
transform 1 0 84732 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_921
timestamp 1666464484
transform 1 0 85836 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_933
timestamp 1666464484
transform 1 0 86940 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_945
timestamp 1666464484
transform 1 0 88044 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_951
timestamp 1666464484
transform 1 0 88596 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_953
timestamp 1666464484
transform 1 0 88780 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_965
timestamp 1666464484
transform 1 0 89884 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_977
timestamp 1666464484
transform 1 0 90988 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_989
timestamp 1666464484
transform 1 0 92092 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1001
timestamp 1666464484
transform 1 0 93196 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1007
timestamp 1666464484
transform 1 0 93748 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1009
timestamp 1666464484
transform 1 0 93932 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1021
timestamp 1666464484
transform 1 0 95036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1033
timestamp 1666464484
transform 1 0 96140 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1045
timestamp 1666464484
transform 1 0 97244 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1057
timestamp 1666464484
transform 1 0 98348 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1063
timestamp 1666464484
transform 1 0 98900 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1065
timestamp 1666464484
transform 1 0 99084 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1077
timestamp 1666464484
transform 1 0 100188 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1089
timestamp 1666464484
transform 1 0 101292 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1101
timestamp 1666464484
transform 1 0 102396 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1113
timestamp 1666464484
transform 1 0 103500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1119
timestamp 1666464484
transform 1 0 104052 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1121
timestamp 1666464484
transform 1 0 104236 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1133
timestamp 1666464484
transform 1 0 105340 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1145
timestamp 1666464484
transform 1 0 106444 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1157
timestamp 1666464484
transform 1 0 107548 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1169
timestamp 1666464484
transform 1 0 108652 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1175
timestamp 1666464484
transform 1 0 109204 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1177
timestamp 1666464484
transform 1 0 109388 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1189
timestamp 1666464484
transform 1 0 110492 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1201
timestamp 1666464484
transform 1 0 111596 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1213
timestamp 1666464484
transform 1 0 112700 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1225
timestamp 1666464484
transform 1 0 113804 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1231
timestamp 1666464484
transform 1 0 114356 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1233
timestamp 1666464484
transform 1 0 114540 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1245
timestamp 1666464484
transform 1 0 115644 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1257
timestamp 1666464484
transform 1 0 116748 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1269
timestamp 1666464484
transform 1 0 117852 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1281
timestamp 1666464484
transform 1 0 118956 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1287
timestamp 1666464484
transform 1 0 119508 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1289
timestamp 1666464484
transform 1 0 119692 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1301
timestamp 1666464484
transform 1 0 120796 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1313
timestamp 1666464484
transform 1 0 121900 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1325
timestamp 1666464484
transform 1 0 123004 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1337
timestamp 1666464484
transform 1 0 124108 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1343
timestamp 1666464484
transform 1 0 124660 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1345
timestamp 1666464484
transform 1 0 124844 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1357
timestamp 1666464484
transform 1 0 125948 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1369
timestamp 1666464484
transform 1 0 127052 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1381
timestamp 1666464484
transform 1 0 128156 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1393
timestamp 1666464484
transform 1 0 129260 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1399
timestamp 1666464484
transform 1 0 129812 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1401
timestamp 1666464484
transform 1 0 129996 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1413
timestamp 1666464484
transform 1 0 131100 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1425
timestamp 1666464484
transform 1 0 132204 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1437
timestamp 1666464484
transform 1 0 133308 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1449
timestamp 1666464484
transform 1 0 134412 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1455
timestamp 1666464484
transform 1 0 134964 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1457
timestamp 1666464484
transform 1 0 135148 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1469
timestamp 1666464484
transform 1 0 136252 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1481
timestamp 1666464484
transform 1 0 137356 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1493
timestamp 1666464484
transform 1 0 138460 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1505
timestamp 1666464484
transform 1 0 139564 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1511
timestamp 1666464484
transform 1 0 140116 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1513
timestamp 1666464484
transform 1 0 140300 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1525
timestamp 1666464484
transform 1 0 141404 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1537
timestamp 1666464484
transform 1 0 142508 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1549
timestamp 1666464484
transform 1 0 143612 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1561
timestamp 1666464484
transform 1 0 144716 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1567
timestamp 1666464484
transform 1 0 145268 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1569
timestamp 1666464484
transform 1 0 145452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1581
timestamp 1666464484
transform 1 0 146556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_1593
timestamp 1666464484
transform 1 0 147660 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_1601
timestamp 1666464484
transform 1 0 148396 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1666464484
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1666464484
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1666464484
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1666464484
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1666464484
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1666464484
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1666464484
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1666464484
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1666464484
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1666464484
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1666464484
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1666464484
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1666464484
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1666464484
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1666464484
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1666464484
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1666464484
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1666464484
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1666464484
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1666464484
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1666464484
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1666464484
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1666464484
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1666464484
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1666464484
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1666464484
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1666464484
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1666464484
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1666464484
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1666464484
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1666464484
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1666464484
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1666464484
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1666464484
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1666464484
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1666464484
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1666464484
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1666464484
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1666464484
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1666464484
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1666464484
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1666464484
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1666464484
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1666464484
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1666464484
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1666464484
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1666464484
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1666464484
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1666464484
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1666464484
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1666464484
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1666464484
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1666464484
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1666464484
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1666464484
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1666464484
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1666464484
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1666464484
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1666464484
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_569
timestamp 1666464484
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1666464484
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1666464484
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1666464484
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_601
timestamp 1666464484
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_613
timestamp 1666464484
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_625
timestamp 1666464484
transform 1 0 58604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_637
timestamp 1666464484
transform 1 0 59708 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_643
timestamp 1666464484
transform 1 0 60260 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_645
timestamp 1666464484
transform 1 0 60444 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_657
timestamp 1666464484
transform 1 0 61548 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_669
timestamp 1666464484
transform 1 0 62652 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_681
timestamp 1666464484
transform 1 0 63756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_693
timestamp 1666464484
transform 1 0 64860 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_699
timestamp 1666464484
transform 1 0 65412 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_701
timestamp 1666464484
transform 1 0 65596 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_713
timestamp 1666464484
transform 1 0 66700 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_725
timestamp 1666464484
transform 1 0 67804 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_737
timestamp 1666464484
transform 1 0 68908 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_749
timestamp 1666464484
transform 1 0 70012 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_755
timestamp 1666464484
transform 1 0 70564 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_757
timestamp 1666464484
transform 1 0 70748 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_769
timestamp 1666464484
transform 1 0 71852 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_781
timestamp 1666464484
transform 1 0 72956 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_793
timestamp 1666464484
transform 1 0 74060 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_805
timestamp 1666464484
transform 1 0 75164 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_811
timestamp 1666464484
transform 1 0 75716 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_813
timestamp 1666464484
transform 1 0 75900 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_825
timestamp 1666464484
transform 1 0 77004 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_837
timestamp 1666464484
transform 1 0 78108 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_849
timestamp 1666464484
transform 1 0 79212 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_861
timestamp 1666464484
transform 1 0 80316 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_867
timestamp 1666464484
transform 1 0 80868 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_869
timestamp 1666464484
transform 1 0 81052 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_881
timestamp 1666464484
transform 1 0 82156 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_893
timestamp 1666464484
transform 1 0 83260 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_905
timestamp 1666464484
transform 1 0 84364 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_917
timestamp 1666464484
transform 1 0 85468 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_923
timestamp 1666464484
transform 1 0 86020 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_925
timestamp 1666464484
transform 1 0 86204 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_937
timestamp 1666464484
transform 1 0 87308 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_949
timestamp 1666464484
transform 1 0 88412 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_961
timestamp 1666464484
transform 1 0 89516 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_973
timestamp 1666464484
transform 1 0 90620 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_979
timestamp 1666464484
transform 1 0 91172 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_981
timestamp 1666464484
transform 1 0 91356 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_993
timestamp 1666464484
transform 1 0 92460 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1005
timestamp 1666464484
transform 1 0 93564 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1017
timestamp 1666464484
transform 1 0 94668 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1029
timestamp 1666464484
transform 1 0 95772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1035
timestamp 1666464484
transform 1 0 96324 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1037
timestamp 1666464484
transform 1 0 96508 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1049
timestamp 1666464484
transform 1 0 97612 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1061
timestamp 1666464484
transform 1 0 98716 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1073
timestamp 1666464484
transform 1 0 99820 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1085
timestamp 1666464484
transform 1 0 100924 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1091
timestamp 1666464484
transform 1 0 101476 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1093
timestamp 1666464484
transform 1 0 101660 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1105
timestamp 1666464484
transform 1 0 102764 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1117
timestamp 1666464484
transform 1 0 103868 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1129
timestamp 1666464484
transform 1 0 104972 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1141
timestamp 1666464484
transform 1 0 106076 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1147
timestamp 1666464484
transform 1 0 106628 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1149
timestamp 1666464484
transform 1 0 106812 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1161
timestamp 1666464484
transform 1 0 107916 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1173
timestamp 1666464484
transform 1 0 109020 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1185
timestamp 1666464484
transform 1 0 110124 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1197
timestamp 1666464484
transform 1 0 111228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1203
timestamp 1666464484
transform 1 0 111780 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1205
timestamp 1666464484
transform 1 0 111964 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1217
timestamp 1666464484
transform 1 0 113068 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1229
timestamp 1666464484
transform 1 0 114172 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1241
timestamp 1666464484
transform 1 0 115276 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1253
timestamp 1666464484
transform 1 0 116380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1259
timestamp 1666464484
transform 1 0 116932 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1261
timestamp 1666464484
transform 1 0 117116 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1273
timestamp 1666464484
transform 1 0 118220 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1285
timestamp 1666464484
transform 1 0 119324 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1297
timestamp 1666464484
transform 1 0 120428 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1309
timestamp 1666464484
transform 1 0 121532 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1315
timestamp 1666464484
transform 1 0 122084 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1317
timestamp 1666464484
transform 1 0 122268 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1329
timestamp 1666464484
transform 1 0 123372 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1341
timestamp 1666464484
transform 1 0 124476 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1353
timestamp 1666464484
transform 1 0 125580 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1365
timestamp 1666464484
transform 1 0 126684 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1371
timestamp 1666464484
transform 1 0 127236 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1373
timestamp 1666464484
transform 1 0 127420 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1385
timestamp 1666464484
transform 1 0 128524 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1397
timestamp 1666464484
transform 1 0 129628 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1409
timestamp 1666464484
transform 1 0 130732 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1421
timestamp 1666464484
transform 1 0 131836 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1427
timestamp 1666464484
transform 1 0 132388 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1429
timestamp 1666464484
transform 1 0 132572 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1441
timestamp 1666464484
transform 1 0 133676 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1453
timestamp 1666464484
transform 1 0 134780 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1465
timestamp 1666464484
transform 1 0 135884 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1477
timestamp 1666464484
transform 1 0 136988 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1483
timestamp 1666464484
transform 1 0 137540 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1485
timestamp 1666464484
transform 1 0 137724 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1497
timestamp 1666464484
transform 1 0 138828 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1509
timestamp 1666464484
transform 1 0 139932 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1521
timestamp 1666464484
transform 1 0 141036 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1533
timestamp 1666464484
transform 1 0 142140 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1539
timestamp 1666464484
transform 1 0 142692 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1541
timestamp 1666464484
transform 1 0 142876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1553
timestamp 1666464484
transform 1 0 143980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1565
timestamp 1666464484
transform 1 0 145084 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1577
timestamp 1666464484
transform 1 0 146188 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1589
timestamp 1666464484
transform 1 0 147292 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1595
timestamp 1666464484
transform 1 0 147844 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1597
timestamp 1666464484
transform 1 0 148028 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1666464484
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1666464484
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1666464484
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1666464484
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1666464484
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1666464484
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1666464484
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1666464484
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1666464484
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1666464484
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1666464484
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1666464484
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1666464484
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1666464484
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1666464484
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1666464484
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1666464484
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1666464484
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1666464484
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1666464484
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1666464484
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1666464484
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1666464484
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1666464484
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1666464484
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1666464484
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1666464484
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1666464484
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1666464484
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1666464484
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1666464484
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1666464484
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1666464484
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1666464484
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1666464484
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1666464484
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1666464484
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1666464484
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1666464484
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1666464484
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1666464484
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1666464484
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1666464484
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1666464484
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1666464484
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1666464484
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1666464484
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1666464484
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1666464484
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1666464484
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1666464484
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1666464484
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1666464484
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1666464484
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1666464484
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1666464484
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1666464484
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1666464484
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1666464484
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1666464484
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1666464484
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_585
timestamp 1666464484
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_597
timestamp 1666464484
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1666464484
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1666464484
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_617
timestamp 1666464484
transform 1 0 57868 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_629
timestamp 1666464484
transform 1 0 58972 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_641
timestamp 1666464484
transform 1 0 60076 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_653
timestamp 1666464484
transform 1 0 61180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_665
timestamp 1666464484
transform 1 0 62284 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_671
timestamp 1666464484
transform 1 0 62836 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_673
timestamp 1666464484
transform 1 0 63020 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_685
timestamp 1666464484
transform 1 0 64124 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_697
timestamp 1666464484
transform 1 0 65228 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_709
timestamp 1666464484
transform 1 0 66332 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_721
timestamp 1666464484
transform 1 0 67436 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_727
timestamp 1666464484
transform 1 0 67988 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_729
timestamp 1666464484
transform 1 0 68172 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_741
timestamp 1666464484
transform 1 0 69276 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_753
timestamp 1666464484
transform 1 0 70380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_765
timestamp 1666464484
transform 1 0 71484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_777
timestamp 1666464484
transform 1 0 72588 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_783
timestamp 1666464484
transform 1 0 73140 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_785
timestamp 1666464484
transform 1 0 73324 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_797
timestamp 1666464484
transform 1 0 74428 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_809
timestamp 1666464484
transform 1 0 75532 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_821
timestamp 1666464484
transform 1 0 76636 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_833
timestamp 1666464484
transform 1 0 77740 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_839
timestamp 1666464484
transform 1 0 78292 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_841
timestamp 1666464484
transform 1 0 78476 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_853
timestamp 1666464484
transform 1 0 79580 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_865
timestamp 1666464484
transform 1 0 80684 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_877
timestamp 1666464484
transform 1 0 81788 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_889
timestamp 1666464484
transform 1 0 82892 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_895
timestamp 1666464484
transform 1 0 83444 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_897
timestamp 1666464484
transform 1 0 83628 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_909
timestamp 1666464484
transform 1 0 84732 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_921
timestamp 1666464484
transform 1 0 85836 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_933
timestamp 1666464484
transform 1 0 86940 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_945
timestamp 1666464484
transform 1 0 88044 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_951
timestamp 1666464484
transform 1 0 88596 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_953
timestamp 1666464484
transform 1 0 88780 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_965
timestamp 1666464484
transform 1 0 89884 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_977
timestamp 1666464484
transform 1 0 90988 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_989
timestamp 1666464484
transform 1 0 92092 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1001
timestamp 1666464484
transform 1 0 93196 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1007
timestamp 1666464484
transform 1 0 93748 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1009
timestamp 1666464484
transform 1 0 93932 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1021
timestamp 1666464484
transform 1 0 95036 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1033
timestamp 1666464484
transform 1 0 96140 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1045
timestamp 1666464484
transform 1 0 97244 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1057
timestamp 1666464484
transform 1 0 98348 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1063
timestamp 1666464484
transform 1 0 98900 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1065
timestamp 1666464484
transform 1 0 99084 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1077
timestamp 1666464484
transform 1 0 100188 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1089
timestamp 1666464484
transform 1 0 101292 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1101
timestamp 1666464484
transform 1 0 102396 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1113
timestamp 1666464484
transform 1 0 103500 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1119
timestamp 1666464484
transform 1 0 104052 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1121
timestamp 1666464484
transform 1 0 104236 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1133
timestamp 1666464484
transform 1 0 105340 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1145
timestamp 1666464484
transform 1 0 106444 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1157
timestamp 1666464484
transform 1 0 107548 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1169
timestamp 1666464484
transform 1 0 108652 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1175
timestamp 1666464484
transform 1 0 109204 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1177
timestamp 1666464484
transform 1 0 109388 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1189
timestamp 1666464484
transform 1 0 110492 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1201
timestamp 1666464484
transform 1 0 111596 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1213
timestamp 1666464484
transform 1 0 112700 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1225
timestamp 1666464484
transform 1 0 113804 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1231
timestamp 1666464484
transform 1 0 114356 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1233
timestamp 1666464484
transform 1 0 114540 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1245
timestamp 1666464484
transform 1 0 115644 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1257
timestamp 1666464484
transform 1 0 116748 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1269
timestamp 1666464484
transform 1 0 117852 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1281
timestamp 1666464484
transform 1 0 118956 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1287
timestamp 1666464484
transform 1 0 119508 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1289
timestamp 1666464484
transform 1 0 119692 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1301
timestamp 1666464484
transform 1 0 120796 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1313
timestamp 1666464484
transform 1 0 121900 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1325
timestamp 1666464484
transform 1 0 123004 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1337
timestamp 1666464484
transform 1 0 124108 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1343
timestamp 1666464484
transform 1 0 124660 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1345
timestamp 1666464484
transform 1 0 124844 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1357
timestamp 1666464484
transform 1 0 125948 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1369
timestamp 1666464484
transform 1 0 127052 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1381
timestamp 1666464484
transform 1 0 128156 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1393
timestamp 1666464484
transform 1 0 129260 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1399
timestamp 1666464484
transform 1 0 129812 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1401
timestamp 1666464484
transform 1 0 129996 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1413
timestamp 1666464484
transform 1 0 131100 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1425
timestamp 1666464484
transform 1 0 132204 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1437
timestamp 1666464484
transform 1 0 133308 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1449
timestamp 1666464484
transform 1 0 134412 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1455
timestamp 1666464484
transform 1 0 134964 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1457
timestamp 1666464484
transform 1 0 135148 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1469
timestamp 1666464484
transform 1 0 136252 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1481
timestamp 1666464484
transform 1 0 137356 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1493
timestamp 1666464484
transform 1 0 138460 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1505
timestamp 1666464484
transform 1 0 139564 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1511
timestamp 1666464484
transform 1 0 140116 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1513
timestamp 1666464484
transform 1 0 140300 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1525
timestamp 1666464484
transform 1 0 141404 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1537
timestamp 1666464484
transform 1 0 142508 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1549
timestamp 1666464484
transform 1 0 143612 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1561
timestamp 1666464484
transform 1 0 144716 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1567
timestamp 1666464484
transform 1 0 145268 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1569
timestamp 1666464484
transform 1 0 145452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1581
timestamp 1666464484
transform 1 0 146556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_1593
timestamp 1666464484
transform 1 0 147660 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_1601
timestamp 1666464484
transform 1 0 148396 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1666464484
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1666464484
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1666464484
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1666464484
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1666464484
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1666464484
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1666464484
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1666464484
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1666464484
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1666464484
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1666464484
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1666464484
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1666464484
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1666464484
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1666464484
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1666464484
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1666464484
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1666464484
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1666464484
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1666464484
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1666464484
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1666464484
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1666464484
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1666464484
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1666464484
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1666464484
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1666464484
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1666464484
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1666464484
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1666464484
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1666464484
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1666464484
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1666464484
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1666464484
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1666464484
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1666464484
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1666464484
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1666464484
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1666464484
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1666464484
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1666464484
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1666464484
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1666464484
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1666464484
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1666464484
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1666464484
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1666464484
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1666464484
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1666464484
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1666464484
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1666464484
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1666464484
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1666464484
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1666464484
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1666464484
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1666464484
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1666464484
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1666464484
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_545
timestamp 1666464484
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_557
timestamp 1666464484
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_569
timestamp 1666464484
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1666464484
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1666464484
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_589
timestamp 1666464484
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_601
timestamp 1666464484
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_613
timestamp 1666464484
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_625
timestamp 1666464484
transform 1 0 58604 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_637
timestamp 1666464484
transform 1 0 59708 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_643
timestamp 1666464484
transform 1 0 60260 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_645
timestamp 1666464484
transform 1 0 60444 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_657
timestamp 1666464484
transform 1 0 61548 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_669
timestamp 1666464484
transform 1 0 62652 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_681
timestamp 1666464484
transform 1 0 63756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_693
timestamp 1666464484
transform 1 0 64860 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_699
timestamp 1666464484
transform 1 0 65412 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_701
timestamp 1666464484
transform 1 0 65596 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_713
timestamp 1666464484
transform 1 0 66700 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_725
timestamp 1666464484
transform 1 0 67804 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_737
timestamp 1666464484
transform 1 0 68908 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_749
timestamp 1666464484
transform 1 0 70012 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_755
timestamp 1666464484
transform 1 0 70564 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_757
timestamp 1666464484
transform 1 0 70748 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_769
timestamp 1666464484
transform 1 0 71852 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_781
timestamp 1666464484
transform 1 0 72956 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_793
timestamp 1666464484
transform 1 0 74060 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_805
timestamp 1666464484
transform 1 0 75164 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_811
timestamp 1666464484
transform 1 0 75716 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_813
timestamp 1666464484
transform 1 0 75900 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_825
timestamp 1666464484
transform 1 0 77004 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_837
timestamp 1666464484
transform 1 0 78108 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_849
timestamp 1666464484
transform 1 0 79212 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_861
timestamp 1666464484
transform 1 0 80316 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_867
timestamp 1666464484
transform 1 0 80868 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_869
timestamp 1666464484
transform 1 0 81052 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_881
timestamp 1666464484
transform 1 0 82156 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_893
timestamp 1666464484
transform 1 0 83260 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_905
timestamp 1666464484
transform 1 0 84364 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_917
timestamp 1666464484
transform 1 0 85468 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_923
timestamp 1666464484
transform 1 0 86020 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_925
timestamp 1666464484
transform 1 0 86204 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_937
timestamp 1666464484
transform 1 0 87308 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_949
timestamp 1666464484
transform 1 0 88412 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_961
timestamp 1666464484
transform 1 0 89516 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_973
timestamp 1666464484
transform 1 0 90620 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_979
timestamp 1666464484
transform 1 0 91172 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_981
timestamp 1666464484
transform 1 0 91356 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_993
timestamp 1666464484
transform 1 0 92460 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1005
timestamp 1666464484
transform 1 0 93564 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1017
timestamp 1666464484
transform 1 0 94668 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1029
timestamp 1666464484
transform 1 0 95772 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1035
timestamp 1666464484
transform 1 0 96324 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1037
timestamp 1666464484
transform 1 0 96508 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1049
timestamp 1666464484
transform 1 0 97612 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1061
timestamp 1666464484
transform 1 0 98716 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1073
timestamp 1666464484
transform 1 0 99820 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1085
timestamp 1666464484
transform 1 0 100924 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1091
timestamp 1666464484
transform 1 0 101476 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1093
timestamp 1666464484
transform 1 0 101660 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1105
timestamp 1666464484
transform 1 0 102764 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1117
timestamp 1666464484
transform 1 0 103868 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1129
timestamp 1666464484
transform 1 0 104972 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1141
timestamp 1666464484
transform 1 0 106076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1147
timestamp 1666464484
transform 1 0 106628 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1149
timestamp 1666464484
transform 1 0 106812 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1161
timestamp 1666464484
transform 1 0 107916 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1173
timestamp 1666464484
transform 1 0 109020 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1185
timestamp 1666464484
transform 1 0 110124 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1197
timestamp 1666464484
transform 1 0 111228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1203
timestamp 1666464484
transform 1 0 111780 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1205
timestamp 1666464484
transform 1 0 111964 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1217
timestamp 1666464484
transform 1 0 113068 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1229
timestamp 1666464484
transform 1 0 114172 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1241
timestamp 1666464484
transform 1 0 115276 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1253
timestamp 1666464484
transform 1 0 116380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1259
timestamp 1666464484
transform 1 0 116932 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1261
timestamp 1666464484
transform 1 0 117116 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1273
timestamp 1666464484
transform 1 0 118220 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1285
timestamp 1666464484
transform 1 0 119324 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1297
timestamp 1666464484
transform 1 0 120428 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1309
timestamp 1666464484
transform 1 0 121532 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1315
timestamp 1666464484
transform 1 0 122084 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1317
timestamp 1666464484
transform 1 0 122268 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1329
timestamp 1666464484
transform 1 0 123372 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1341
timestamp 1666464484
transform 1 0 124476 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1353
timestamp 1666464484
transform 1 0 125580 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1365
timestamp 1666464484
transform 1 0 126684 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1371
timestamp 1666464484
transform 1 0 127236 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1373
timestamp 1666464484
transform 1 0 127420 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1385
timestamp 1666464484
transform 1 0 128524 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1397
timestamp 1666464484
transform 1 0 129628 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1409
timestamp 1666464484
transform 1 0 130732 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1421
timestamp 1666464484
transform 1 0 131836 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1427
timestamp 1666464484
transform 1 0 132388 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1429
timestamp 1666464484
transform 1 0 132572 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1441
timestamp 1666464484
transform 1 0 133676 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1453
timestamp 1666464484
transform 1 0 134780 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1465
timestamp 1666464484
transform 1 0 135884 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1477
timestamp 1666464484
transform 1 0 136988 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1483
timestamp 1666464484
transform 1 0 137540 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1485
timestamp 1666464484
transform 1 0 137724 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1497
timestamp 1666464484
transform 1 0 138828 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1509
timestamp 1666464484
transform 1 0 139932 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1521
timestamp 1666464484
transform 1 0 141036 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1533
timestamp 1666464484
transform 1 0 142140 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1539
timestamp 1666464484
transform 1 0 142692 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1541
timestamp 1666464484
transform 1 0 142876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1553
timestamp 1666464484
transform 1 0 143980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1565
timestamp 1666464484
transform 1 0 145084 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1577
timestamp 1666464484
transform 1 0 146188 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1589
timestamp 1666464484
transform 1 0 147292 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1595
timestamp 1666464484
transform 1 0 147844 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1597
timestamp 1666464484
transform 1 0 148028 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1666464484
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1666464484
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1666464484
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1666464484
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1666464484
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1666464484
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1666464484
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1666464484
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1666464484
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1666464484
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1666464484
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1666464484
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1666464484
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1666464484
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1666464484
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1666464484
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1666464484
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1666464484
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1666464484
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1666464484
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1666464484
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1666464484
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1666464484
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1666464484
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1666464484
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1666464484
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1666464484
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1666464484
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1666464484
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1666464484
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1666464484
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1666464484
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1666464484
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1666464484
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1666464484
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1666464484
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1666464484
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1666464484
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1666464484
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1666464484
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1666464484
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1666464484
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1666464484
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1666464484
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1666464484
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1666464484
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1666464484
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1666464484
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1666464484
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1666464484
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1666464484
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1666464484
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1666464484
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1666464484
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1666464484
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1666464484
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1666464484
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1666464484
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1666464484
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1666464484
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1666464484
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_573
timestamp 1666464484
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_585
timestamp 1666464484
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_597
timestamp 1666464484
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1666464484
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1666464484
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_617
timestamp 1666464484
transform 1 0 57868 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_629
timestamp 1666464484
transform 1 0 58972 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_641
timestamp 1666464484
transform 1 0 60076 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_653
timestamp 1666464484
transform 1 0 61180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_665
timestamp 1666464484
transform 1 0 62284 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_671
timestamp 1666464484
transform 1 0 62836 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_673
timestamp 1666464484
transform 1 0 63020 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_685
timestamp 1666464484
transform 1 0 64124 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_697
timestamp 1666464484
transform 1 0 65228 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_709
timestamp 1666464484
transform 1 0 66332 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_721
timestamp 1666464484
transform 1 0 67436 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_727
timestamp 1666464484
transform 1 0 67988 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_729
timestamp 1666464484
transform 1 0 68172 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_741
timestamp 1666464484
transform 1 0 69276 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_753
timestamp 1666464484
transform 1 0 70380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_765
timestamp 1666464484
transform 1 0 71484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_777
timestamp 1666464484
transform 1 0 72588 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_783
timestamp 1666464484
transform 1 0 73140 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_785
timestamp 1666464484
transform 1 0 73324 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_797
timestamp 1666464484
transform 1 0 74428 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_809
timestamp 1666464484
transform 1 0 75532 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_821
timestamp 1666464484
transform 1 0 76636 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_833
timestamp 1666464484
transform 1 0 77740 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_839
timestamp 1666464484
transform 1 0 78292 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_841
timestamp 1666464484
transform 1 0 78476 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_853
timestamp 1666464484
transform 1 0 79580 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_865
timestamp 1666464484
transform 1 0 80684 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_877
timestamp 1666464484
transform 1 0 81788 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_889
timestamp 1666464484
transform 1 0 82892 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_895
timestamp 1666464484
transform 1 0 83444 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_897
timestamp 1666464484
transform 1 0 83628 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_909
timestamp 1666464484
transform 1 0 84732 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_921
timestamp 1666464484
transform 1 0 85836 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_933
timestamp 1666464484
transform 1 0 86940 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_945
timestamp 1666464484
transform 1 0 88044 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_951
timestamp 1666464484
transform 1 0 88596 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_953
timestamp 1666464484
transform 1 0 88780 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_965
timestamp 1666464484
transform 1 0 89884 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_977
timestamp 1666464484
transform 1 0 90988 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_989
timestamp 1666464484
transform 1 0 92092 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1001
timestamp 1666464484
transform 1 0 93196 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1007
timestamp 1666464484
transform 1 0 93748 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1009
timestamp 1666464484
transform 1 0 93932 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1021
timestamp 1666464484
transform 1 0 95036 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1033
timestamp 1666464484
transform 1 0 96140 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1045
timestamp 1666464484
transform 1 0 97244 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1057
timestamp 1666464484
transform 1 0 98348 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1063
timestamp 1666464484
transform 1 0 98900 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1065
timestamp 1666464484
transform 1 0 99084 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1077
timestamp 1666464484
transform 1 0 100188 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1089
timestamp 1666464484
transform 1 0 101292 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1101
timestamp 1666464484
transform 1 0 102396 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1113
timestamp 1666464484
transform 1 0 103500 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1119
timestamp 1666464484
transform 1 0 104052 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1121
timestamp 1666464484
transform 1 0 104236 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1133
timestamp 1666464484
transform 1 0 105340 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1145
timestamp 1666464484
transform 1 0 106444 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1157
timestamp 1666464484
transform 1 0 107548 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1169
timestamp 1666464484
transform 1 0 108652 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1175
timestamp 1666464484
transform 1 0 109204 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1177
timestamp 1666464484
transform 1 0 109388 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1189
timestamp 1666464484
transform 1 0 110492 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1201
timestamp 1666464484
transform 1 0 111596 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1213
timestamp 1666464484
transform 1 0 112700 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1225
timestamp 1666464484
transform 1 0 113804 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1231
timestamp 1666464484
transform 1 0 114356 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1233
timestamp 1666464484
transform 1 0 114540 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1245
timestamp 1666464484
transform 1 0 115644 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1257
timestamp 1666464484
transform 1 0 116748 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1269
timestamp 1666464484
transform 1 0 117852 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1281
timestamp 1666464484
transform 1 0 118956 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1287
timestamp 1666464484
transform 1 0 119508 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1289
timestamp 1666464484
transform 1 0 119692 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1301
timestamp 1666464484
transform 1 0 120796 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1313
timestamp 1666464484
transform 1 0 121900 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1325
timestamp 1666464484
transform 1 0 123004 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1337
timestamp 1666464484
transform 1 0 124108 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1343
timestamp 1666464484
transform 1 0 124660 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1345
timestamp 1666464484
transform 1 0 124844 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1357
timestamp 1666464484
transform 1 0 125948 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1369
timestamp 1666464484
transform 1 0 127052 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1381
timestamp 1666464484
transform 1 0 128156 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1393
timestamp 1666464484
transform 1 0 129260 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1399
timestamp 1666464484
transform 1 0 129812 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1401
timestamp 1666464484
transform 1 0 129996 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1413
timestamp 1666464484
transform 1 0 131100 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1425
timestamp 1666464484
transform 1 0 132204 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1437
timestamp 1666464484
transform 1 0 133308 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1449
timestamp 1666464484
transform 1 0 134412 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1455
timestamp 1666464484
transform 1 0 134964 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1457
timestamp 1666464484
transform 1 0 135148 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1469
timestamp 1666464484
transform 1 0 136252 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1481
timestamp 1666464484
transform 1 0 137356 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1493
timestamp 1666464484
transform 1 0 138460 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1505
timestamp 1666464484
transform 1 0 139564 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1511
timestamp 1666464484
transform 1 0 140116 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1513
timestamp 1666464484
transform 1 0 140300 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1525
timestamp 1666464484
transform 1 0 141404 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1537
timestamp 1666464484
transform 1 0 142508 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1549
timestamp 1666464484
transform 1 0 143612 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1561
timestamp 1666464484
transform 1 0 144716 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1567
timestamp 1666464484
transform 1 0 145268 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1569
timestamp 1666464484
transform 1 0 145452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1581
timestamp 1666464484
transform 1 0 146556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_1593
timestamp 1666464484
transform 1 0 147660 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_1601
timestamp 1666464484
transform 1 0 148396 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1666464484
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1666464484
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1666464484
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1666464484
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1666464484
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1666464484
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1666464484
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1666464484
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1666464484
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1666464484
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1666464484
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1666464484
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1666464484
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1666464484
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1666464484
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1666464484
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1666464484
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1666464484
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1666464484
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1666464484
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1666464484
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1666464484
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1666464484
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1666464484
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1666464484
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1666464484
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1666464484
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1666464484
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1666464484
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1666464484
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1666464484
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1666464484
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1666464484
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1666464484
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1666464484
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1666464484
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1666464484
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1666464484
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1666464484
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1666464484
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1666464484
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1666464484
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1666464484
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1666464484
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1666464484
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1666464484
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1666464484
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1666464484
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1666464484
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1666464484
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1666464484
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1666464484
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1666464484
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1666464484
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1666464484
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1666464484
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1666464484
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1666464484
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1666464484
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1666464484
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1666464484
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1666464484
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1666464484
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1666464484
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_601
timestamp 1666464484
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_613
timestamp 1666464484
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_625
timestamp 1666464484
transform 1 0 58604 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_637
timestamp 1666464484
transform 1 0 59708 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_643
timestamp 1666464484
transform 1 0 60260 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_645
timestamp 1666464484
transform 1 0 60444 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_657
timestamp 1666464484
transform 1 0 61548 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_669
timestamp 1666464484
transform 1 0 62652 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_681
timestamp 1666464484
transform 1 0 63756 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_693
timestamp 1666464484
transform 1 0 64860 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_699
timestamp 1666464484
transform 1 0 65412 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_701
timestamp 1666464484
transform 1 0 65596 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_713
timestamp 1666464484
transform 1 0 66700 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_725
timestamp 1666464484
transform 1 0 67804 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_737
timestamp 1666464484
transform 1 0 68908 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_749
timestamp 1666464484
transform 1 0 70012 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_755
timestamp 1666464484
transform 1 0 70564 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_757
timestamp 1666464484
transform 1 0 70748 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_769
timestamp 1666464484
transform 1 0 71852 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_781
timestamp 1666464484
transform 1 0 72956 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_793
timestamp 1666464484
transform 1 0 74060 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_805
timestamp 1666464484
transform 1 0 75164 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_811
timestamp 1666464484
transform 1 0 75716 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_813
timestamp 1666464484
transform 1 0 75900 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_825
timestamp 1666464484
transform 1 0 77004 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_837
timestamp 1666464484
transform 1 0 78108 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_849
timestamp 1666464484
transform 1 0 79212 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_861
timestamp 1666464484
transform 1 0 80316 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_867
timestamp 1666464484
transform 1 0 80868 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_869
timestamp 1666464484
transform 1 0 81052 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_881
timestamp 1666464484
transform 1 0 82156 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_893
timestamp 1666464484
transform 1 0 83260 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_905
timestamp 1666464484
transform 1 0 84364 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_917
timestamp 1666464484
transform 1 0 85468 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_923
timestamp 1666464484
transform 1 0 86020 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_925
timestamp 1666464484
transform 1 0 86204 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_937
timestamp 1666464484
transform 1 0 87308 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_949
timestamp 1666464484
transform 1 0 88412 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_961
timestamp 1666464484
transform 1 0 89516 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_973
timestamp 1666464484
transform 1 0 90620 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_979
timestamp 1666464484
transform 1 0 91172 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_981
timestamp 1666464484
transform 1 0 91356 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_993
timestamp 1666464484
transform 1 0 92460 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1005
timestamp 1666464484
transform 1 0 93564 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1017
timestamp 1666464484
transform 1 0 94668 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1029
timestamp 1666464484
transform 1 0 95772 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1035
timestamp 1666464484
transform 1 0 96324 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1037
timestamp 1666464484
transform 1 0 96508 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1049
timestamp 1666464484
transform 1 0 97612 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1061
timestamp 1666464484
transform 1 0 98716 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1073
timestamp 1666464484
transform 1 0 99820 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1085
timestamp 1666464484
transform 1 0 100924 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1091
timestamp 1666464484
transform 1 0 101476 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1093
timestamp 1666464484
transform 1 0 101660 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1105
timestamp 1666464484
transform 1 0 102764 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1117
timestamp 1666464484
transform 1 0 103868 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1129
timestamp 1666464484
transform 1 0 104972 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1141
timestamp 1666464484
transform 1 0 106076 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1147
timestamp 1666464484
transform 1 0 106628 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1149
timestamp 1666464484
transform 1 0 106812 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1161
timestamp 1666464484
transform 1 0 107916 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1173
timestamp 1666464484
transform 1 0 109020 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1185
timestamp 1666464484
transform 1 0 110124 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1197
timestamp 1666464484
transform 1 0 111228 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1203
timestamp 1666464484
transform 1 0 111780 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1205
timestamp 1666464484
transform 1 0 111964 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1217
timestamp 1666464484
transform 1 0 113068 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1229
timestamp 1666464484
transform 1 0 114172 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1241
timestamp 1666464484
transform 1 0 115276 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1253
timestamp 1666464484
transform 1 0 116380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1259
timestamp 1666464484
transform 1 0 116932 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1261
timestamp 1666464484
transform 1 0 117116 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1273
timestamp 1666464484
transform 1 0 118220 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1285
timestamp 1666464484
transform 1 0 119324 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1297
timestamp 1666464484
transform 1 0 120428 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1309
timestamp 1666464484
transform 1 0 121532 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1315
timestamp 1666464484
transform 1 0 122084 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1317
timestamp 1666464484
transform 1 0 122268 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1329
timestamp 1666464484
transform 1 0 123372 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1341
timestamp 1666464484
transform 1 0 124476 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1353
timestamp 1666464484
transform 1 0 125580 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1365
timestamp 1666464484
transform 1 0 126684 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1371
timestamp 1666464484
transform 1 0 127236 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1373
timestamp 1666464484
transform 1 0 127420 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1385
timestamp 1666464484
transform 1 0 128524 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1397
timestamp 1666464484
transform 1 0 129628 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1409
timestamp 1666464484
transform 1 0 130732 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1421
timestamp 1666464484
transform 1 0 131836 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1427
timestamp 1666464484
transform 1 0 132388 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1429
timestamp 1666464484
transform 1 0 132572 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1441
timestamp 1666464484
transform 1 0 133676 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1453
timestamp 1666464484
transform 1 0 134780 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1465
timestamp 1666464484
transform 1 0 135884 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1477
timestamp 1666464484
transform 1 0 136988 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1483
timestamp 1666464484
transform 1 0 137540 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1485
timestamp 1666464484
transform 1 0 137724 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1497
timestamp 1666464484
transform 1 0 138828 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1509
timestamp 1666464484
transform 1 0 139932 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1521
timestamp 1666464484
transform 1 0 141036 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1533
timestamp 1666464484
transform 1 0 142140 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1539
timestamp 1666464484
transform 1 0 142692 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1541
timestamp 1666464484
transform 1 0 142876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1553
timestamp 1666464484
transform 1 0 143980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1565
timestamp 1666464484
transform 1 0 145084 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1577
timestamp 1666464484
transform 1 0 146188 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1589
timestamp 1666464484
transform 1 0 147292 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1595
timestamp 1666464484
transform 1 0 147844 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1597
timestamp 1666464484
transform 1 0 148028 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1666464484
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1666464484
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1666464484
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1666464484
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1666464484
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1666464484
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1666464484
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1666464484
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1666464484
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1666464484
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1666464484
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1666464484
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1666464484
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1666464484
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1666464484
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1666464484
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1666464484
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1666464484
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1666464484
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1666464484
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1666464484
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1666464484
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1666464484
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1666464484
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1666464484
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1666464484
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1666464484
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1666464484
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1666464484
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1666464484
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1666464484
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1666464484
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1666464484
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1666464484
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1666464484
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1666464484
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1666464484
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1666464484
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1666464484
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1666464484
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1666464484
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1666464484
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1666464484
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1666464484
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1666464484
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1666464484
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1666464484
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1666464484
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1666464484
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1666464484
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1666464484
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1666464484
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1666464484
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1666464484
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1666464484
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1666464484
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1666464484
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1666464484
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1666464484
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1666464484
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1666464484
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1666464484
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_585
timestamp 1666464484
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_597
timestamp 1666464484
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1666464484
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1666464484
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_617
timestamp 1666464484
transform 1 0 57868 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_629
timestamp 1666464484
transform 1 0 58972 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_641
timestamp 1666464484
transform 1 0 60076 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_653
timestamp 1666464484
transform 1 0 61180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_665
timestamp 1666464484
transform 1 0 62284 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_671
timestamp 1666464484
transform 1 0 62836 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_673
timestamp 1666464484
transform 1 0 63020 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_685
timestamp 1666464484
transform 1 0 64124 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_697
timestamp 1666464484
transform 1 0 65228 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_709
timestamp 1666464484
transform 1 0 66332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_721
timestamp 1666464484
transform 1 0 67436 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_727
timestamp 1666464484
transform 1 0 67988 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_729
timestamp 1666464484
transform 1 0 68172 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_741
timestamp 1666464484
transform 1 0 69276 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_753
timestamp 1666464484
transform 1 0 70380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_765
timestamp 1666464484
transform 1 0 71484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_777
timestamp 1666464484
transform 1 0 72588 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_783
timestamp 1666464484
transform 1 0 73140 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_785
timestamp 1666464484
transform 1 0 73324 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_797
timestamp 1666464484
transform 1 0 74428 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_809
timestamp 1666464484
transform 1 0 75532 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_821
timestamp 1666464484
transform 1 0 76636 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_833
timestamp 1666464484
transform 1 0 77740 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_839
timestamp 1666464484
transform 1 0 78292 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_841
timestamp 1666464484
transform 1 0 78476 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_853
timestamp 1666464484
transform 1 0 79580 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_865
timestamp 1666464484
transform 1 0 80684 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_877
timestamp 1666464484
transform 1 0 81788 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_889
timestamp 1666464484
transform 1 0 82892 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_895
timestamp 1666464484
transform 1 0 83444 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_897
timestamp 1666464484
transform 1 0 83628 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_909
timestamp 1666464484
transform 1 0 84732 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_921
timestamp 1666464484
transform 1 0 85836 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_933
timestamp 1666464484
transform 1 0 86940 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_945
timestamp 1666464484
transform 1 0 88044 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_951
timestamp 1666464484
transform 1 0 88596 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_953
timestamp 1666464484
transform 1 0 88780 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_965
timestamp 1666464484
transform 1 0 89884 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_977
timestamp 1666464484
transform 1 0 90988 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_989
timestamp 1666464484
transform 1 0 92092 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1001
timestamp 1666464484
transform 1 0 93196 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1007
timestamp 1666464484
transform 1 0 93748 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1009
timestamp 1666464484
transform 1 0 93932 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1021
timestamp 1666464484
transform 1 0 95036 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1033
timestamp 1666464484
transform 1 0 96140 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1045
timestamp 1666464484
transform 1 0 97244 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1057
timestamp 1666464484
transform 1 0 98348 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1063
timestamp 1666464484
transform 1 0 98900 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1065
timestamp 1666464484
transform 1 0 99084 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1077
timestamp 1666464484
transform 1 0 100188 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1089
timestamp 1666464484
transform 1 0 101292 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1101
timestamp 1666464484
transform 1 0 102396 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1113
timestamp 1666464484
transform 1 0 103500 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1119
timestamp 1666464484
transform 1 0 104052 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1121
timestamp 1666464484
transform 1 0 104236 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1133
timestamp 1666464484
transform 1 0 105340 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1145
timestamp 1666464484
transform 1 0 106444 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1157
timestamp 1666464484
transform 1 0 107548 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1169
timestamp 1666464484
transform 1 0 108652 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1175
timestamp 1666464484
transform 1 0 109204 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1177
timestamp 1666464484
transform 1 0 109388 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1189
timestamp 1666464484
transform 1 0 110492 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1201
timestamp 1666464484
transform 1 0 111596 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1213
timestamp 1666464484
transform 1 0 112700 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1225
timestamp 1666464484
transform 1 0 113804 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1231
timestamp 1666464484
transform 1 0 114356 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1233
timestamp 1666464484
transform 1 0 114540 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1245
timestamp 1666464484
transform 1 0 115644 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1257
timestamp 1666464484
transform 1 0 116748 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1269
timestamp 1666464484
transform 1 0 117852 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1281
timestamp 1666464484
transform 1 0 118956 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1287
timestamp 1666464484
transform 1 0 119508 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1289
timestamp 1666464484
transform 1 0 119692 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1301
timestamp 1666464484
transform 1 0 120796 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1313
timestamp 1666464484
transform 1 0 121900 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1325
timestamp 1666464484
transform 1 0 123004 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1337
timestamp 1666464484
transform 1 0 124108 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1343
timestamp 1666464484
transform 1 0 124660 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1345
timestamp 1666464484
transform 1 0 124844 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1357
timestamp 1666464484
transform 1 0 125948 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1369
timestamp 1666464484
transform 1 0 127052 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1381
timestamp 1666464484
transform 1 0 128156 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1393
timestamp 1666464484
transform 1 0 129260 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1399
timestamp 1666464484
transform 1 0 129812 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1401
timestamp 1666464484
transform 1 0 129996 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1413
timestamp 1666464484
transform 1 0 131100 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1425
timestamp 1666464484
transform 1 0 132204 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1437
timestamp 1666464484
transform 1 0 133308 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1449
timestamp 1666464484
transform 1 0 134412 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1455
timestamp 1666464484
transform 1 0 134964 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1457
timestamp 1666464484
transform 1 0 135148 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1469
timestamp 1666464484
transform 1 0 136252 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1481
timestamp 1666464484
transform 1 0 137356 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1493
timestamp 1666464484
transform 1 0 138460 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1505
timestamp 1666464484
transform 1 0 139564 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1511
timestamp 1666464484
transform 1 0 140116 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1513
timestamp 1666464484
transform 1 0 140300 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1525
timestamp 1666464484
transform 1 0 141404 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1537
timestamp 1666464484
transform 1 0 142508 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1549
timestamp 1666464484
transform 1 0 143612 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1561
timestamp 1666464484
transform 1 0 144716 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1567
timestamp 1666464484
transform 1 0 145268 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1569
timestamp 1666464484
transform 1 0 145452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1581
timestamp 1666464484
transform 1 0 146556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_1593
timestamp 1666464484
transform 1 0 147660 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_1601
timestamp 1666464484
transform 1 0 148396 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1666464484
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1666464484
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1666464484
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1666464484
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1666464484
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1666464484
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1666464484
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1666464484
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1666464484
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1666464484
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1666464484
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1666464484
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1666464484
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1666464484
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1666464484
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1666464484
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1666464484
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1666464484
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1666464484
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1666464484
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1666464484
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1666464484
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1666464484
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1666464484
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1666464484
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1666464484
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1666464484
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1666464484
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1666464484
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1666464484
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1666464484
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1666464484
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1666464484
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1666464484
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1666464484
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1666464484
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1666464484
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1666464484
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1666464484
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1666464484
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1666464484
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1666464484
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1666464484
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1666464484
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1666464484
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1666464484
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1666464484
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1666464484
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1666464484
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1666464484
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1666464484
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1666464484
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1666464484
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1666464484
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1666464484
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1666464484
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1666464484
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1666464484
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1666464484
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1666464484
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_569
timestamp 1666464484
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1666464484
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1666464484
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1666464484
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_601
timestamp 1666464484
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_613
timestamp 1666464484
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_625
timestamp 1666464484
transform 1 0 58604 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_637
timestamp 1666464484
transform 1 0 59708 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_643
timestamp 1666464484
transform 1 0 60260 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_645
timestamp 1666464484
transform 1 0 60444 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_657
timestamp 1666464484
transform 1 0 61548 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_669
timestamp 1666464484
transform 1 0 62652 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_681
timestamp 1666464484
transform 1 0 63756 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_693
timestamp 1666464484
transform 1 0 64860 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_699
timestamp 1666464484
transform 1 0 65412 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_701
timestamp 1666464484
transform 1 0 65596 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_713
timestamp 1666464484
transform 1 0 66700 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_725
timestamp 1666464484
transform 1 0 67804 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_737
timestamp 1666464484
transform 1 0 68908 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_749
timestamp 1666464484
transform 1 0 70012 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_755
timestamp 1666464484
transform 1 0 70564 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_757
timestamp 1666464484
transform 1 0 70748 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_769
timestamp 1666464484
transform 1 0 71852 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_781
timestamp 1666464484
transform 1 0 72956 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_793
timestamp 1666464484
transform 1 0 74060 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_805
timestamp 1666464484
transform 1 0 75164 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_811
timestamp 1666464484
transform 1 0 75716 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_813
timestamp 1666464484
transform 1 0 75900 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_825
timestamp 1666464484
transform 1 0 77004 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_837
timestamp 1666464484
transform 1 0 78108 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_849
timestamp 1666464484
transform 1 0 79212 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_861
timestamp 1666464484
transform 1 0 80316 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_867
timestamp 1666464484
transform 1 0 80868 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_869
timestamp 1666464484
transform 1 0 81052 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_881
timestamp 1666464484
transform 1 0 82156 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_893
timestamp 1666464484
transform 1 0 83260 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_905
timestamp 1666464484
transform 1 0 84364 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_917
timestamp 1666464484
transform 1 0 85468 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_923
timestamp 1666464484
transform 1 0 86020 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_925
timestamp 1666464484
transform 1 0 86204 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_937
timestamp 1666464484
transform 1 0 87308 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_949
timestamp 1666464484
transform 1 0 88412 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_961
timestamp 1666464484
transform 1 0 89516 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_973
timestamp 1666464484
transform 1 0 90620 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_979
timestamp 1666464484
transform 1 0 91172 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_981
timestamp 1666464484
transform 1 0 91356 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_993
timestamp 1666464484
transform 1 0 92460 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1005
timestamp 1666464484
transform 1 0 93564 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1017
timestamp 1666464484
transform 1 0 94668 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1029
timestamp 1666464484
transform 1 0 95772 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1035
timestamp 1666464484
transform 1 0 96324 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1037
timestamp 1666464484
transform 1 0 96508 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1049
timestamp 1666464484
transform 1 0 97612 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1061
timestamp 1666464484
transform 1 0 98716 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1073
timestamp 1666464484
transform 1 0 99820 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1085
timestamp 1666464484
transform 1 0 100924 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1091
timestamp 1666464484
transform 1 0 101476 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1093
timestamp 1666464484
transform 1 0 101660 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1105
timestamp 1666464484
transform 1 0 102764 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1117
timestamp 1666464484
transform 1 0 103868 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1129
timestamp 1666464484
transform 1 0 104972 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1141
timestamp 1666464484
transform 1 0 106076 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1147
timestamp 1666464484
transform 1 0 106628 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1149
timestamp 1666464484
transform 1 0 106812 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1161
timestamp 1666464484
transform 1 0 107916 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1173
timestamp 1666464484
transform 1 0 109020 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1185
timestamp 1666464484
transform 1 0 110124 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1197
timestamp 1666464484
transform 1 0 111228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1203
timestamp 1666464484
transform 1 0 111780 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1205
timestamp 1666464484
transform 1 0 111964 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1217
timestamp 1666464484
transform 1 0 113068 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1229
timestamp 1666464484
transform 1 0 114172 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1241
timestamp 1666464484
transform 1 0 115276 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1253
timestamp 1666464484
transform 1 0 116380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1259
timestamp 1666464484
transform 1 0 116932 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1261
timestamp 1666464484
transform 1 0 117116 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1273
timestamp 1666464484
transform 1 0 118220 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1285
timestamp 1666464484
transform 1 0 119324 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1297
timestamp 1666464484
transform 1 0 120428 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1309
timestamp 1666464484
transform 1 0 121532 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1315
timestamp 1666464484
transform 1 0 122084 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1317
timestamp 1666464484
transform 1 0 122268 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1329
timestamp 1666464484
transform 1 0 123372 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1341
timestamp 1666464484
transform 1 0 124476 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1353
timestamp 1666464484
transform 1 0 125580 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1365
timestamp 1666464484
transform 1 0 126684 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1371
timestamp 1666464484
transform 1 0 127236 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1373
timestamp 1666464484
transform 1 0 127420 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1385
timestamp 1666464484
transform 1 0 128524 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1397
timestamp 1666464484
transform 1 0 129628 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1409
timestamp 1666464484
transform 1 0 130732 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1421
timestamp 1666464484
transform 1 0 131836 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1427
timestamp 1666464484
transform 1 0 132388 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1429
timestamp 1666464484
transform 1 0 132572 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1441
timestamp 1666464484
transform 1 0 133676 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1453
timestamp 1666464484
transform 1 0 134780 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1465
timestamp 1666464484
transform 1 0 135884 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1477
timestamp 1666464484
transform 1 0 136988 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1483
timestamp 1666464484
transform 1 0 137540 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1485
timestamp 1666464484
transform 1 0 137724 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1497
timestamp 1666464484
transform 1 0 138828 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1509
timestamp 1666464484
transform 1 0 139932 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1521
timestamp 1666464484
transform 1 0 141036 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1533
timestamp 1666464484
transform 1 0 142140 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1539
timestamp 1666464484
transform 1 0 142692 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1541
timestamp 1666464484
transform 1 0 142876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1553
timestamp 1666464484
transform 1 0 143980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1565
timestamp 1666464484
transform 1 0 145084 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1577
timestamp 1666464484
transform 1 0 146188 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1589
timestamp 1666464484
transform 1 0 147292 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1595
timestamp 1666464484
transform 1 0 147844 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1597
timestamp 1666464484
transform 1 0 148028 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1666464484
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1666464484
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1666464484
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1666464484
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1666464484
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1666464484
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1666464484
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1666464484
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1666464484
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1666464484
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1666464484
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1666464484
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1666464484
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1666464484
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1666464484
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1666464484
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1666464484
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1666464484
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1666464484
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1666464484
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1666464484
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1666464484
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1666464484
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1666464484
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1666464484
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1666464484
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1666464484
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1666464484
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1666464484
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1666464484
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1666464484
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1666464484
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1666464484
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1666464484
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1666464484
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1666464484
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1666464484
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1666464484
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1666464484
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1666464484
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1666464484
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1666464484
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1666464484
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1666464484
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1666464484
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1666464484
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1666464484
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1666464484
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1666464484
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1666464484
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1666464484
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1666464484
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1666464484
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1666464484
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1666464484
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1666464484
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1666464484
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1666464484
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1666464484
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1666464484
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_561
timestamp 1666464484
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_573
timestamp 1666464484
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_585
timestamp 1666464484
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_597
timestamp 1666464484
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1666464484
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1666464484
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_617
timestamp 1666464484
transform 1 0 57868 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_629
timestamp 1666464484
transform 1 0 58972 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_641
timestamp 1666464484
transform 1 0 60076 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_653
timestamp 1666464484
transform 1 0 61180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_665
timestamp 1666464484
transform 1 0 62284 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_671
timestamp 1666464484
transform 1 0 62836 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_673
timestamp 1666464484
transform 1 0 63020 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_685
timestamp 1666464484
transform 1 0 64124 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_697
timestamp 1666464484
transform 1 0 65228 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_709
timestamp 1666464484
transform 1 0 66332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_721
timestamp 1666464484
transform 1 0 67436 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_727
timestamp 1666464484
transform 1 0 67988 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_729
timestamp 1666464484
transform 1 0 68172 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_741
timestamp 1666464484
transform 1 0 69276 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_753
timestamp 1666464484
transform 1 0 70380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_765
timestamp 1666464484
transform 1 0 71484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_777
timestamp 1666464484
transform 1 0 72588 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_783
timestamp 1666464484
transform 1 0 73140 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_785
timestamp 1666464484
transform 1 0 73324 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_797
timestamp 1666464484
transform 1 0 74428 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_809
timestamp 1666464484
transform 1 0 75532 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_821
timestamp 1666464484
transform 1 0 76636 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_833
timestamp 1666464484
transform 1 0 77740 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_839
timestamp 1666464484
transform 1 0 78292 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_841
timestamp 1666464484
transform 1 0 78476 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_853
timestamp 1666464484
transform 1 0 79580 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_865
timestamp 1666464484
transform 1 0 80684 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_877
timestamp 1666464484
transform 1 0 81788 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_889
timestamp 1666464484
transform 1 0 82892 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_895
timestamp 1666464484
transform 1 0 83444 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_897
timestamp 1666464484
transform 1 0 83628 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_909
timestamp 1666464484
transform 1 0 84732 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_921
timestamp 1666464484
transform 1 0 85836 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_933
timestamp 1666464484
transform 1 0 86940 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_945
timestamp 1666464484
transform 1 0 88044 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_951
timestamp 1666464484
transform 1 0 88596 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_953
timestamp 1666464484
transform 1 0 88780 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_965
timestamp 1666464484
transform 1 0 89884 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_977
timestamp 1666464484
transform 1 0 90988 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_989
timestamp 1666464484
transform 1 0 92092 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1001
timestamp 1666464484
transform 1 0 93196 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1007
timestamp 1666464484
transform 1 0 93748 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1009
timestamp 1666464484
transform 1 0 93932 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1021
timestamp 1666464484
transform 1 0 95036 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1033
timestamp 1666464484
transform 1 0 96140 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1045
timestamp 1666464484
transform 1 0 97244 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1057
timestamp 1666464484
transform 1 0 98348 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1063
timestamp 1666464484
transform 1 0 98900 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1065
timestamp 1666464484
transform 1 0 99084 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1077
timestamp 1666464484
transform 1 0 100188 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1089
timestamp 1666464484
transform 1 0 101292 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1101
timestamp 1666464484
transform 1 0 102396 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1113
timestamp 1666464484
transform 1 0 103500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1119
timestamp 1666464484
transform 1 0 104052 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1121
timestamp 1666464484
transform 1 0 104236 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1133
timestamp 1666464484
transform 1 0 105340 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1145
timestamp 1666464484
transform 1 0 106444 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1157
timestamp 1666464484
transform 1 0 107548 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1169
timestamp 1666464484
transform 1 0 108652 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1175
timestamp 1666464484
transform 1 0 109204 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1177
timestamp 1666464484
transform 1 0 109388 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1189
timestamp 1666464484
transform 1 0 110492 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1201
timestamp 1666464484
transform 1 0 111596 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1213
timestamp 1666464484
transform 1 0 112700 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1225
timestamp 1666464484
transform 1 0 113804 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1231
timestamp 1666464484
transform 1 0 114356 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1233
timestamp 1666464484
transform 1 0 114540 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1245
timestamp 1666464484
transform 1 0 115644 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1257
timestamp 1666464484
transform 1 0 116748 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1269
timestamp 1666464484
transform 1 0 117852 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1281
timestamp 1666464484
transform 1 0 118956 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1287
timestamp 1666464484
transform 1 0 119508 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1289
timestamp 1666464484
transform 1 0 119692 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1301
timestamp 1666464484
transform 1 0 120796 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1313
timestamp 1666464484
transform 1 0 121900 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1325
timestamp 1666464484
transform 1 0 123004 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1337
timestamp 1666464484
transform 1 0 124108 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1343
timestamp 1666464484
transform 1 0 124660 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1345
timestamp 1666464484
transform 1 0 124844 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1357
timestamp 1666464484
transform 1 0 125948 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1369
timestamp 1666464484
transform 1 0 127052 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1381
timestamp 1666464484
transform 1 0 128156 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1393
timestamp 1666464484
transform 1 0 129260 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1399
timestamp 1666464484
transform 1 0 129812 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1401
timestamp 1666464484
transform 1 0 129996 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1413
timestamp 1666464484
transform 1 0 131100 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1425
timestamp 1666464484
transform 1 0 132204 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1437
timestamp 1666464484
transform 1 0 133308 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1449
timestamp 1666464484
transform 1 0 134412 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1455
timestamp 1666464484
transform 1 0 134964 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1457
timestamp 1666464484
transform 1 0 135148 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1469
timestamp 1666464484
transform 1 0 136252 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1481
timestamp 1666464484
transform 1 0 137356 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1493
timestamp 1666464484
transform 1 0 138460 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1505
timestamp 1666464484
transform 1 0 139564 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1511
timestamp 1666464484
transform 1 0 140116 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1513
timestamp 1666464484
transform 1 0 140300 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1525
timestamp 1666464484
transform 1 0 141404 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1537
timestamp 1666464484
transform 1 0 142508 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1549
timestamp 1666464484
transform 1 0 143612 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1561
timestamp 1666464484
transform 1 0 144716 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1567
timestamp 1666464484
transform 1 0 145268 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1569
timestamp 1666464484
transform 1 0 145452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1581
timestamp 1666464484
transform 1 0 146556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_1593
timestamp 1666464484
transform 1 0 147660 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_1601
timestamp 1666464484
transform 1 0 148396 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1666464484
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1666464484
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1666464484
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1666464484
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1666464484
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1666464484
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1666464484
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1666464484
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1666464484
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1666464484
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1666464484
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1666464484
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1666464484
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1666464484
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1666464484
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1666464484
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1666464484
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1666464484
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1666464484
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1666464484
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1666464484
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1666464484
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1666464484
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1666464484
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1666464484
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1666464484
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1666464484
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1666464484
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1666464484
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1666464484
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1666464484
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1666464484
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1666464484
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1666464484
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1666464484
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1666464484
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1666464484
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1666464484
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1666464484
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1666464484
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1666464484
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1666464484
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1666464484
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1666464484
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1666464484
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1666464484
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1666464484
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1666464484
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1666464484
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1666464484
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1666464484
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1666464484
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1666464484
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1666464484
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1666464484
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1666464484
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1666464484
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1666464484
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1666464484
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1666464484
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_569
timestamp 1666464484
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1666464484
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1666464484
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_589
timestamp 1666464484
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_601
timestamp 1666464484
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_613
timestamp 1666464484
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_625
timestamp 1666464484
transform 1 0 58604 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_637
timestamp 1666464484
transform 1 0 59708 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_643
timestamp 1666464484
transform 1 0 60260 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_645
timestamp 1666464484
transform 1 0 60444 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_657
timestamp 1666464484
transform 1 0 61548 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_669
timestamp 1666464484
transform 1 0 62652 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_681
timestamp 1666464484
transform 1 0 63756 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_693
timestamp 1666464484
transform 1 0 64860 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_699
timestamp 1666464484
transform 1 0 65412 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_701
timestamp 1666464484
transform 1 0 65596 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_713
timestamp 1666464484
transform 1 0 66700 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_725
timestamp 1666464484
transform 1 0 67804 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_737
timestamp 1666464484
transform 1 0 68908 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_749
timestamp 1666464484
transform 1 0 70012 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_755
timestamp 1666464484
transform 1 0 70564 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_757
timestamp 1666464484
transform 1 0 70748 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_769
timestamp 1666464484
transform 1 0 71852 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_781
timestamp 1666464484
transform 1 0 72956 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_793
timestamp 1666464484
transform 1 0 74060 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_805
timestamp 1666464484
transform 1 0 75164 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_811
timestamp 1666464484
transform 1 0 75716 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_813
timestamp 1666464484
transform 1 0 75900 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_825
timestamp 1666464484
transform 1 0 77004 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_837
timestamp 1666464484
transform 1 0 78108 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_849
timestamp 1666464484
transform 1 0 79212 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_861
timestamp 1666464484
transform 1 0 80316 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_867
timestamp 1666464484
transform 1 0 80868 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_869
timestamp 1666464484
transform 1 0 81052 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_881
timestamp 1666464484
transform 1 0 82156 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_893
timestamp 1666464484
transform 1 0 83260 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_905
timestamp 1666464484
transform 1 0 84364 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_917
timestamp 1666464484
transform 1 0 85468 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_923
timestamp 1666464484
transform 1 0 86020 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_925
timestamp 1666464484
transform 1 0 86204 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_937
timestamp 1666464484
transform 1 0 87308 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_949
timestamp 1666464484
transform 1 0 88412 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_961
timestamp 1666464484
transform 1 0 89516 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_973
timestamp 1666464484
transform 1 0 90620 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_979
timestamp 1666464484
transform 1 0 91172 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_981
timestamp 1666464484
transform 1 0 91356 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_993
timestamp 1666464484
transform 1 0 92460 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1005
timestamp 1666464484
transform 1 0 93564 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1017
timestamp 1666464484
transform 1 0 94668 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1029
timestamp 1666464484
transform 1 0 95772 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1035
timestamp 1666464484
transform 1 0 96324 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1037
timestamp 1666464484
transform 1 0 96508 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1049
timestamp 1666464484
transform 1 0 97612 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1061
timestamp 1666464484
transform 1 0 98716 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1073
timestamp 1666464484
transform 1 0 99820 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1085
timestamp 1666464484
transform 1 0 100924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1091
timestamp 1666464484
transform 1 0 101476 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1093
timestamp 1666464484
transform 1 0 101660 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1105
timestamp 1666464484
transform 1 0 102764 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1117
timestamp 1666464484
transform 1 0 103868 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1129
timestamp 1666464484
transform 1 0 104972 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1141
timestamp 1666464484
transform 1 0 106076 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1147
timestamp 1666464484
transform 1 0 106628 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1149
timestamp 1666464484
transform 1 0 106812 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1161
timestamp 1666464484
transform 1 0 107916 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1173
timestamp 1666464484
transform 1 0 109020 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1185
timestamp 1666464484
transform 1 0 110124 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1197
timestamp 1666464484
transform 1 0 111228 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1203
timestamp 1666464484
transform 1 0 111780 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1205
timestamp 1666464484
transform 1 0 111964 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1217
timestamp 1666464484
transform 1 0 113068 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1229
timestamp 1666464484
transform 1 0 114172 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1241
timestamp 1666464484
transform 1 0 115276 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1253
timestamp 1666464484
transform 1 0 116380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1259
timestamp 1666464484
transform 1 0 116932 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1261
timestamp 1666464484
transform 1 0 117116 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1273
timestamp 1666464484
transform 1 0 118220 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1285
timestamp 1666464484
transform 1 0 119324 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1297
timestamp 1666464484
transform 1 0 120428 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1309
timestamp 1666464484
transform 1 0 121532 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1315
timestamp 1666464484
transform 1 0 122084 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1317
timestamp 1666464484
transform 1 0 122268 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1329
timestamp 1666464484
transform 1 0 123372 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1341
timestamp 1666464484
transform 1 0 124476 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1353
timestamp 1666464484
transform 1 0 125580 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1365
timestamp 1666464484
transform 1 0 126684 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1371
timestamp 1666464484
transform 1 0 127236 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1373
timestamp 1666464484
transform 1 0 127420 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1385
timestamp 1666464484
transform 1 0 128524 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1397
timestamp 1666464484
transform 1 0 129628 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1409
timestamp 1666464484
transform 1 0 130732 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1421
timestamp 1666464484
transform 1 0 131836 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1427
timestamp 1666464484
transform 1 0 132388 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1429
timestamp 1666464484
transform 1 0 132572 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1441
timestamp 1666464484
transform 1 0 133676 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1453
timestamp 1666464484
transform 1 0 134780 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1465
timestamp 1666464484
transform 1 0 135884 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1477
timestamp 1666464484
transform 1 0 136988 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1483
timestamp 1666464484
transform 1 0 137540 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1485
timestamp 1666464484
transform 1 0 137724 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1497
timestamp 1666464484
transform 1 0 138828 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1509
timestamp 1666464484
transform 1 0 139932 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1521
timestamp 1666464484
transform 1 0 141036 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1533
timestamp 1666464484
transform 1 0 142140 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1539
timestamp 1666464484
transform 1 0 142692 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1541
timestamp 1666464484
transform 1 0 142876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1553
timestamp 1666464484
transform 1 0 143980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1565
timestamp 1666464484
transform 1 0 145084 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1577
timestamp 1666464484
transform 1 0 146188 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1589
timestamp 1666464484
transform 1 0 147292 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1595
timestamp 1666464484
transform 1 0 147844 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1597
timestamp 1666464484
transform 1 0 148028 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1666464484
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1666464484
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1666464484
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1666464484
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1666464484
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1666464484
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1666464484
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1666464484
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1666464484
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1666464484
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1666464484
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1666464484
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1666464484
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1666464484
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1666464484
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1666464484
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1666464484
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1666464484
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1666464484
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1666464484
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1666464484
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1666464484
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1666464484
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1666464484
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1666464484
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1666464484
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1666464484
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1666464484
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1666464484
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1666464484
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1666464484
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1666464484
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1666464484
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1666464484
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1666464484
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1666464484
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1666464484
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1666464484
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1666464484
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1666464484
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1666464484
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1666464484
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1666464484
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1666464484
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1666464484
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1666464484
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1666464484
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1666464484
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1666464484
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1666464484
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1666464484
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1666464484
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1666464484
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1666464484
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1666464484
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1666464484
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1666464484
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1666464484
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1666464484
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1666464484
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1666464484
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1666464484
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1666464484
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1666464484
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1666464484
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1666464484
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_617
timestamp 1666464484
transform 1 0 57868 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_629
timestamp 1666464484
transform 1 0 58972 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_641
timestamp 1666464484
transform 1 0 60076 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_653
timestamp 1666464484
transform 1 0 61180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_665
timestamp 1666464484
transform 1 0 62284 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_671
timestamp 1666464484
transform 1 0 62836 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_673
timestamp 1666464484
transform 1 0 63020 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_685
timestamp 1666464484
transform 1 0 64124 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_697
timestamp 1666464484
transform 1 0 65228 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_709
timestamp 1666464484
transform 1 0 66332 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_721
timestamp 1666464484
transform 1 0 67436 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_727
timestamp 1666464484
transform 1 0 67988 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_729
timestamp 1666464484
transform 1 0 68172 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_741
timestamp 1666464484
transform 1 0 69276 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_753
timestamp 1666464484
transform 1 0 70380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_765
timestamp 1666464484
transform 1 0 71484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_777
timestamp 1666464484
transform 1 0 72588 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_783
timestamp 1666464484
transform 1 0 73140 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_785
timestamp 1666464484
transform 1 0 73324 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_797
timestamp 1666464484
transform 1 0 74428 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_809
timestamp 1666464484
transform 1 0 75532 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_821
timestamp 1666464484
transform 1 0 76636 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_833
timestamp 1666464484
transform 1 0 77740 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_839
timestamp 1666464484
transform 1 0 78292 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_841
timestamp 1666464484
transform 1 0 78476 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_853
timestamp 1666464484
transform 1 0 79580 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_865
timestamp 1666464484
transform 1 0 80684 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_877
timestamp 1666464484
transform 1 0 81788 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_889
timestamp 1666464484
transform 1 0 82892 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_895
timestamp 1666464484
transform 1 0 83444 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_897
timestamp 1666464484
transform 1 0 83628 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_909
timestamp 1666464484
transform 1 0 84732 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_921
timestamp 1666464484
transform 1 0 85836 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_933
timestamp 1666464484
transform 1 0 86940 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_945
timestamp 1666464484
transform 1 0 88044 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_951
timestamp 1666464484
transform 1 0 88596 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_953
timestamp 1666464484
transform 1 0 88780 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_965
timestamp 1666464484
transform 1 0 89884 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_977
timestamp 1666464484
transform 1 0 90988 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_989
timestamp 1666464484
transform 1 0 92092 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1001
timestamp 1666464484
transform 1 0 93196 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1007
timestamp 1666464484
transform 1 0 93748 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1009
timestamp 1666464484
transform 1 0 93932 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1021
timestamp 1666464484
transform 1 0 95036 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1033
timestamp 1666464484
transform 1 0 96140 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1045
timestamp 1666464484
transform 1 0 97244 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1057
timestamp 1666464484
transform 1 0 98348 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1063
timestamp 1666464484
transform 1 0 98900 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1065
timestamp 1666464484
transform 1 0 99084 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1077
timestamp 1666464484
transform 1 0 100188 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1089
timestamp 1666464484
transform 1 0 101292 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1101
timestamp 1666464484
transform 1 0 102396 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1113
timestamp 1666464484
transform 1 0 103500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1119
timestamp 1666464484
transform 1 0 104052 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1121
timestamp 1666464484
transform 1 0 104236 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1133
timestamp 1666464484
transform 1 0 105340 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1145
timestamp 1666464484
transform 1 0 106444 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1157
timestamp 1666464484
transform 1 0 107548 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1169
timestamp 1666464484
transform 1 0 108652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1175
timestamp 1666464484
transform 1 0 109204 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1177
timestamp 1666464484
transform 1 0 109388 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1189
timestamp 1666464484
transform 1 0 110492 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1201
timestamp 1666464484
transform 1 0 111596 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1213
timestamp 1666464484
transform 1 0 112700 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1225
timestamp 1666464484
transform 1 0 113804 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1231
timestamp 1666464484
transform 1 0 114356 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1233
timestamp 1666464484
transform 1 0 114540 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1245
timestamp 1666464484
transform 1 0 115644 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1257
timestamp 1666464484
transform 1 0 116748 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1269
timestamp 1666464484
transform 1 0 117852 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1281
timestamp 1666464484
transform 1 0 118956 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1287
timestamp 1666464484
transform 1 0 119508 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1289
timestamp 1666464484
transform 1 0 119692 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1301
timestamp 1666464484
transform 1 0 120796 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1313
timestamp 1666464484
transform 1 0 121900 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1325
timestamp 1666464484
transform 1 0 123004 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1337
timestamp 1666464484
transform 1 0 124108 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1343
timestamp 1666464484
transform 1 0 124660 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1345
timestamp 1666464484
transform 1 0 124844 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1357
timestamp 1666464484
transform 1 0 125948 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1369
timestamp 1666464484
transform 1 0 127052 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1381
timestamp 1666464484
transform 1 0 128156 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1393
timestamp 1666464484
transform 1 0 129260 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1399
timestamp 1666464484
transform 1 0 129812 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1401
timestamp 1666464484
transform 1 0 129996 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1413
timestamp 1666464484
transform 1 0 131100 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1425
timestamp 1666464484
transform 1 0 132204 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1437
timestamp 1666464484
transform 1 0 133308 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1449
timestamp 1666464484
transform 1 0 134412 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1455
timestamp 1666464484
transform 1 0 134964 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1457
timestamp 1666464484
transform 1 0 135148 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1469
timestamp 1666464484
transform 1 0 136252 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1481
timestamp 1666464484
transform 1 0 137356 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1493
timestamp 1666464484
transform 1 0 138460 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1505
timestamp 1666464484
transform 1 0 139564 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1511
timestamp 1666464484
transform 1 0 140116 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1513
timestamp 1666464484
transform 1 0 140300 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1525
timestamp 1666464484
transform 1 0 141404 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1537
timestamp 1666464484
transform 1 0 142508 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1549
timestamp 1666464484
transform 1 0 143612 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1561
timestamp 1666464484
transform 1 0 144716 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1567
timestamp 1666464484
transform 1 0 145268 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1569
timestamp 1666464484
transform 1 0 145452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1581
timestamp 1666464484
transform 1 0 146556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_1593
timestamp 1666464484
transform 1 0 147660 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_1601
timestamp 1666464484
transform 1 0 148396 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1666464484
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1666464484
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1666464484
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1666464484
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1666464484
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1666464484
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1666464484
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1666464484
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1666464484
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1666464484
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1666464484
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1666464484
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1666464484
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1666464484
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1666464484
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1666464484
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1666464484
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1666464484
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1666464484
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1666464484
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1666464484
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1666464484
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1666464484
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1666464484
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1666464484
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1666464484
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1666464484
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1666464484
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1666464484
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1666464484
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1666464484
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1666464484
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1666464484
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1666464484
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1666464484
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1666464484
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1666464484
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1666464484
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1666464484
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1666464484
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1666464484
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1666464484
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1666464484
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1666464484
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1666464484
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1666464484
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1666464484
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1666464484
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1666464484
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1666464484
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1666464484
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1666464484
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1666464484
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1666464484
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1666464484
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1666464484
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1666464484
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1666464484
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1666464484
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1666464484
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_569
timestamp 1666464484
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1666464484
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1666464484
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1666464484
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1666464484
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_613
timestamp 1666464484
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_625
timestamp 1666464484
transform 1 0 58604 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_637
timestamp 1666464484
transform 1 0 59708 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_643
timestamp 1666464484
transform 1 0 60260 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_645
timestamp 1666464484
transform 1 0 60444 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_657
timestamp 1666464484
transform 1 0 61548 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_669
timestamp 1666464484
transform 1 0 62652 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_681
timestamp 1666464484
transform 1 0 63756 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_693
timestamp 1666464484
transform 1 0 64860 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_699
timestamp 1666464484
transform 1 0 65412 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_701
timestamp 1666464484
transform 1 0 65596 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_713
timestamp 1666464484
transform 1 0 66700 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_725
timestamp 1666464484
transform 1 0 67804 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_737
timestamp 1666464484
transform 1 0 68908 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_749
timestamp 1666464484
transform 1 0 70012 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_755
timestamp 1666464484
transform 1 0 70564 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_757
timestamp 1666464484
transform 1 0 70748 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_769
timestamp 1666464484
transform 1 0 71852 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_781
timestamp 1666464484
transform 1 0 72956 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_793
timestamp 1666464484
transform 1 0 74060 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_805
timestamp 1666464484
transform 1 0 75164 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_811
timestamp 1666464484
transform 1 0 75716 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_813
timestamp 1666464484
transform 1 0 75900 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_825
timestamp 1666464484
transform 1 0 77004 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_837
timestamp 1666464484
transform 1 0 78108 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_849
timestamp 1666464484
transform 1 0 79212 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_861
timestamp 1666464484
transform 1 0 80316 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_867
timestamp 1666464484
transform 1 0 80868 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_869
timestamp 1666464484
transform 1 0 81052 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_881
timestamp 1666464484
transform 1 0 82156 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_893
timestamp 1666464484
transform 1 0 83260 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_905
timestamp 1666464484
transform 1 0 84364 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_917
timestamp 1666464484
transform 1 0 85468 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_923
timestamp 1666464484
transform 1 0 86020 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_925
timestamp 1666464484
transform 1 0 86204 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_937
timestamp 1666464484
transform 1 0 87308 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_949
timestamp 1666464484
transform 1 0 88412 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_961
timestamp 1666464484
transform 1 0 89516 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_973
timestamp 1666464484
transform 1 0 90620 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_979
timestamp 1666464484
transform 1 0 91172 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_981
timestamp 1666464484
transform 1 0 91356 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_993
timestamp 1666464484
transform 1 0 92460 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1005
timestamp 1666464484
transform 1 0 93564 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1017
timestamp 1666464484
transform 1 0 94668 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1029
timestamp 1666464484
transform 1 0 95772 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1035
timestamp 1666464484
transform 1 0 96324 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1037
timestamp 1666464484
transform 1 0 96508 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1049
timestamp 1666464484
transform 1 0 97612 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1061
timestamp 1666464484
transform 1 0 98716 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1073
timestamp 1666464484
transform 1 0 99820 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1085
timestamp 1666464484
transform 1 0 100924 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1091
timestamp 1666464484
transform 1 0 101476 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1093
timestamp 1666464484
transform 1 0 101660 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1105
timestamp 1666464484
transform 1 0 102764 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1117
timestamp 1666464484
transform 1 0 103868 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1129
timestamp 1666464484
transform 1 0 104972 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1141
timestamp 1666464484
transform 1 0 106076 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1147
timestamp 1666464484
transform 1 0 106628 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1149
timestamp 1666464484
transform 1 0 106812 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1161
timestamp 1666464484
transform 1 0 107916 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1173
timestamp 1666464484
transform 1 0 109020 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1185
timestamp 1666464484
transform 1 0 110124 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1197
timestamp 1666464484
transform 1 0 111228 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1203
timestamp 1666464484
transform 1 0 111780 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1205
timestamp 1666464484
transform 1 0 111964 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1217
timestamp 1666464484
transform 1 0 113068 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1229
timestamp 1666464484
transform 1 0 114172 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1241
timestamp 1666464484
transform 1 0 115276 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1253
timestamp 1666464484
transform 1 0 116380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1259
timestamp 1666464484
transform 1 0 116932 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1261
timestamp 1666464484
transform 1 0 117116 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1273
timestamp 1666464484
transform 1 0 118220 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1285
timestamp 1666464484
transform 1 0 119324 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1297
timestamp 1666464484
transform 1 0 120428 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1309
timestamp 1666464484
transform 1 0 121532 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1315
timestamp 1666464484
transform 1 0 122084 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1317
timestamp 1666464484
transform 1 0 122268 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1329
timestamp 1666464484
transform 1 0 123372 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1341
timestamp 1666464484
transform 1 0 124476 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1353
timestamp 1666464484
transform 1 0 125580 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1365
timestamp 1666464484
transform 1 0 126684 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1371
timestamp 1666464484
transform 1 0 127236 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1373
timestamp 1666464484
transform 1 0 127420 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1385
timestamp 1666464484
transform 1 0 128524 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1397
timestamp 1666464484
transform 1 0 129628 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1409
timestamp 1666464484
transform 1 0 130732 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1421
timestamp 1666464484
transform 1 0 131836 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1427
timestamp 1666464484
transform 1 0 132388 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1429
timestamp 1666464484
transform 1 0 132572 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1441
timestamp 1666464484
transform 1 0 133676 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1453
timestamp 1666464484
transform 1 0 134780 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1465
timestamp 1666464484
transform 1 0 135884 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1477
timestamp 1666464484
transform 1 0 136988 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1483
timestamp 1666464484
transform 1 0 137540 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1485
timestamp 1666464484
transform 1 0 137724 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1497
timestamp 1666464484
transform 1 0 138828 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1509
timestamp 1666464484
transform 1 0 139932 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1521
timestamp 1666464484
transform 1 0 141036 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1533
timestamp 1666464484
transform 1 0 142140 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1539
timestamp 1666464484
transform 1 0 142692 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1541
timestamp 1666464484
transform 1 0 142876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1553
timestamp 1666464484
transform 1 0 143980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1565
timestamp 1666464484
transform 1 0 145084 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1577
timestamp 1666464484
transform 1 0 146188 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1589
timestamp 1666464484
transform 1 0 147292 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1595
timestamp 1666464484
transform 1 0 147844 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1597
timestamp 1666464484
transform 1 0 148028 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1666464484
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1666464484
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1666464484
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1666464484
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1666464484
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1666464484
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1666464484
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1666464484
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1666464484
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1666464484
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1666464484
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1666464484
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1666464484
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1666464484
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1666464484
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1666464484
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1666464484
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1666464484
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1666464484
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1666464484
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1666464484
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1666464484
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1666464484
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1666464484
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1666464484
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1666464484
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1666464484
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1666464484
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1666464484
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1666464484
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1666464484
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1666464484
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1666464484
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1666464484
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1666464484
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1666464484
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1666464484
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1666464484
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1666464484
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1666464484
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1666464484
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1666464484
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1666464484
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1666464484
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1666464484
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1666464484
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1666464484
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1666464484
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1666464484
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1666464484
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1666464484
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1666464484
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1666464484
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1666464484
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1666464484
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1666464484
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1666464484
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1666464484
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1666464484
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1666464484
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1666464484
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1666464484
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1666464484
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1666464484
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1666464484
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1666464484
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_617
timestamp 1666464484
transform 1 0 57868 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_629
timestamp 1666464484
transform 1 0 58972 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_641
timestamp 1666464484
transform 1 0 60076 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_653
timestamp 1666464484
transform 1 0 61180 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_665
timestamp 1666464484
transform 1 0 62284 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_671
timestamp 1666464484
transform 1 0 62836 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_673
timestamp 1666464484
transform 1 0 63020 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_685
timestamp 1666464484
transform 1 0 64124 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_697
timestamp 1666464484
transform 1 0 65228 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_709
timestamp 1666464484
transform 1 0 66332 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_721
timestamp 1666464484
transform 1 0 67436 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_727
timestamp 1666464484
transform 1 0 67988 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_729
timestamp 1666464484
transform 1 0 68172 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_741
timestamp 1666464484
transform 1 0 69276 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_753
timestamp 1666464484
transform 1 0 70380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_765
timestamp 1666464484
transform 1 0 71484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_777
timestamp 1666464484
transform 1 0 72588 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_783
timestamp 1666464484
transform 1 0 73140 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_785
timestamp 1666464484
transform 1 0 73324 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_797
timestamp 1666464484
transform 1 0 74428 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_809
timestamp 1666464484
transform 1 0 75532 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_821
timestamp 1666464484
transform 1 0 76636 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_833
timestamp 1666464484
transform 1 0 77740 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_839
timestamp 1666464484
transform 1 0 78292 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_841
timestamp 1666464484
transform 1 0 78476 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_853
timestamp 1666464484
transform 1 0 79580 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_865
timestamp 1666464484
transform 1 0 80684 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_877
timestamp 1666464484
transform 1 0 81788 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_889
timestamp 1666464484
transform 1 0 82892 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_895
timestamp 1666464484
transform 1 0 83444 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_897
timestamp 1666464484
transform 1 0 83628 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_909
timestamp 1666464484
transform 1 0 84732 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_921
timestamp 1666464484
transform 1 0 85836 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_933
timestamp 1666464484
transform 1 0 86940 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_945
timestamp 1666464484
transform 1 0 88044 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_951
timestamp 1666464484
transform 1 0 88596 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_953
timestamp 1666464484
transform 1 0 88780 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_965
timestamp 1666464484
transform 1 0 89884 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_977
timestamp 1666464484
transform 1 0 90988 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_989
timestamp 1666464484
transform 1 0 92092 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_1001
timestamp 1666464484
transform 1 0 93196 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1007
timestamp 1666464484
transform 1 0 93748 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1009
timestamp 1666464484
transform 1 0 93932 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1021
timestamp 1666464484
transform 1 0 95036 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1033
timestamp 1666464484
transform 1 0 96140 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1045
timestamp 1666464484
transform 1 0 97244 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_1057
timestamp 1666464484
transform 1 0 98348 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1063
timestamp 1666464484
transform 1 0 98900 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1065
timestamp 1666464484
transform 1 0 99084 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1077
timestamp 1666464484
transform 1 0 100188 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1089
timestamp 1666464484
transform 1 0 101292 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1101
timestamp 1666464484
transform 1 0 102396 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_1113
timestamp 1666464484
transform 1 0 103500 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1119
timestamp 1666464484
transform 1 0 104052 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1121
timestamp 1666464484
transform 1 0 104236 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1133
timestamp 1666464484
transform 1 0 105340 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1145
timestamp 1666464484
transform 1 0 106444 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1157
timestamp 1666464484
transform 1 0 107548 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_1169
timestamp 1666464484
transform 1 0 108652 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1175
timestamp 1666464484
transform 1 0 109204 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1177
timestamp 1666464484
transform 1 0 109388 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1189
timestamp 1666464484
transform 1 0 110492 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1201
timestamp 1666464484
transform 1 0 111596 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1213
timestamp 1666464484
transform 1 0 112700 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_1225
timestamp 1666464484
transform 1 0 113804 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1231
timestamp 1666464484
transform 1 0 114356 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1233
timestamp 1666464484
transform 1 0 114540 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1245
timestamp 1666464484
transform 1 0 115644 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1257
timestamp 1666464484
transform 1 0 116748 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1269
timestamp 1666464484
transform 1 0 117852 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_1281
timestamp 1666464484
transform 1 0 118956 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1287
timestamp 1666464484
transform 1 0 119508 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1289
timestamp 1666464484
transform 1 0 119692 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1301
timestamp 1666464484
transform 1 0 120796 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1313
timestamp 1666464484
transform 1 0 121900 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1325
timestamp 1666464484
transform 1 0 123004 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_1337
timestamp 1666464484
transform 1 0 124108 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1343
timestamp 1666464484
transform 1 0 124660 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1345
timestamp 1666464484
transform 1 0 124844 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1357
timestamp 1666464484
transform 1 0 125948 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1369
timestamp 1666464484
transform 1 0 127052 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1381
timestamp 1666464484
transform 1 0 128156 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_1393
timestamp 1666464484
transform 1 0 129260 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1399
timestamp 1666464484
transform 1 0 129812 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1401
timestamp 1666464484
transform 1 0 129996 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1413
timestamp 1666464484
transform 1 0 131100 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1425
timestamp 1666464484
transform 1 0 132204 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1437
timestamp 1666464484
transform 1 0 133308 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_1449
timestamp 1666464484
transform 1 0 134412 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1455
timestamp 1666464484
transform 1 0 134964 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1457
timestamp 1666464484
transform 1 0 135148 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1469
timestamp 1666464484
transform 1 0 136252 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1481
timestamp 1666464484
transform 1 0 137356 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1493
timestamp 1666464484
transform 1 0 138460 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_1505
timestamp 1666464484
transform 1 0 139564 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1511
timestamp 1666464484
transform 1 0 140116 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1513
timestamp 1666464484
transform 1 0 140300 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1525
timestamp 1666464484
transform 1 0 141404 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1537
timestamp 1666464484
transform 1 0 142508 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1549
timestamp 1666464484
transform 1 0 143612 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_1561
timestamp 1666464484
transform 1 0 144716 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1567
timestamp 1666464484
transform 1 0 145268 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1569
timestamp 1666464484
transform 1 0 145452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1581
timestamp 1666464484
transform 1 0 146556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_1593
timestamp 1666464484
transform 1 0 147660 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_1601
timestamp 1666464484
transform 1 0 148396 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1666464484
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1666464484
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1666464484
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1666464484
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1666464484
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1666464484
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1666464484
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1666464484
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1666464484
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1666464484
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1666464484
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1666464484
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1666464484
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1666464484
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1666464484
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1666464484
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1666464484
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1666464484
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1666464484
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1666464484
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1666464484
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1666464484
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1666464484
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1666464484
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1666464484
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1666464484
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1666464484
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1666464484
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1666464484
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1666464484
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1666464484
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1666464484
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1666464484
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1666464484
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1666464484
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1666464484
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1666464484
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1666464484
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1666464484
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1666464484
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1666464484
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1666464484
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1666464484
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1666464484
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1666464484
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1666464484
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1666464484
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1666464484
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1666464484
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1666464484
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1666464484
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1666464484
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1666464484
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1666464484
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1666464484
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1666464484
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1666464484
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1666464484
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1666464484
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1666464484
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1666464484
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1666464484
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1666464484
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1666464484
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1666464484
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_613
timestamp 1666464484
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_625
timestamp 1666464484
transform 1 0 58604 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_637
timestamp 1666464484
transform 1 0 59708 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_643
timestamp 1666464484
transform 1 0 60260 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_645
timestamp 1666464484
transform 1 0 60444 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_657
timestamp 1666464484
transform 1 0 61548 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_669
timestamp 1666464484
transform 1 0 62652 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_681
timestamp 1666464484
transform 1 0 63756 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_693
timestamp 1666464484
transform 1 0 64860 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_699
timestamp 1666464484
transform 1 0 65412 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_701
timestamp 1666464484
transform 1 0 65596 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_713
timestamp 1666464484
transform 1 0 66700 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_725
timestamp 1666464484
transform 1 0 67804 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_737
timestamp 1666464484
transform 1 0 68908 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_749
timestamp 1666464484
transform 1 0 70012 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_755
timestamp 1666464484
transform 1 0 70564 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_757
timestamp 1666464484
transform 1 0 70748 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_769
timestamp 1666464484
transform 1 0 71852 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_781
timestamp 1666464484
transform 1 0 72956 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_793
timestamp 1666464484
transform 1 0 74060 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_805
timestamp 1666464484
transform 1 0 75164 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_811
timestamp 1666464484
transform 1 0 75716 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_813
timestamp 1666464484
transform 1 0 75900 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_825
timestamp 1666464484
transform 1 0 77004 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_837
timestamp 1666464484
transform 1 0 78108 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_849
timestamp 1666464484
transform 1 0 79212 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_861
timestamp 1666464484
transform 1 0 80316 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_867
timestamp 1666464484
transform 1 0 80868 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_869
timestamp 1666464484
transform 1 0 81052 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_881
timestamp 1666464484
transform 1 0 82156 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_893
timestamp 1666464484
transform 1 0 83260 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_905
timestamp 1666464484
transform 1 0 84364 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_917
timestamp 1666464484
transform 1 0 85468 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_923
timestamp 1666464484
transform 1 0 86020 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_925
timestamp 1666464484
transform 1 0 86204 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_937
timestamp 1666464484
transform 1 0 87308 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_949
timestamp 1666464484
transform 1 0 88412 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_961
timestamp 1666464484
transform 1 0 89516 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_973
timestamp 1666464484
transform 1 0 90620 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_979
timestamp 1666464484
transform 1 0 91172 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_981
timestamp 1666464484
transform 1 0 91356 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_993
timestamp 1666464484
transform 1 0 92460 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1005
timestamp 1666464484
transform 1 0 93564 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1017
timestamp 1666464484
transform 1 0 94668 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1029
timestamp 1666464484
transform 1 0 95772 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1035
timestamp 1666464484
transform 1 0 96324 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1037
timestamp 1666464484
transform 1 0 96508 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1049
timestamp 1666464484
transform 1 0 97612 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1061
timestamp 1666464484
transform 1 0 98716 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1073
timestamp 1666464484
transform 1 0 99820 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1085
timestamp 1666464484
transform 1 0 100924 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1091
timestamp 1666464484
transform 1 0 101476 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1093
timestamp 1666464484
transform 1 0 101660 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1105
timestamp 1666464484
transform 1 0 102764 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1117
timestamp 1666464484
transform 1 0 103868 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1129
timestamp 1666464484
transform 1 0 104972 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1141
timestamp 1666464484
transform 1 0 106076 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1147
timestamp 1666464484
transform 1 0 106628 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1149
timestamp 1666464484
transform 1 0 106812 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1161
timestamp 1666464484
transform 1 0 107916 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1173
timestamp 1666464484
transform 1 0 109020 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1185
timestamp 1666464484
transform 1 0 110124 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1197
timestamp 1666464484
transform 1 0 111228 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1203
timestamp 1666464484
transform 1 0 111780 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1205
timestamp 1666464484
transform 1 0 111964 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1217
timestamp 1666464484
transform 1 0 113068 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1229
timestamp 1666464484
transform 1 0 114172 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1241
timestamp 1666464484
transform 1 0 115276 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1253
timestamp 1666464484
transform 1 0 116380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1259
timestamp 1666464484
transform 1 0 116932 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1261
timestamp 1666464484
transform 1 0 117116 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1273
timestamp 1666464484
transform 1 0 118220 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1285
timestamp 1666464484
transform 1 0 119324 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1297
timestamp 1666464484
transform 1 0 120428 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1309
timestamp 1666464484
transform 1 0 121532 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1315
timestamp 1666464484
transform 1 0 122084 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1317
timestamp 1666464484
transform 1 0 122268 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1329
timestamp 1666464484
transform 1 0 123372 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1341
timestamp 1666464484
transform 1 0 124476 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1353
timestamp 1666464484
transform 1 0 125580 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1365
timestamp 1666464484
transform 1 0 126684 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1371
timestamp 1666464484
transform 1 0 127236 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1373
timestamp 1666464484
transform 1 0 127420 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1385
timestamp 1666464484
transform 1 0 128524 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1397
timestamp 1666464484
transform 1 0 129628 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1409
timestamp 1666464484
transform 1 0 130732 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1421
timestamp 1666464484
transform 1 0 131836 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1427
timestamp 1666464484
transform 1 0 132388 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1429
timestamp 1666464484
transform 1 0 132572 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1441
timestamp 1666464484
transform 1 0 133676 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1453
timestamp 1666464484
transform 1 0 134780 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1465
timestamp 1666464484
transform 1 0 135884 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1477
timestamp 1666464484
transform 1 0 136988 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1483
timestamp 1666464484
transform 1 0 137540 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1485
timestamp 1666464484
transform 1 0 137724 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1497
timestamp 1666464484
transform 1 0 138828 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1509
timestamp 1666464484
transform 1 0 139932 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1521
timestamp 1666464484
transform 1 0 141036 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1533
timestamp 1666464484
transform 1 0 142140 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1539
timestamp 1666464484
transform 1 0 142692 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1541
timestamp 1666464484
transform 1 0 142876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1553
timestamp 1666464484
transform 1 0 143980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1565
timestamp 1666464484
transform 1 0 145084 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1577
timestamp 1666464484
transform 1 0 146188 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1589
timestamp 1666464484
transform 1 0 147292 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1595
timestamp 1666464484
transform 1 0 147844 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1597
timestamp 1666464484
transform 1 0 148028 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1666464484
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1666464484
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1666464484
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1666464484
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1666464484
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1666464484
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1666464484
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1666464484
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1666464484
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1666464484
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1666464484
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1666464484
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1666464484
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1666464484
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1666464484
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1666464484
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1666464484
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1666464484
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1666464484
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1666464484
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1666464484
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1666464484
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1666464484
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1666464484
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1666464484
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1666464484
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1666464484
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1666464484
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1666464484
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1666464484
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1666464484
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1666464484
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1666464484
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1666464484
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1666464484
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1666464484
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1666464484
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1666464484
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1666464484
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1666464484
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1666464484
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1666464484
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1666464484
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1666464484
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1666464484
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1666464484
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1666464484
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1666464484
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1666464484
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1666464484
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1666464484
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1666464484
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1666464484
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1666464484
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1666464484
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1666464484
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1666464484
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1666464484
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1666464484
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1666464484
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1666464484
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1666464484
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1666464484
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1666464484
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1666464484
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1666464484
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_617
timestamp 1666464484
transform 1 0 57868 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_629
timestamp 1666464484
transform 1 0 58972 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_641
timestamp 1666464484
transform 1 0 60076 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_653
timestamp 1666464484
transform 1 0 61180 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_665
timestamp 1666464484
transform 1 0 62284 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_671
timestamp 1666464484
transform 1 0 62836 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_673
timestamp 1666464484
transform 1 0 63020 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_685
timestamp 1666464484
transform 1 0 64124 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_697
timestamp 1666464484
transform 1 0 65228 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_709
timestamp 1666464484
transform 1 0 66332 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_721
timestamp 1666464484
transform 1 0 67436 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_727
timestamp 1666464484
transform 1 0 67988 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_729
timestamp 1666464484
transform 1 0 68172 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_741
timestamp 1666464484
transform 1 0 69276 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_753
timestamp 1666464484
transform 1 0 70380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_765
timestamp 1666464484
transform 1 0 71484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_777
timestamp 1666464484
transform 1 0 72588 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_783
timestamp 1666464484
transform 1 0 73140 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_785
timestamp 1666464484
transform 1 0 73324 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_797
timestamp 1666464484
transform 1 0 74428 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_809
timestamp 1666464484
transform 1 0 75532 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_821
timestamp 1666464484
transform 1 0 76636 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_833
timestamp 1666464484
transform 1 0 77740 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_839
timestamp 1666464484
transform 1 0 78292 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_841
timestamp 1666464484
transform 1 0 78476 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_853
timestamp 1666464484
transform 1 0 79580 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_865
timestamp 1666464484
transform 1 0 80684 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_877
timestamp 1666464484
transform 1 0 81788 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_889
timestamp 1666464484
transform 1 0 82892 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_895
timestamp 1666464484
transform 1 0 83444 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_897
timestamp 1666464484
transform 1 0 83628 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_909
timestamp 1666464484
transform 1 0 84732 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_921
timestamp 1666464484
transform 1 0 85836 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_933
timestamp 1666464484
transform 1 0 86940 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_945
timestamp 1666464484
transform 1 0 88044 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_951
timestamp 1666464484
transform 1 0 88596 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_953
timestamp 1666464484
transform 1 0 88780 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_965
timestamp 1666464484
transform 1 0 89884 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_977
timestamp 1666464484
transform 1 0 90988 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_989
timestamp 1666464484
transform 1 0 92092 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1001
timestamp 1666464484
transform 1 0 93196 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1007
timestamp 1666464484
transform 1 0 93748 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1009
timestamp 1666464484
transform 1 0 93932 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1021
timestamp 1666464484
transform 1 0 95036 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1033
timestamp 1666464484
transform 1 0 96140 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1045
timestamp 1666464484
transform 1 0 97244 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1057
timestamp 1666464484
transform 1 0 98348 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1063
timestamp 1666464484
transform 1 0 98900 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1065
timestamp 1666464484
transform 1 0 99084 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1077
timestamp 1666464484
transform 1 0 100188 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1089
timestamp 1666464484
transform 1 0 101292 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1101
timestamp 1666464484
transform 1 0 102396 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1113
timestamp 1666464484
transform 1 0 103500 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1119
timestamp 1666464484
transform 1 0 104052 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1121
timestamp 1666464484
transform 1 0 104236 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1133
timestamp 1666464484
transform 1 0 105340 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1145
timestamp 1666464484
transform 1 0 106444 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1157
timestamp 1666464484
transform 1 0 107548 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1169
timestamp 1666464484
transform 1 0 108652 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1175
timestamp 1666464484
transform 1 0 109204 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1177
timestamp 1666464484
transform 1 0 109388 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1189
timestamp 1666464484
transform 1 0 110492 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1201
timestamp 1666464484
transform 1 0 111596 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1213
timestamp 1666464484
transform 1 0 112700 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1225
timestamp 1666464484
transform 1 0 113804 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1231
timestamp 1666464484
transform 1 0 114356 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1233
timestamp 1666464484
transform 1 0 114540 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1245
timestamp 1666464484
transform 1 0 115644 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1257
timestamp 1666464484
transform 1 0 116748 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1269
timestamp 1666464484
transform 1 0 117852 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1281
timestamp 1666464484
transform 1 0 118956 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1287
timestamp 1666464484
transform 1 0 119508 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1289
timestamp 1666464484
transform 1 0 119692 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1301
timestamp 1666464484
transform 1 0 120796 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1313
timestamp 1666464484
transform 1 0 121900 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1325
timestamp 1666464484
transform 1 0 123004 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1337
timestamp 1666464484
transform 1 0 124108 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1343
timestamp 1666464484
transform 1 0 124660 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1345
timestamp 1666464484
transform 1 0 124844 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1357
timestamp 1666464484
transform 1 0 125948 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1369
timestamp 1666464484
transform 1 0 127052 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1381
timestamp 1666464484
transform 1 0 128156 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1393
timestamp 1666464484
transform 1 0 129260 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1399
timestamp 1666464484
transform 1 0 129812 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1401
timestamp 1666464484
transform 1 0 129996 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1413
timestamp 1666464484
transform 1 0 131100 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1425
timestamp 1666464484
transform 1 0 132204 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1437
timestamp 1666464484
transform 1 0 133308 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1449
timestamp 1666464484
transform 1 0 134412 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1455
timestamp 1666464484
transform 1 0 134964 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1457
timestamp 1666464484
transform 1 0 135148 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1469
timestamp 1666464484
transform 1 0 136252 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1481
timestamp 1666464484
transform 1 0 137356 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1493
timestamp 1666464484
transform 1 0 138460 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1505
timestamp 1666464484
transform 1 0 139564 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1511
timestamp 1666464484
transform 1 0 140116 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1513
timestamp 1666464484
transform 1 0 140300 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1525
timestamp 1666464484
transform 1 0 141404 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1537
timestamp 1666464484
transform 1 0 142508 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1549
timestamp 1666464484
transform 1 0 143612 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1561
timestamp 1666464484
transform 1 0 144716 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1567
timestamp 1666464484
transform 1 0 145268 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1569
timestamp 1666464484
transform 1 0 145452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1581
timestamp 1666464484
transform 1 0 146556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_1593
timestamp 1666464484
transform 1 0 147660 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_1601
timestamp 1666464484
transform 1 0 148396 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1666464484
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1666464484
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1666464484
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1666464484
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1666464484
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1666464484
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1666464484
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1666464484
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1666464484
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1666464484
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1666464484
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1666464484
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1666464484
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1666464484
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1666464484
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1666464484
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1666464484
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1666464484
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1666464484
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1666464484
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1666464484
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1666464484
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1666464484
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1666464484
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1666464484
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1666464484
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1666464484
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1666464484
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1666464484
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1666464484
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1666464484
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1666464484
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1666464484
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1666464484
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1666464484
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1666464484
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1666464484
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1666464484
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1666464484
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1666464484
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1666464484
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1666464484
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1666464484
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1666464484
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1666464484
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1666464484
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1666464484
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1666464484
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1666464484
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1666464484
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1666464484
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1666464484
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1666464484
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1666464484
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1666464484
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1666464484
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1666464484
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1666464484
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1666464484
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1666464484
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1666464484
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1666464484
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1666464484
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1666464484
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1666464484
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_613
timestamp 1666464484
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_625
timestamp 1666464484
transform 1 0 58604 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_637
timestamp 1666464484
transform 1 0 59708 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_643
timestamp 1666464484
transform 1 0 60260 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_645
timestamp 1666464484
transform 1 0 60444 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_657
timestamp 1666464484
transform 1 0 61548 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_669
timestamp 1666464484
transform 1 0 62652 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_681
timestamp 1666464484
transform 1 0 63756 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_693
timestamp 1666464484
transform 1 0 64860 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_699
timestamp 1666464484
transform 1 0 65412 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_701
timestamp 1666464484
transform 1 0 65596 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_713
timestamp 1666464484
transform 1 0 66700 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_725
timestamp 1666464484
transform 1 0 67804 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_737
timestamp 1666464484
transform 1 0 68908 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_749
timestamp 1666464484
transform 1 0 70012 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_755
timestamp 1666464484
transform 1 0 70564 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_757
timestamp 1666464484
transform 1 0 70748 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_769
timestamp 1666464484
transform 1 0 71852 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_781
timestamp 1666464484
transform 1 0 72956 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_793
timestamp 1666464484
transform 1 0 74060 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_805
timestamp 1666464484
transform 1 0 75164 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_811
timestamp 1666464484
transform 1 0 75716 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_813
timestamp 1666464484
transform 1 0 75900 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_825
timestamp 1666464484
transform 1 0 77004 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_837
timestamp 1666464484
transform 1 0 78108 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_849
timestamp 1666464484
transform 1 0 79212 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_861
timestamp 1666464484
transform 1 0 80316 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_867
timestamp 1666464484
transform 1 0 80868 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_869
timestamp 1666464484
transform 1 0 81052 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_881
timestamp 1666464484
transform 1 0 82156 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_893
timestamp 1666464484
transform 1 0 83260 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_905
timestamp 1666464484
transform 1 0 84364 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_917
timestamp 1666464484
transform 1 0 85468 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_923
timestamp 1666464484
transform 1 0 86020 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_925
timestamp 1666464484
transform 1 0 86204 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_937
timestamp 1666464484
transform 1 0 87308 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_949
timestamp 1666464484
transform 1 0 88412 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_961
timestamp 1666464484
transform 1 0 89516 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_973
timestamp 1666464484
transform 1 0 90620 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_979
timestamp 1666464484
transform 1 0 91172 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_981
timestamp 1666464484
transform 1 0 91356 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_993
timestamp 1666464484
transform 1 0 92460 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1005
timestamp 1666464484
transform 1 0 93564 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1017
timestamp 1666464484
transform 1 0 94668 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1029
timestamp 1666464484
transform 1 0 95772 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1035
timestamp 1666464484
transform 1 0 96324 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1037
timestamp 1666464484
transform 1 0 96508 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1049
timestamp 1666464484
transform 1 0 97612 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1061
timestamp 1666464484
transform 1 0 98716 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1073
timestamp 1666464484
transform 1 0 99820 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1085
timestamp 1666464484
transform 1 0 100924 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1091
timestamp 1666464484
transform 1 0 101476 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1093
timestamp 1666464484
transform 1 0 101660 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1105
timestamp 1666464484
transform 1 0 102764 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1117
timestamp 1666464484
transform 1 0 103868 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1129
timestamp 1666464484
transform 1 0 104972 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1141
timestamp 1666464484
transform 1 0 106076 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1147
timestamp 1666464484
transform 1 0 106628 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1149
timestamp 1666464484
transform 1 0 106812 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1161
timestamp 1666464484
transform 1 0 107916 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1173
timestamp 1666464484
transform 1 0 109020 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1185
timestamp 1666464484
transform 1 0 110124 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1197
timestamp 1666464484
transform 1 0 111228 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1203
timestamp 1666464484
transform 1 0 111780 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1205
timestamp 1666464484
transform 1 0 111964 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1217
timestamp 1666464484
transform 1 0 113068 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1229
timestamp 1666464484
transform 1 0 114172 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1241
timestamp 1666464484
transform 1 0 115276 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1253
timestamp 1666464484
transform 1 0 116380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1259
timestamp 1666464484
transform 1 0 116932 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1261
timestamp 1666464484
transform 1 0 117116 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1273
timestamp 1666464484
transform 1 0 118220 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1285
timestamp 1666464484
transform 1 0 119324 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1297
timestamp 1666464484
transform 1 0 120428 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1309
timestamp 1666464484
transform 1 0 121532 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1315
timestamp 1666464484
transform 1 0 122084 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1317
timestamp 1666464484
transform 1 0 122268 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1329
timestamp 1666464484
transform 1 0 123372 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1341
timestamp 1666464484
transform 1 0 124476 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1353
timestamp 1666464484
transform 1 0 125580 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1365
timestamp 1666464484
transform 1 0 126684 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1371
timestamp 1666464484
transform 1 0 127236 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1373
timestamp 1666464484
transform 1 0 127420 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1385
timestamp 1666464484
transform 1 0 128524 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1397
timestamp 1666464484
transform 1 0 129628 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1409
timestamp 1666464484
transform 1 0 130732 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1421
timestamp 1666464484
transform 1 0 131836 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1427
timestamp 1666464484
transform 1 0 132388 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1429
timestamp 1666464484
transform 1 0 132572 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1441
timestamp 1666464484
transform 1 0 133676 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1453
timestamp 1666464484
transform 1 0 134780 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1465
timestamp 1666464484
transform 1 0 135884 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1477
timestamp 1666464484
transform 1 0 136988 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1483
timestamp 1666464484
transform 1 0 137540 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1485
timestamp 1666464484
transform 1 0 137724 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1497
timestamp 1666464484
transform 1 0 138828 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1509
timestamp 1666464484
transform 1 0 139932 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1521
timestamp 1666464484
transform 1 0 141036 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1533
timestamp 1666464484
transform 1 0 142140 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1539
timestamp 1666464484
transform 1 0 142692 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1541
timestamp 1666464484
transform 1 0 142876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1553
timestamp 1666464484
transform 1 0 143980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1565
timestamp 1666464484
transform 1 0 145084 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1577
timestamp 1666464484
transform 1 0 146188 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1589
timestamp 1666464484
transform 1 0 147292 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1595
timestamp 1666464484
transform 1 0 147844 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1597
timestamp 1666464484
transform 1 0 148028 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1666464484
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1666464484
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1666464484
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1666464484
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1666464484
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1666464484
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1666464484
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1666464484
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1666464484
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1666464484
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1666464484
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1666464484
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1666464484
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1666464484
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1666464484
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1666464484
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1666464484
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1666464484
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1666464484
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1666464484
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1666464484
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1666464484
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1666464484
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1666464484
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1666464484
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1666464484
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1666464484
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1666464484
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1666464484
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1666464484
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1666464484
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1666464484
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1666464484
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1666464484
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1666464484
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1666464484
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1666464484
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1666464484
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1666464484
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1666464484
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1666464484
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1666464484
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1666464484
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1666464484
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1666464484
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1666464484
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1666464484
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1666464484
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1666464484
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1666464484
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1666464484
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1666464484
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1666464484
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1666464484
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1666464484
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1666464484
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1666464484
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1666464484
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1666464484
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1666464484
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1666464484
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1666464484
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1666464484
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_597
timestamp 1666464484
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1666464484
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1666464484
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_617
timestamp 1666464484
transform 1 0 57868 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_629
timestamp 1666464484
transform 1 0 58972 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_641
timestamp 1666464484
transform 1 0 60076 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_653
timestamp 1666464484
transform 1 0 61180 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_665
timestamp 1666464484
transform 1 0 62284 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_671
timestamp 1666464484
transform 1 0 62836 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_673
timestamp 1666464484
transform 1 0 63020 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_685
timestamp 1666464484
transform 1 0 64124 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_697
timestamp 1666464484
transform 1 0 65228 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_709
timestamp 1666464484
transform 1 0 66332 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_721
timestamp 1666464484
transform 1 0 67436 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_727
timestamp 1666464484
transform 1 0 67988 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_729
timestamp 1666464484
transform 1 0 68172 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_741
timestamp 1666464484
transform 1 0 69276 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_753
timestamp 1666464484
transform 1 0 70380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_765
timestamp 1666464484
transform 1 0 71484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_777
timestamp 1666464484
transform 1 0 72588 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_783
timestamp 1666464484
transform 1 0 73140 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_785
timestamp 1666464484
transform 1 0 73324 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_797
timestamp 1666464484
transform 1 0 74428 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_809
timestamp 1666464484
transform 1 0 75532 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_821
timestamp 1666464484
transform 1 0 76636 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_833
timestamp 1666464484
transform 1 0 77740 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_839
timestamp 1666464484
transform 1 0 78292 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_841
timestamp 1666464484
transform 1 0 78476 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_853
timestamp 1666464484
transform 1 0 79580 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_865
timestamp 1666464484
transform 1 0 80684 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_877
timestamp 1666464484
transform 1 0 81788 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_889
timestamp 1666464484
transform 1 0 82892 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_895
timestamp 1666464484
transform 1 0 83444 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_897
timestamp 1666464484
transform 1 0 83628 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_909
timestamp 1666464484
transform 1 0 84732 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_921
timestamp 1666464484
transform 1 0 85836 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_933
timestamp 1666464484
transform 1 0 86940 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_945
timestamp 1666464484
transform 1 0 88044 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_951
timestamp 1666464484
transform 1 0 88596 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_953
timestamp 1666464484
transform 1 0 88780 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_965
timestamp 1666464484
transform 1 0 89884 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_977
timestamp 1666464484
transform 1 0 90988 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_989
timestamp 1666464484
transform 1 0 92092 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1001
timestamp 1666464484
transform 1 0 93196 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1007
timestamp 1666464484
transform 1 0 93748 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1009
timestamp 1666464484
transform 1 0 93932 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1021
timestamp 1666464484
transform 1 0 95036 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1033
timestamp 1666464484
transform 1 0 96140 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1045
timestamp 1666464484
transform 1 0 97244 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1057
timestamp 1666464484
transform 1 0 98348 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1063
timestamp 1666464484
transform 1 0 98900 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1065
timestamp 1666464484
transform 1 0 99084 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1077
timestamp 1666464484
transform 1 0 100188 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1089
timestamp 1666464484
transform 1 0 101292 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1101
timestamp 1666464484
transform 1 0 102396 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1113
timestamp 1666464484
transform 1 0 103500 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1119
timestamp 1666464484
transform 1 0 104052 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1121
timestamp 1666464484
transform 1 0 104236 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1133
timestamp 1666464484
transform 1 0 105340 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1145
timestamp 1666464484
transform 1 0 106444 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1157
timestamp 1666464484
transform 1 0 107548 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1169
timestamp 1666464484
transform 1 0 108652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1175
timestamp 1666464484
transform 1 0 109204 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1177
timestamp 1666464484
transform 1 0 109388 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1189
timestamp 1666464484
transform 1 0 110492 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1201
timestamp 1666464484
transform 1 0 111596 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1213
timestamp 1666464484
transform 1 0 112700 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1225
timestamp 1666464484
transform 1 0 113804 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1231
timestamp 1666464484
transform 1 0 114356 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1233
timestamp 1666464484
transform 1 0 114540 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1245
timestamp 1666464484
transform 1 0 115644 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1257
timestamp 1666464484
transform 1 0 116748 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1269
timestamp 1666464484
transform 1 0 117852 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1281
timestamp 1666464484
transform 1 0 118956 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1287
timestamp 1666464484
transform 1 0 119508 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1289
timestamp 1666464484
transform 1 0 119692 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1301
timestamp 1666464484
transform 1 0 120796 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1313
timestamp 1666464484
transform 1 0 121900 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1325
timestamp 1666464484
transform 1 0 123004 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1337
timestamp 1666464484
transform 1 0 124108 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1343
timestamp 1666464484
transform 1 0 124660 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1345
timestamp 1666464484
transform 1 0 124844 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1357
timestamp 1666464484
transform 1 0 125948 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1369
timestamp 1666464484
transform 1 0 127052 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1381
timestamp 1666464484
transform 1 0 128156 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1393
timestamp 1666464484
transform 1 0 129260 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1399
timestamp 1666464484
transform 1 0 129812 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1401
timestamp 1666464484
transform 1 0 129996 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1413
timestamp 1666464484
transform 1 0 131100 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1425
timestamp 1666464484
transform 1 0 132204 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1437
timestamp 1666464484
transform 1 0 133308 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1449
timestamp 1666464484
transform 1 0 134412 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1455
timestamp 1666464484
transform 1 0 134964 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1457
timestamp 1666464484
transform 1 0 135148 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1469
timestamp 1666464484
transform 1 0 136252 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1481
timestamp 1666464484
transform 1 0 137356 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1493
timestamp 1666464484
transform 1 0 138460 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1505
timestamp 1666464484
transform 1 0 139564 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1511
timestamp 1666464484
transform 1 0 140116 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1513
timestamp 1666464484
transform 1 0 140300 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1525
timestamp 1666464484
transform 1 0 141404 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1537
timestamp 1666464484
transform 1 0 142508 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1549
timestamp 1666464484
transform 1 0 143612 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1561
timestamp 1666464484
transform 1 0 144716 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1567
timestamp 1666464484
transform 1 0 145268 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1569
timestamp 1666464484
transform 1 0 145452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1581
timestamp 1666464484
transform 1 0 146556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_1593
timestamp 1666464484
transform 1 0 147660 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_1601
timestamp 1666464484
transform 1 0 148396 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1666464484
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1666464484
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1666464484
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1666464484
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1666464484
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1666464484
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1666464484
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1666464484
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1666464484
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1666464484
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1666464484
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1666464484
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1666464484
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1666464484
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1666464484
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1666464484
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1666464484
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1666464484
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1666464484
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1666464484
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1666464484
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1666464484
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1666464484
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1666464484
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1666464484
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1666464484
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1666464484
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1666464484
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1666464484
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1666464484
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1666464484
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1666464484
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1666464484
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1666464484
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1666464484
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1666464484
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1666464484
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1666464484
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1666464484
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1666464484
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1666464484
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1666464484
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1666464484
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1666464484
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1666464484
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1666464484
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1666464484
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1666464484
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1666464484
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1666464484
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1666464484
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1666464484
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1666464484
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1666464484
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1666464484
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1666464484
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1666464484
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1666464484
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1666464484
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1666464484
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1666464484
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1666464484
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1666464484
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1666464484
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1666464484
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_613
timestamp 1666464484
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_625
timestamp 1666464484
transform 1 0 58604 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_637
timestamp 1666464484
transform 1 0 59708 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_643
timestamp 1666464484
transform 1 0 60260 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_645
timestamp 1666464484
transform 1 0 60444 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_657
timestamp 1666464484
transform 1 0 61548 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_669
timestamp 1666464484
transform 1 0 62652 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_681
timestamp 1666464484
transform 1 0 63756 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_693
timestamp 1666464484
transform 1 0 64860 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_699
timestamp 1666464484
transform 1 0 65412 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_701
timestamp 1666464484
transform 1 0 65596 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_713
timestamp 1666464484
transform 1 0 66700 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_725
timestamp 1666464484
transform 1 0 67804 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_737
timestamp 1666464484
transform 1 0 68908 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_749
timestamp 1666464484
transform 1 0 70012 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_755
timestamp 1666464484
transform 1 0 70564 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_757
timestamp 1666464484
transform 1 0 70748 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_769
timestamp 1666464484
transform 1 0 71852 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_781
timestamp 1666464484
transform 1 0 72956 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_793
timestamp 1666464484
transform 1 0 74060 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_805
timestamp 1666464484
transform 1 0 75164 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_811
timestamp 1666464484
transform 1 0 75716 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_813
timestamp 1666464484
transform 1 0 75900 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_825
timestamp 1666464484
transform 1 0 77004 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_837
timestamp 1666464484
transform 1 0 78108 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_849
timestamp 1666464484
transform 1 0 79212 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_861
timestamp 1666464484
transform 1 0 80316 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_867
timestamp 1666464484
transform 1 0 80868 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_869
timestamp 1666464484
transform 1 0 81052 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_881
timestamp 1666464484
transform 1 0 82156 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_893
timestamp 1666464484
transform 1 0 83260 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_905
timestamp 1666464484
transform 1 0 84364 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_917
timestamp 1666464484
transform 1 0 85468 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_923
timestamp 1666464484
transform 1 0 86020 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_925
timestamp 1666464484
transform 1 0 86204 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_937
timestamp 1666464484
transform 1 0 87308 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_949
timestamp 1666464484
transform 1 0 88412 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_961
timestamp 1666464484
transform 1 0 89516 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_973
timestamp 1666464484
transform 1 0 90620 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_979
timestamp 1666464484
transform 1 0 91172 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_981
timestamp 1666464484
transform 1 0 91356 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_993
timestamp 1666464484
transform 1 0 92460 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1005
timestamp 1666464484
transform 1 0 93564 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1017
timestamp 1666464484
transform 1 0 94668 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1029
timestamp 1666464484
transform 1 0 95772 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1035
timestamp 1666464484
transform 1 0 96324 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1037
timestamp 1666464484
transform 1 0 96508 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1049
timestamp 1666464484
transform 1 0 97612 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1061
timestamp 1666464484
transform 1 0 98716 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1073
timestamp 1666464484
transform 1 0 99820 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1085
timestamp 1666464484
transform 1 0 100924 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1091
timestamp 1666464484
transform 1 0 101476 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1093
timestamp 1666464484
transform 1 0 101660 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1105
timestamp 1666464484
transform 1 0 102764 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1117
timestamp 1666464484
transform 1 0 103868 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1129
timestamp 1666464484
transform 1 0 104972 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1141
timestamp 1666464484
transform 1 0 106076 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1147
timestamp 1666464484
transform 1 0 106628 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1149
timestamp 1666464484
transform 1 0 106812 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1161
timestamp 1666464484
transform 1 0 107916 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1173
timestamp 1666464484
transform 1 0 109020 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1185
timestamp 1666464484
transform 1 0 110124 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1197
timestamp 1666464484
transform 1 0 111228 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1203
timestamp 1666464484
transform 1 0 111780 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1205
timestamp 1666464484
transform 1 0 111964 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1217
timestamp 1666464484
transform 1 0 113068 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1229
timestamp 1666464484
transform 1 0 114172 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1241
timestamp 1666464484
transform 1 0 115276 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1253
timestamp 1666464484
transform 1 0 116380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1259
timestamp 1666464484
transform 1 0 116932 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1261
timestamp 1666464484
transform 1 0 117116 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1273
timestamp 1666464484
transform 1 0 118220 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1285
timestamp 1666464484
transform 1 0 119324 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1297
timestamp 1666464484
transform 1 0 120428 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1309
timestamp 1666464484
transform 1 0 121532 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1315
timestamp 1666464484
transform 1 0 122084 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1317
timestamp 1666464484
transform 1 0 122268 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1329
timestamp 1666464484
transform 1 0 123372 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1341
timestamp 1666464484
transform 1 0 124476 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1353
timestamp 1666464484
transform 1 0 125580 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1365
timestamp 1666464484
transform 1 0 126684 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1371
timestamp 1666464484
transform 1 0 127236 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1373
timestamp 1666464484
transform 1 0 127420 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1385
timestamp 1666464484
transform 1 0 128524 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1397
timestamp 1666464484
transform 1 0 129628 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1409
timestamp 1666464484
transform 1 0 130732 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1421
timestamp 1666464484
transform 1 0 131836 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1427
timestamp 1666464484
transform 1 0 132388 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1429
timestamp 1666464484
transform 1 0 132572 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1441
timestamp 1666464484
transform 1 0 133676 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1453
timestamp 1666464484
transform 1 0 134780 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1465
timestamp 1666464484
transform 1 0 135884 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1477
timestamp 1666464484
transform 1 0 136988 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1483
timestamp 1666464484
transform 1 0 137540 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1485
timestamp 1666464484
transform 1 0 137724 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1497
timestamp 1666464484
transform 1 0 138828 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1509
timestamp 1666464484
transform 1 0 139932 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1521
timestamp 1666464484
transform 1 0 141036 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1533
timestamp 1666464484
transform 1 0 142140 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1539
timestamp 1666464484
transform 1 0 142692 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1541
timestamp 1666464484
transform 1 0 142876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1553
timestamp 1666464484
transform 1 0 143980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1565
timestamp 1666464484
transform 1 0 145084 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1577
timestamp 1666464484
transform 1 0 146188 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1589
timestamp 1666464484
transform 1 0 147292 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1595
timestamp 1666464484
transform 1 0 147844 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1597
timestamp 1666464484
transform 1 0 148028 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1666464484
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1666464484
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1666464484
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1666464484
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1666464484
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1666464484
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1666464484
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1666464484
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1666464484
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1666464484
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1666464484
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1666464484
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1666464484
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1666464484
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1666464484
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1666464484
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1666464484
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1666464484
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1666464484
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1666464484
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1666464484
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1666464484
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1666464484
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1666464484
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1666464484
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1666464484
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1666464484
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1666464484
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1666464484
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1666464484
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1666464484
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1666464484
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1666464484
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1666464484
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1666464484
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1666464484
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1666464484
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1666464484
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1666464484
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1666464484
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1666464484
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1666464484
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1666464484
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1666464484
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1666464484
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1666464484
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1666464484
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1666464484
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1666464484
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1666464484
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1666464484
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1666464484
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1666464484
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1666464484
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1666464484
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1666464484
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1666464484
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1666464484
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1666464484
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1666464484
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1666464484
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1666464484
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1666464484
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1666464484
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1666464484
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1666464484
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_617
timestamp 1666464484
transform 1 0 57868 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_629
timestamp 1666464484
transform 1 0 58972 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_641
timestamp 1666464484
transform 1 0 60076 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_653
timestamp 1666464484
transform 1 0 61180 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_665
timestamp 1666464484
transform 1 0 62284 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_671
timestamp 1666464484
transform 1 0 62836 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_673
timestamp 1666464484
transform 1 0 63020 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_685
timestamp 1666464484
transform 1 0 64124 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_697
timestamp 1666464484
transform 1 0 65228 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_709
timestamp 1666464484
transform 1 0 66332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_721
timestamp 1666464484
transform 1 0 67436 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_727
timestamp 1666464484
transform 1 0 67988 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_729
timestamp 1666464484
transform 1 0 68172 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_741
timestamp 1666464484
transform 1 0 69276 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_753
timestamp 1666464484
transform 1 0 70380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_765
timestamp 1666464484
transform 1 0 71484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_777
timestamp 1666464484
transform 1 0 72588 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_783
timestamp 1666464484
transform 1 0 73140 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_785
timestamp 1666464484
transform 1 0 73324 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_797
timestamp 1666464484
transform 1 0 74428 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_809
timestamp 1666464484
transform 1 0 75532 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_821
timestamp 1666464484
transform 1 0 76636 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_833
timestamp 1666464484
transform 1 0 77740 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_839
timestamp 1666464484
transform 1 0 78292 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_841
timestamp 1666464484
transform 1 0 78476 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_853
timestamp 1666464484
transform 1 0 79580 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_865
timestamp 1666464484
transform 1 0 80684 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_877
timestamp 1666464484
transform 1 0 81788 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_889
timestamp 1666464484
transform 1 0 82892 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_895
timestamp 1666464484
transform 1 0 83444 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_897
timestamp 1666464484
transform 1 0 83628 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_909
timestamp 1666464484
transform 1 0 84732 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_921
timestamp 1666464484
transform 1 0 85836 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_933
timestamp 1666464484
transform 1 0 86940 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_945
timestamp 1666464484
transform 1 0 88044 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_951
timestamp 1666464484
transform 1 0 88596 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_953
timestamp 1666464484
transform 1 0 88780 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_965
timestamp 1666464484
transform 1 0 89884 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_977
timestamp 1666464484
transform 1 0 90988 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_989
timestamp 1666464484
transform 1 0 92092 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_1001
timestamp 1666464484
transform 1 0 93196 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1007
timestamp 1666464484
transform 1 0 93748 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1009
timestamp 1666464484
transform 1 0 93932 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1021
timestamp 1666464484
transform 1 0 95036 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1033
timestamp 1666464484
transform 1 0 96140 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1045
timestamp 1666464484
transform 1 0 97244 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_1057
timestamp 1666464484
transform 1 0 98348 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1063
timestamp 1666464484
transform 1 0 98900 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1065
timestamp 1666464484
transform 1 0 99084 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1077
timestamp 1666464484
transform 1 0 100188 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1089
timestamp 1666464484
transform 1 0 101292 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1101
timestamp 1666464484
transform 1 0 102396 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_1113
timestamp 1666464484
transform 1 0 103500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1119
timestamp 1666464484
transform 1 0 104052 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1121
timestamp 1666464484
transform 1 0 104236 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1133
timestamp 1666464484
transform 1 0 105340 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1145
timestamp 1666464484
transform 1 0 106444 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1157
timestamp 1666464484
transform 1 0 107548 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_1169
timestamp 1666464484
transform 1 0 108652 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1175
timestamp 1666464484
transform 1 0 109204 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1177
timestamp 1666464484
transform 1 0 109388 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1189
timestamp 1666464484
transform 1 0 110492 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1201
timestamp 1666464484
transform 1 0 111596 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1213
timestamp 1666464484
transform 1 0 112700 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_1225
timestamp 1666464484
transform 1 0 113804 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1231
timestamp 1666464484
transform 1 0 114356 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1233
timestamp 1666464484
transform 1 0 114540 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1245
timestamp 1666464484
transform 1 0 115644 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1257
timestamp 1666464484
transform 1 0 116748 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1269
timestamp 1666464484
transform 1 0 117852 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_1281
timestamp 1666464484
transform 1 0 118956 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1287
timestamp 1666464484
transform 1 0 119508 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1289
timestamp 1666464484
transform 1 0 119692 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1301
timestamp 1666464484
transform 1 0 120796 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1313
timestamp 1666464484
transform 1 0 121900 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1325
timestamp 1666464484
transform 1 0 123004 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_1337
timestamp 1666464484
transform 1 0 124108 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1343
timestamp 1666464484
transform 1 0 124660 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1345
timestamp 1666464484
transform 1 0 124844 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1357
timestamp 1666464484
transform 1 0 125948 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1369
timestamp 1666464484
transform 1 0 127052 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1381
timestamp 1666464484
transform 1 0 128156 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_1393
timestamp 1666464484
transform 1 0 129260 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1399
timestamp 1666464484
transform 1 0 129812 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1401
timestamp 1666464484
transform 1 0 129996 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1413
timestamp 1666464484
transform 1 0 131100 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1425
timestamp 1666464484
transform 1 0 132204 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1437
timestamp 1666464484
transform 1 0 133308 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_1449
timestamp 1666464484
transform 1 0 134412 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1455
timestamp 1666464484
transform 1 0 134964 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1457
timestamp 1666464484
transform 1 0 135148 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1469
timestamp 1666464484
transform 1 0 136252 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1481
timestamp 1666464484
transform 1 0 137356 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1493
timestamp 1666464484
transform 1 0 138460 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_1505
timestamp 1666464484
transform 1 0 139564 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1511
timestamp 1666464484
transform 1 0 140116 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1513
timestamp 1666464484
transform 1 0 140300 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1525
timestamp 1666464484
transform 1 0 141404 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1537
timestamp 1666464484
transform 1 0 142508 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1549
timestamp 1666464484
transform 1 0 143612 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_1561
timestamp 1666464484
transform 1 0 144716 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1567
timestamp 1666464484
transform 1 0 145268 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1569
timestamp 1666464484
transform 1 0 145452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1581
timestamp 1666464484
transform 1 0 146556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_1593
timestamp 1666464484
transform 1 0 147660 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_1601
timestamp 1666464484
transform 1 0 148396 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1666464484
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1666464484
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1666464484
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1666464484
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1666464484
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1666464484
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1666464484
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1666464484
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1666464484
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1666464484
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1666464484
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1666464484
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1666464484
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1666464484
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1666464484
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1666464484
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1666464484
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1666464484
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1666464484
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1666464484
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1666464484
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1666464484
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1666464484
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1666464484
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1666464484
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1666464484
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1666464484
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1666464484
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1666464484
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1666464484
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1666464484
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1666464484
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1666464484
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1666464484
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1666464484
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1666464484
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1666464484
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1666464484
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1666464484
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1666464484
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1666464484
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1666464484
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1666464484
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1666464484
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1666464484
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1666464484
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1666464484
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1666464484
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1666464484
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1666464484
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1666464484
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1666464484
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1666464484
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1666464484
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1666464484
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1666464484
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1666464484
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1666464484
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1666464484
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1666464484
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1666464484
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1666464484
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1666464484
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1666464484
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_601
timestamp 1666464484
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_613
timestamp 1666464484
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_625
timestamp 1666464484
transform 1 0 58604 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_637
timestamp 1666464484
transform 1 0 59708 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_643
timestamp 1666464484
transform 1 0 60260 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_645
timestamp 1666464484
transform 1 0 60444 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_657
timestamp 1666464484
transform 1 0 61548 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_669
timestamp 1666464484
transform 1 0 62652 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_681
timestamp 1666464484
transform 1 0 63756 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_693
timestamp 1666464484
transform 1 0 64860 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_699
timestamp 1666464484
transform 1 0 65412 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_701
timestamp 1666464484
transform 1 0 65596 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_713
timestamp 1666464484
transform 1 0 66700 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_725
timestamp 1666464484
transform 1 0 67804 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_737
timestamp 1666464484
transform 1 0 68908 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_749
timestamp 1666464484
transform 1 0 70012 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_755
timestamp 1666464484
transform 1 0 70564 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_757
timestamp 1666464484
transform 1 0 70748 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_769
timestamp 1666464484
transform 1 0 71852 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_781
timestamp 1666464484
transform 1 0 72956 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_793
timestamp 1666464484
transform 1 0 74060 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_805
timestamp 1666464484
transform 1 0 75164 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_811
timestamp 1666464484
transform 1 0 75716 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_813
timestamp 1666464484
transform 1 0 75900 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_825
timestamp 1666464484
transform 1 0 77004 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_837
timestamp 1666464484
transform 1 0 78108 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_849
timestamp 1666464484
transform 1 0 79212 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_861
timestamp 1666464484
transform 1 0 80316 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_867
timestamp 1666464484
transform 1 0 80868 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_869
timestamp 1666464484
transform 1 0 81052 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_881
timestamp 1666464484
transform 1 0 82156 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_893
timestamp 1666464484
transform 1 0 83260 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_905
timestamp 1666464484
transform 1 0 84364 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_917
timestamp 1666464484
transform 1 0 85468 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_923
timestamp 1666464484
transform 1 0 86020 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_925
timestamp 1666464484
transform 1 0 86204 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_937
timestamp 1666464484
transform 1 0 87308 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_949
timestamp 1666464484
transform 1 0 88412 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_961
timestamp 1666464484
transform 1 0 89516 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_973
timestamp 1666464484
transform 1 0 90620 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_979
timestamp 1666464484
transform 1 0 91172 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_981
timestamp 1666464484
transform 1 0 91356 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_993
timestamp 1666464484
transform 1 0 92460 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1005
timestamp 1666464484
transform 1 0 93564 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1017
timestamp 1666464484
transform 1 0 94668 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1029
timestamp 1666464484
transform 1 0 95772 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1035
timestamp 1666464484
transform 1 0 96324 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1037
timestamp 1666464484
transform 1 0 96508 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1049
timestamp 1666464484
transform 1 0 97612 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1061
timestamp 1666464484
transform 1 0 98716 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1073
timestamp 1666464484
transform 1 0 99820 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1085
timestamp 1666464484
transform 1 0 100924 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1091
timestamp 1666464484
transform 1 0 101476 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1093
timestamp 1666464484
transform 1 0 101660 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1105
timestamp 1666464484
transform 1 0 102764 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1117
timestamp 1666464484
transform 1 0 103868 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1129
timestamp 1666464484
transform 1 0 104972 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1141
timestamp 1666464484
transform 1 0 106076 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1147
timestamp 1666464484
transform 1 0 106628 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1149
timestamp 1666464484
transform 1 0 106812 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1161
timestamp 1666464484
transform 1 0 107916 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1173
timestamp 1666464484
transform 1 0 109020 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1185
timestamp 1666464484
transform 1 0 110124 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1197
timestamp 1666464484
transform 1 0 111228 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1203
timestamp 1666464484
transform 1 0 111780 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1205
timestamp 1666464484
transform 1 0 111964 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1217
timestamp 1666464484
transform 1 0 113068 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1229
timestamp 1666464484
transform 1 0 114172 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1241
timestamp 1666464484
transform 1 0 115276 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1253
timestamp 1666464484
transform 1 0 116380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1259
timestamp 1666464484
transform 1 0 116932 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1261
timestamp 1666464484
transform 1 0 117116 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1273
timestamp 1666464484
transform 1 0 118220 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1285
timestamp 1666464484
transform 1 0 119324 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1297
timestamp 1666464484
transform 1 0 120428 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1309
timestamp 1666464484
transform 1 0 121532 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1315
timestamp 1666464484
transform 1 0 122084 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1317
timestamp 1666464484
transform 1 0 122268 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1329
timestamp 1666464484
transform 1 0 123372 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1341
timestamp 1666464484
transform 1 0 124476 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1353
timestamp 1666464484
transform 1 0 125580 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1365
timestamp 1666464484
transform 1 0 126684 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1371
timestamp 1666464484
transform 1 0 127236 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1373
timestamp 1666464484
transform 1 0 127420 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1385
timestamp 1666464484
transform 1 0 128524 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1397
timestamp 1666464484
transform 1 0 129628 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1409
timestamp 1666464484
transform 1 0 130732 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1421
timestamp 1666464484
transform 1 0 131836 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1427
timestamp 1666464484
transform 1 0 132388 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1429
timestamp 1666464484
transform 1 0 132572 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1441
timestamp 1666464484
transform 1 0 133676 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1453
timestamp 1666464484
transform 1 0 134780 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1465
timestamp 1666464484
transform 1 0 135884 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1477
timestamp 1666464484
transform 1 0 136988 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1483
timestamp 1666464484
transform 1 0 137540 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1485
timestamp 1666464484
transform 1 0 137724 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1497
timestamp 1666464484
transform 1 0 138828 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1509
timestamp 1666464484
transform 1 0 139932 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1521
timestamp 1666464484
transform 1 0 141036 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1533
timestamp 1666464484
transform 1 0 142140 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1539
timestamp 1666464484
transform 1 0 142692 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1541
timestamp 1666464484
transform 1 0 142876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1553
timestamp 1666464484
transform 1 0 143980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1565
timestamp 1666464484
transform 1 0 145084 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1577
timestamp 1666464484
transform 1 0 146188 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1589
timestamp 1666464484
transform 1 0 147292 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1595
timestamp 1666464484
transform 1 0 147844 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1597
timestamp 1666464484
transform 1 0 148028 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1666464484
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1666464484
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1666464484
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1666464484
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1666464484
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1666464484
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1666464484
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1666464484
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1666464484
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1666464484
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1666464484
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1666464484
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1666464484
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1666464484
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1666464484
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1666464484
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1666464484
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1666464484
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1666464484
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1666464484
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1666464484
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1666464484
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1666464484
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1666464484
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1666464484
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1666464484
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1666464484
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1666464484
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1666464484
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1666464484
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1666464484
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1666464484
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1666464484
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1666464484
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1666464484
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1666464484
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1666464484
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1666464484
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1666464484
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1666464484
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1666464484
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1666464484
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1666464484
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1666464484
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1666464484
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1666464484
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1666464484
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1666464484
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1666464484
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1666464484
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1666464484
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1666464484
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1666464484
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1666464484
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1666464484
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1666464484
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1666464484
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1666464484
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1666464484
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1666464484
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1666464484
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1666464484
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1666464484
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_597
timestamp 1666464484
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1666464484
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1666464484
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_617
timestamp 1666464484
transform 1 0 57868 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_629
timestamp 1666464484
transform 1 0 58972 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_641
timestamp 1666464484
transform 1 0 60076 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_653
timestamp 1666464484
transform 1 0 61180 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_665
timestamp 1666464484
transform 1 0 62284 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_671
timestamp 1666464484
transform 1 0 62836 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_673
timestamp 1666464484
transform 1 0 63020 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_685
timestamp 1666464484
transform 1 0 64124 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_697
timestamp 1666464484
transform 1 0 65228 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_709
timestamp 1666464484
transform 1 0 66332 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_721
timestamp 1666464484
transform 1 0 67436 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_727
timestamp 1666464484
transform 1 0 67988 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_729
timestamp 1666464484
transform 1 0 68172 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_741
timestamp 1666464484
transform 1 0 69276 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_753
timestamp 1666464484
transform 1 0 70380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_765
timestamp 1666464484
transform 1 0 71484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_777
timestamp 1666464484
transform 1 0 72588 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_783
timestamp 1666464484
transform 1 0 73140 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_785
timestamp 1666464484
transform 1 0 73324 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_797
timestamp 1666464484
transform 1 0 74428 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_809
timestamp 1666464484
transform 1 0 75532 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_821
timestamp 1666464484
transform 1 0 76636 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_833
timestamp 1666464484
transform 1 0 77740 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_839
timestamp 1666464484
transform 1 0 78292 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_841
timestamp 1666464484
transform 1 0 78476 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_853
timestamp 1666464484
transform 1 0 79580 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_865
timestamp 1666464484
transform 1 0 80684 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_877
timestamp 1666464484
transform 1 0 81788 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_889
timestamp 1666464484
transform 1 0 82892 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_895
timestamp 1666464484
transform 1 0 83444 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_897
timestamp 1666464484
transform 1 0 83628 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_909
timestamp 1666464484
transform 1 0 84732 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_921
timestamp 1666464484
transform 1 0 85836 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_933
timestamp 1666464484
transform 1 0 86940 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_945
timestamp 1666464484
transform 1 0 88044 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_951
timestamp 1666464484
transform 1 0 88596 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_953
timestamp 1666464484
transform 1 0 88780 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_965
timestamp 1666464484
transform 1 0 89884 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_977
timestamp 1666464484
transform 1 0 90988 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_989
timestamp 1666464484
transform 1 0 92092 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_1001
timestamp 1666464484
transform 1 0 93196 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1007
timestamp 1666464484
transform 1 0 93748 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1009
timestamp 1666464484
transform 1 0 93932 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1021
timestamp 1666464484
transform 1 0 95036 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1033
timestamp 1666464484
transform 1 0 96140 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1045
timestamp 1666464484
transform 1 0 97244 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_1057
timestamp 1666464484
transform 1 0 98348 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1063
timestamp 1666464484
transform 1 0 98900 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1065
timestamp 1666464484
transform 1 0 99084 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1077
timestamp 1666464484
transform 1 0 100188 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1089
timestamp 1666464484
transform 1 0 101292 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1101
timestamp 1666464484
transform 1 0 102396 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_1113
timestamp 1666464484
transform 1 0 103500 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1119
timestamp 1666464484
transform 1 0 104052 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1121
timestamp 1666464484
transform 1 0 104236 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1133
timestamp 1666464484
transform 1 0 105340 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1145
timestamp 1666464484
transform 1 0 106444 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1157
timestamp 1666464484
transform 1 0 107548 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_1169
timestamp 1666464484
transform 1 0 108652 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1175
timestamp 1666464484
transform 1 0 109204 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1177
timestamp 1666464484
transform 1 0 109388 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1189
timestamp 1666464484
transform 1 0 110492 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1201
timestamp 1666464484
transform 1 0 111596 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1213
timestamp 1666464484
transform 1 0 112700 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_1225
timestamp 1666464484
transform 1 0 113804 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1231
timestamp 1666464484
transform 1 0 114356 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1233
timestamp 1666464484
transform 1 0 114540 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1245
timestamp 1666464484
transform 1 0 115644 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1257
timestamp 1666464484
transform 1 0 116748 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1269
timestamp 1666464484
transform 1 0 117852 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_1281
timestamp 1666464484
transform 1 0 118956 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1287
timestamp 1666464484
transform 1 0 119508 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1289
timestamp 1666464484
transform 1 0 119692 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1301
timestamp 1666464484
transform 1 0 120796 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1313
timestamp 1666464484
transform 1 0 121900 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1325
timestamp 1666464484
transform 1 0 123004 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_1337
timestamp 1666464484
transform 1 0 124108 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1343
timestamp 1666464484
transform 1 0 124660 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1345
timestamp 1666464484
transform 1 0 124844 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1357
timestamp 1666464484
transform 1 0 125948 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1369
timestamp 1666464484
transform 1 0 127052 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1381
timestamp 1666464484
transform 1 0 128156 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_1393
timestamp 1666464484
transform 1 0 129260 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1399
timestamp 1666464484
transform 1 0 129812 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1401
timestamp 1666464484
transform 1 0 129996 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1413
timestamp 1666464484
transform 1 0 131100 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1425
timestamp 1666464484
transform 1 0 132204 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1437
timestamp 1666464484
transform 1 0 133308 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_1449
timestamp 1666464484
transform 1 0 134412 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1455
timestamp 1666464484
transform 1 0 134964 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1457
timestamp 1666464484
transform 1 0 135148 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1469
timestamp 1666464484
transform 1 0 136252 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1481
timestamp 1666464484
transform 1 0 137356 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1493
timestamp 1666464484
transform 1 0 138460 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_1505
timestamp 1666464484
transform 1 0 139564 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1511
timestamp 1666464484
transform 1 0 140116 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1513
timestamp 1666464484
transform 1 0 140300 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1525
timestamp 1666464484
transform 1 0 141404 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1537
timestamp 1666464484
transform 1 0 142508 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1549
timestamp 1666464484
transform 1 0 143612 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_1561
timestamp 1666464484
transform 1 0 144716 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1567
timestamp 1666464484
transform 1 0 145268 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1569
timestamp 1666464484
transform 1 0 145452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1581
timestamp 1666464484
transform 1 0 146556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_1593
timestamp 1666464484
transform 1 0 147660 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_1601
timestamp 1666464484
transform 1 0 148396 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1666464484
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1666464484
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1666464484
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1666464484
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1666464484
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1666464484
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1666464484
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1666464484
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1666464484
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1666464484
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1666464484
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1666464484
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1666464484
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1666464484
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1666464484
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1666464484
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1666464484
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1666464484
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1666464484
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1666464484
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1666464484
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1666464484
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1666464484
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1666464484
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1666464484
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1666464484
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1666464484
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1666464484
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1666464484
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1666464484
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1666464484
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1666464484
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1666464484
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1666464484
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1666464484
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1666464484
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1666464484
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1666464484
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1666464484
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1666464484
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1666464484
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1666464484
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1666464484
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1666464484
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1666464484
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1666464484
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1666464484
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1666464484
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1666464484
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1666464484
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1666464484
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1666464484
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1666464484
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1666464484
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1666464484
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1666464484
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1666464484
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1666464484
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1666464484
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1666464484
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1666464484
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1666464484
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1666464484
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1666464484
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_601
timestamp 1666464484
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_613
timestamp 1666464484
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_625
timestamp 1666464484
transform 1 0 58604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_637
timestamp 1666464484
transform 1 0 59708 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_643
timestamp 1666464484
transform 1 0 60260 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_645
timestamp 1666464484
transform 1 0 60444 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_657
timestamp 1666464484
transform 1 0 61548 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_669
timestamp 1666464484
transform 1 0 62652 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_681
timestamp 1666464484
transform 1 0 63756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_693
timestamp 1666464484
transform 1 0 64860 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_699
timestamp 1666464484
transform 1 0 65412 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_701
timestamp 1666464484
transform 1 0 65596 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_713
timestamp 1666464484
transform 1 0 66700 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_725
timestamp 1666464484
transform 1 0 67804 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_737
timestamp 1666464484
transform 1 0 68908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_749
timestamp 1666464484
transform 1 0 70012 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_755
timestamp 1666464484
transform 1 0 70564 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_757
timestamp 1666464484
transform 1 0 70748 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_769
timestamp 1666464484
transform 1 0 71852 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_781
timestamp 1666464484
transform 1 0 72956 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_793
timestamp 1666464484
transform 1 0 74060 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_805
timestamp 1666464484
transform 1 0 75164 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_811
timestamp 1666464484
transform 1 0 75716 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_813
timestamp 1666464484
transform 1 0 75900 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_825
timestamp 1666464484
transform 1 0 77004 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_837
timestamp 1666464484
transform 1 0 78108 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_849
timestamp 1666464484
transform 1 0 79212 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_861
timestamp 1666464484
transform 1 0 80316 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_867
timestamp 1666464484
transform 1 0 80868 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_869
timestamp 1666464484
transform 1 0 81052 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_881
timestamp 1666464484
transform 1 0 82156 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_893
timestamp 1666464484
transform 1 0 83260 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_905
timestamp 1666464484
transform 1 0 84364 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_917
timestamp 1666464484
transform 1 0 85468 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_923
timestamp 1666464484
transform 1 0 86020 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_925
timestamp 1666464484
transform 1 0 86204 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_937
timestamp 1666464484
transform 1 0 87308 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_949
timestamp 1666464484
transform 1 0 88412 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_961
timestamp 1666464484
transform 1 0 89516 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_973
timestamp 1666464484
transform 1 0 90620 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_979
timestamp 1666464484
transform 1 0 91172 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_981
timestamp 1666464484
transform 1 0 91356 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_993
timestamp 1666464484
transform 1 0 92460 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1005
timestamp 1666464484
transform 1 0 93564 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1017
timestamp 1666464484
transform 1 0 94668 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1029
timestamp 1666464484
transform 1 0 95772 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1035
timestamp 1666464484
transform 1 0 96324 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1037
timestamp 1666464484
transform 1 0 96508 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1049
timestamp 1666464484
transform 1 0 97612 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1061
timestamp 1666464484
transform 1 0 98716 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1073
timestamp 1666464484
transform 1 0 99820 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1085
timestamp 1666464484
transform 1 0 100924 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1091
timestamp 1666464484
transform 1 0 101476 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1093
timestamp 1666464484
transform 1 0 101660 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1105
timestamp 1666464484
transform 1 0 102764 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1117
timestamp 1666464484
transform 1 0 103868 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1129
timestamp 1666464484
transform 1 0 104972 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1141
timestamp 1666464484
transform 1 0 106076 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1147
timestamp 1666464484
transform 1 0 106628 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1149
timestamp 1666464484
transform 1 0 106812 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1161
timestamp 1666464484
transform 1 0 107916 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1173
timestamp 1666464484
transform 1 0 109020 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1185
timestamp 1666464484
transform 1 0 110124 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1197
timestamp 1666464484
transform 1 0 111228 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1203
timestamp 1666464484
transform 1 0 111780 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1205
timestamp 1666464484
transform 1 0 111964 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1217
timestamp 1666464484
transform 1 0 113068 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1229
timestamp 1666464484
transform 1 0 114172 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1241
timestamp 1666464484
transform 1 0 115276 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1253
timestamp 1666464484
transform 1 0 116380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1259
timestamp 1666464484
transform 1 0 116932 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1261
timestamp 1666464484
transform 1 0 117116 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1273
timestamp 1666464484
transform 1 0 118220 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1285
timestamp 1666464484
transform 1 0 119324 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1297
timestamp 1666464484
transform 1 0 120428 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1309
timestamp 1666464484
transform 1 0 121532 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1315
timestamp 1666464484
transform 1 0 122084 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1317
timestamp 1666464484
transform 1 0 122268 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1329
timestamp 1666464484
transform 1 0 123372 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1341
timestamp 1666464484
transform 1 0 124476 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1353
timestamp 1666464484
transform 1 0 125580 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1365
timestamp 1666464484
transform 1 0 126684 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1371
timestamp 1666464484
transform 1 0 127236 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1373
timestamp 1666464484
transform 1 0 127420 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1385
timestamp 1666464484
transform 1 0 128524 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1397
timestamp 1666464484
transform 1 0 129628 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1409
timestamp 1666464484
transform 1 0 130732 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1421
timestamp 1666464484
transform 1 0 131836 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1427
timestamp 1666464484
transform 1 0 132388 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1429
timestamp 1666464484
transform 1 0 132572 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1441
timestamp 1666464484
transform 1 0 133676 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1453
timestamp 1666464484
transform 1 0 134780 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1465
timestamp 1666464484
transform 1 0 135884 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1477
timestamp 1666464484
transform 1 0 136988 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1483
timestamp 1666464484
transform 1 0 137540 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1485
timestamp 1666464484
transform 1 0 137724 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1497
timestamp 1666464484
transform 1 0 138828 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1509
timestamp 1666464484
transform 1 0 139932 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1521
timestamp 1666464484
transform 1 0 141036 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1533
timestamp 1666464484
transform 1 0 142140 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1539
timestamp 1666464484
transform 1 0 142692 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1541
timestamp 1666464484
transform 1 0 142876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1553
timestamp 1666464484
transform 1 0 143980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1565
timestamp 1666464484
transform 1 0 145084 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1577
timestamp 1666464484
transform 1 0 146188 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1589
timestamp 1666464484
transform 1 0 147292 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1595
timestamp 1666464484
transform 1 0 147844 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1597
timestamp 1666464484
transform 1 0 148028 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1666464484
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1666464484
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1666464484
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1666464484
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1666464484
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1666464484
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1666464484
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1666464484
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1666464484
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1666464484
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1666464484
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1666464484
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1666464484
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1666464484
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1666464484
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1666464484
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1666464484
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1666464484
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1666464484
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1666464484
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1666464484
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1666464484
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1666464484
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1666464484
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1666464484
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1666464484
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1666464484
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1666464484
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1666464484
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1666464484
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1666464484
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1666464484
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1666464484
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1666464484
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1666464484
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1666464484
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1666464484
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1666464484
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1666464484
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1666464484
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1666464484
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1666464484
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1666464484
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1666464484
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1666464484
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1666464484
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1666464484
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1666464484
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1666464484
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1666464484
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1666464484
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1666464484
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1666464484
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1666464484
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1666464484
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1666464484
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1666464484
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1666464484
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1666464484
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1666464484
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1666464484
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_573
timestamp 1666464484
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_585
timestamp 1666464484
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_597
timestamp 1666464484
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1666464484
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1666464484
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_617
timestamp 1666464484
transform 1 0 57868 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_629
timestamp 1666464484
transform 1 0 58972 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_641
timestamp 1666464484
transform 1 0 60076 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_653
timestamp 1666464484
transform 1 0 61180 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_665
timestamp 1666464484
transform 1 0 62284 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_671
timestamp 1666464484
transform 1 0 62836 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_673
timestamp 1666464484
transform 1 0 63020 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_685
timestamp 1666464484
transform 1 0 64124 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_697
timestamp 1666464484
transform 1 0 65228 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_709
timestamp 1666464484
transform 1 0 66332 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_721
timestamp 1666464484
transform 1 0 67436 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_727
timestamp 1666464484
transform 1 0 67988 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_729
timestamp 1666464484
transform 1 0 68172 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_741
timestamp 1666464484
transform 1 0 69276 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_753
timestamp 1666464484
transform 1 0 70380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_765
timestamp 1666464484
transform 1 0 71484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_777
timestamp 1666464484
transform 1 0 72588 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_783
timestamp 1666464484
transform 1 0 73140 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_785
timestamp 1666464484
transform 1 0 73324 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_797
timestamp 1666464484
transform 1 0 74428 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_809
timestamp 1666464484
transform 1 0 75532 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_821
timestamp 1666464484
transform 1 0 76636 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_833
timestamp 1666464484
transform 1 0 77740 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_839
timestamp 1666464484
transform 1 0 78292 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_841
timestamp 1666464484
transform 1 0 78476 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_853
timestamp 1666464484
transform 1 0 79580 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_865
timestamp 1666464484
transform 1 0 80684 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_877
timestamp 1666464484
transform 1 0 81788 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_889
timestamp 1666464484
transform 1 0 82892 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_895
timestamp 1666464484
transform 1 0 83444 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_897
timestamp 1666464484
transform 1 0 83628 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_909
timestamp 1666464484
transform 1 0 84732 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_921
timestamp 1666464484
transform 1 0 85836 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_933
timestamp 1666464484
transform 1 0 86940 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_945
timestamp 1666464484
transform 1 0 88044 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_951
timestamp 1666464484
transform 1 0 88596 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_953
timestamp 1666464484
transform 1 0 88780 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_965
timestamp 1666464484
transform 1 0 89884 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_977
timestamp 1666464484
transform 1 0 90988 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_989
timestamp 1666464484
transform 1 0 92092 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_1001
timestamp 1666464484
transform 1 0 93196 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_1007
timestamp 1666464484
transform 1 0 93748 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1009
timestamp 1666464484
transform 1 0 93932 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1021
timestamp 1666464484
transform 1 0 95036 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1033
timestamp 1666464484
transform 1 0 96140 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1045
timestamp 1666464484
transform 1 0 97244 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_1057
timestamp 1666464484
transform 1 0 98348 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_1063
timestamp 1666464484
transform 1 0 98900 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1065
timestamp 1666464484
transform 1 0 99084 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1077
timestamp 1666464484
transform 1 0 100188 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1089
timestamp 1666464484
transform 1 0 101292 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1101
timestamp 1666464484
transform 1 0 102396 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_1113
timestamp 1666464484
transform 1 0 103500 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_1119
timestamp 1666464484
transform 1 0 104052 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1121
timestamp 1666464484
transform 1 0 104236 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1133
timestamp 1666464484
transform 1 0 105340 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1145
timestamp 1666464484
transform 1 0 106444 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1157
timestamp 1666464484
transform 1 0 107548 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_1169
timestamp 1666464484
transform 1 0 108652 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_1175
timestamp 1666464484
transform 1 0 109204 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1177
timestamp 1666464484
transform 1 0 109388 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1189
timestamp 1666464484
transform 1 0 110492 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1201
timestamp 1666464484
transform 1 0 111596 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1213
timestamp 1666464484
transform 1 0 112700 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_1225
timestamp 1666464484
transform 1 0 113804 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_1231
timestamp 1666464484
transform 1 0 114356 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1233
timestamp 1666464484
transform 1 0 114540 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1245
timestamp 1666464484
transform 1 0 115644 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1257
timestamp 1666464484
transform 1 0 116748 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1269
timestamp 1666464484
transform 1 0 117852 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_1281
timestamp 1666464484
transform 1 0 118956 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_1287
timestamp 1666464484
transform 1 0 119508 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1289
timestamp 1666464484
transform 1 0 119692 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1301
timestamp 1666464484
transform 1 0 120796 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1313
timestamp 1666464484
transform 1 0 121900 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1325
timestamp 1666464484
transform 1 0 123004 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_1337
timestamp 1666464484
transform 1 0 124108 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_1343
timestamp 1666464484
transform 1 0 124660 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1345
timestamp 1666464484
transform 1 0 124844 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1357
timestamp 1666464484
transform 1 0 125948 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1369
timestamp 1666464484
transform 1 0 127052 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1381
timestamp 1666464484
transform 1 0 128156 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_1393
timestamp 1666464484
transform 1 0 129260 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_1399
timestamp 1666464484
transform 1 0 129812 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1401
timestamp 1666464484
transform 1 0 129996 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1413
timestamp 1666464484
transform 1 0 131100 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1425
timestamp 1666464484
transform 1 0 132204 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1437
timestamp 1666464484
transform 1 0 133308 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_1449
timestamp 1666464484
transform 1 0 134412 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_1455
timestamp 1666464484
transform 1 0 134964 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1457
timestamp 1666464484
transform 1 0 135148 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1469
timestamp 1666464484
transform 1 0 136252 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1481
timestamp 1666464484
transform 1 0 137356 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1493
timestamp 1666464484
transform 1 0 138460 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_1505
timestamp 1666464484
transform 1 0 139564 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_1511
timestamp 1666464484
transform 1 0 140116 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1513
timestamp 1666464484
transform 1 0 140300 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1525
timestamp 1666464484
transform 1 0 141404 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1537
timestamp 1666464484
transform 1 0 142508 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1549
timestamp 1666464484
transform 1 0 143612 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_1561
timestamp 1666464484
transform 1 0 144716 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_1567
timestamp 1666464484
transform 1 0 145268 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1569
timestamp 1666464484
transform 1 0 145452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1581
timestamp 1666464484
transform 1 0 146556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_1593
timestamp 1666464484
transform 1 0 147660 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_1601
timestamp 1666464484
transform 1 0 148396 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1666464484
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1666464484
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1666464484
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1666464484
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1666464484
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1666464484
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1666464484
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1666464484
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1666464484
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1666464484
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1666464484
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1666464484
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1666464484
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1666464484
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1666464484
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1666464484
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1666464484
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1666464484
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1666464484
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1666464484
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1666464484
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1666464484
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1666464484
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1666464484
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1666464484
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1666464484
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1666464484
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1666464484
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1666464484
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1666464484
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1666464484
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1666464484
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1666464484
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1666464484
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1666464484
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1666464484
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1666464484
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1666464484
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1666464484
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1666464484
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1666464484
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1666464484
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1666464484
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1666464484
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1666464484
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1666464484
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1666464484
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1666464484
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1666464484
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1666464484
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1666464484
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1666464484
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1666464484
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1666464484
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1666464484
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1666464484
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1666464484
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1666464484
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1666464484
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1666464484
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_569
timestamp 1666464484
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1666464484
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1666464484
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1666464484
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_601
timestamp 1666464484
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_613
timestamp 1666464484
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_625
timestamp 1666464484
transform 1 0 58604 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_637
timestamp 1666464484
transform 1 0 59708 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_643
timestamp 1666464484
transform 1 0 60260 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_645
timestamp 1666464484
transform 1 0 60444 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_657
timestamp 1666464484
transform 1 0 61548 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_669
timestamp 1666464484
transform 1 0 62652 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_681
timestamp 1666464484
transform 1 0 63756 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_693
timestamp 1666464484
transform 1 0 64860 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_699
timestamp 1666464484
transform 1 0 65412 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_701
timestamp 1666464484
transform 1 0 65596 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_713
timestamp 1666464484
transform 1 0 66700 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_725
timestamp 1666464484
transform 1 0 67804 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_737
timestamp 1666464484
transform 1 0 68908 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_749
timestamp 1666464484
transform 1 0 70012 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_755
timestamp 1666464484
transform 1 0 70564 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_757
timestamp 1666464484
transform 1 0 70748 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_769
timestamp 1666464484
transform 1 0 71852 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_781
timestamp 1666464484
transform 1 0 72956 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_793
timestamp 1666464484
transform 1 0 74060 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_805
timestamp 1666464484
transform 1 0 75164 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_811
timestamp 1666464484
transform 1 0 75716 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_813
timestamp 1666464484
transform 1 0 75900 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_825
timestamp 1666464484
transform 1 0 77004 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_837
timestamp 1666464484
transform 1 0 78108 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_849
timestamp 1666464484
transform 1 0 79212 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_861
timestamp 1666464484
transform 1 0 80316 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_867
timestamp 1666464484
transform 1 0 80868 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_869
timestamp 1666464484
transform 1 0 81052 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_881
timestamp 1666464484
transform 1 0 82156 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_893
timestamp 1666464484
transform 1 0 83260 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_905
timestamp 1666464484
transform 1 0 84364 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_917
timestamp 1666464484
transform 1 0 85468 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_923
timestamp 1666464484
transform 1 0 86020 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_925
timestamp 1666464484
transform 1 0 86204 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_937
timestamp 1666464484
transform 1 0 87308 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_949
timestamp 1666464484
transform 1 0 88412 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_961
timestamp 1666464484
transform 1 0 89516 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_973
timestamp 1666464484
transform 1 0 90620 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_979
timestamp 1666464484
transform 1 0 91172 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_981
timestamp 1666464484
transform 1 0 91356 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_993
timestamp 1666464484
transform 1 0 92460 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1005
timestamp 1666464484
transform 1 0 93564 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1017
timestamp 1666464484
transform 1 0 94668 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_1029
timestamp 1666464484
transform 1 0 95772 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1035
timestamp 1666464484
transform 1 0 96324 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1037
timestamp 1666464484
transform 1 0 96508 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1049
timestamp 1666464484
transform 1 0 97612 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1061
timestamp 1666464484
transform 1 0 98716 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1073
timestamp 1666464484
transform 1 0 99820 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_1085
timestamp 1666464484
transform 1 0 100924 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1091
timestamp 1666464484
transform 1 0 101476 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1093
timestamp 1666464484
transform 1 0 101660 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1105
timestamp 1666464484
transform 1 0 102764 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1117
timestamp 1666464484
transform 1 0 103868 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1129
timestamp 1666464484
transform 1 0 104972 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_1141
timestamp 1666464484
transform 1 0 106076 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1147
timestamp 1666464484
transform 1 0 106628 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1149
timestamp 1666464484
transform 1 0 106812 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1161
timestamp 1666464484
transform 1 0 107916 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1173
timestamp 1666464484
transform 1 0 109020 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1185
timestamp 1666464484
transform 1 0 110124 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_1197
timestamp 1666464484
transform 1 0 111228 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1203
timestamp 1666464484
transform 1 0 111780 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1205
timestamp 1666464484
transform 1 0 111964 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1217
timestamp 1666464484
transform 1 0 113068 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1229
timestamp 1666464484
transform 1 0 114172 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1241
timestamp 1666464484
transform 1 0 115276 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_1253
timestamp 1666464484
transform 1 0 116380 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1259
timestamp 1666464484
transform 1 0 116932 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1261
timestamp 1666464484
transform 1 0 117116 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1273
timestamp 1666464484
transform 1 0 118220 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1285
timestamp 1666464484
transform 1 0 119324 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1297
timestamp 1666464484
transform 1 0 120428 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_1309
timestamp 1666464484
transform 1 0 121532 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1315
timestamp 1666464484
transform 1 0 122084 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1317
timestamp 1666464484
transform 1 0 122268 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1329
timestamp 1666464484
transform 1 0 123372 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1341
timestamp 1666464484
transform 1 0 124476 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1353
timestamp 1666464484
transform 1 0 125580 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_1365
timestamp 1666464484
transform 1 0 126684 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1371
timestamp 1666464484
transform 1 0 127236 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1373
timestamp 1666464484
transform 1 0 127420 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1385
timestamp 1666464484
transform 1 0 128524 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1397
timestamp 1666464484
transform 1 0 129628 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1409
timestamp 1666464484
transform 1 0 130732 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_1421
timestamp 1666464484
transform 1 0 131836 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1427
timestamp 1666464484
transform 1 0 132388 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1429
timestamp 1666464484
transform 1 0 132572 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1441
timestamp 1666464484
transform 1 0 133676 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1453
timestamp 1666464484
transform 1 0 134780 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1465
timestamp 1666464484
transform 1 0 135884 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_1477
timestamp 1666464484
transform 1 0 136988 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1483
timestamp 1666464484
transform 1 0 137540 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1485
timestamp 1666464484
transform 1 0 137724 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1497
timestamp 1666464484
transform 1 0 138828 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1509
timestamp 1666464484
transform 1 0 139932 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1521
timestamp 1666464484
transform 1 0 141036 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_1533
timestamp 1666464484
transform 1 0 142140 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1539
timestamp 1666464484
transform 1 0 142692 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1541
timestamp 1666464484
transform 1 0 142876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1553
timestamp 1666464484
transform 1 0 143980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1565
timestamp 1666464484
transform 1 0 145084 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1577
timestamp 1666464484
transform 1 0 146188 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_1589
timestamp 1666464484
transform 1 0 147292 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1595
timestamp 1666464484
transform 1 0 147844 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_1597
timestamp 1666464484
transform 1 0 148028 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1666464484
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1666464484
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1666464484
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1666464484
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1666464484
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1666464484
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1666464484
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1666464484
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1666464484
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1666464484
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1666464484
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1666464484
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1666464484
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1666464484
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1666464484
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1666464484
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1666464484
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1666464484
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1666464484
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1666464484
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1666464484
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1666464484
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1666464484
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1666464484
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1666464484
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1666464484
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1666464484
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1666464484
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1666464484
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1666464484
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1666464484
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1666464484
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1666464484
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1666464484
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1666464484
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1666464484
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1666464484
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1666464484
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1666464484
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1666464484
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1666464484
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1666464484
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1666464484
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1666464484
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1666464484
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1666464484
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1666464484
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1666464484
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1666464484
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1666464484
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1666464484
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1666464484
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1666464484
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1666464484
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1666464484
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1666464484
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1666464484
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1666464484
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1666464484
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1666464484
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1666464484
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1666464484
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1666464484
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_597
timestamp 1666464484
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1666464484
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1666464484
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_617
timestamp 1666464484
transform 1 0 57868 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_629
timestamp 1666464484
transform 1 0 58972 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_641
timestamp 1666464484
transform 1 0 60076 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_653
timestamp 1666464484
transform 1 0 61180 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_665
timestamp 1666464484
transform 1 0 62284 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_671
timestamp 1666464484
transform 1 0 62836 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_673
timestamp 1666464484
transform 1 0 63020 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_685
timestamp 1666464484
transform 1 0 64124 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_697
timestamp 1666464484
transform 1 0 65228 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_709
timestamp 1666464484
transform 1 0 66332 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_721
timestamp 1666464484
transform 1 0 67436 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_727
timestamp 1666464484
transform 1 0 67988 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_729
timestamp 1666464484
transform 1 0 68172 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_741
timestamp 1666464484
transform 1 0 69276 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_753
timestamp 1666464484
transform 1 0 70380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_765
timestamp 1666464484
transform 1 0 71484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_777
timestamp 1666464484
transform 1 0 72588 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_783
timestamp 1666464484
transform 1 0 73140 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_785
timestamp 1666464484
transform 1 0 73324 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_797
timestamp 1666464484
transform 1 0 74428 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_809
timestamp 1666464484
transform 1 0 75532 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_821
timestamp 1666464484
transform 1 0 76636 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_833
timestamp 1666464484
transform 1 0 77740 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_839
timestamp 1666464484
transform 1 0 78292 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_841
timestamp 1666464484
transform 1 0 78476 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_853
timestamp 1666464484
transform 1 0 79580 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_865
timestamp 1666464484
transform 1 0 80684 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_877
timestamp 1666464484
transform 1 0 81788 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_889
timestamp 1666464484
transform 1 0 82892 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_895
timestamp 1666464484
transform 1 0 83444 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_897
timestamp 1666464484
transform 1 0 83628 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_909
timestamp 1666464484
transform 1 0 84732 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_921
timestamp 1666464484
transform 1 0 85836 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_933
timestamp 1666464484
transform 1 0 86940 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_945
timestamp 1666464484
transform 1 0 88044 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_951
timestamp 1666464484
transform 1 0 88596 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_953
timestamp 1666464484
transform 1 0 88780 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_965
timestamp 1666464484
transform 1 0 89884 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_977
timestamp 1666464484
transform 1 0 90988 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_989
timestamp 1666464484
transform 1 0 92092 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_1001
timestamp 1666464484
transform 1 0 93196 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1007
timestamp 1666464484
transform 1 0 93748 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1009
timestamp 1666464484
transform 1 0 93932 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1021
timestamp 1666464484
transform 1 0 95036 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1033
timestamp 1666464484
transform 1 0 96140 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1045
timestamp 1666464484
transform 1 0 97244 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_1057
timestamp 1666464484
transform 1 0 98348 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1063
timestamp 1666464484
transform 1 0 98900 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1065
timestamp 1666464484
transform 1 0 99084 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1077
timestamp 1666464484
transform 1 0 100188 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1089
timestamp 1666464484
transform 1 0 101292 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1101
timestamp 1666464484
transform 1 0 102396 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_1113
timestamp 1666464484
transform 1 0 103500 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1119
timestamp 1666464484
transform 1 0 104052 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1121
timestamp 1666464484
transform 1 0 104236 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1133
timestamp 1666464484
transform 1 0 105340 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1145
timestamp 1666464484
transform 1 0 106444 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1157
timestamp 1666464484
transform 1 0 107548 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_1169
timestamp 1666464484
transform 1 0 108652 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1175
timestamp 1666464484
transform 1 0 109204 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1177
timestamp 1666464484
transform 1 0 109388 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1189
timestamp 1666464484
transform 1 0 110492 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1201
timestamp 1666464484
transform 1 0 111596 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1213
timestamp 1666464484
transform 1 0 112700 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_1225
timestamp 1666464484
transform 1 0 113804 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1231
timestamp 1666464484
transform 1 0 114356 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1233
timestamp 1666464484
transform 1 0 114540 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1245
timestamp 1666464484
transform 1 0 115644 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1257
timestamp 1666464484
transform 1 0 116748 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1269
timestamp 1666464484
transform 1 0 117852 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_1281
timestamp 1666464484
transform 1 0 118956 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1287
timestamp 1666464484
transform 1 0 119508 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1289
timestamp 1666464484
transform 1 0 119692 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1301
timestamp 1666464484
transform 1 0 120796 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1313
timestamp 1666464484
transform 1 0 121900 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1325
timestamp 1666464484
transform 1 0 123004 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_1337
timestamp 1666464484
transform 1 0 124108 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1343
timestamp 1666464484
transform 1 0 124660 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1345
timestamp 1666464484
transform 1 0 124844 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1357
timestamp 1666464484
transform 1 0 125948 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1369
timestamp 1666464484
transform 1 0 127052 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1381
timestamp 1666464484
transform 1 0 128156 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_1393
timestamp 1666464484
transform 1 0 129260 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1399
timestamp 1666464484
transform 1 0 129812 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1401
timestamp 1666464484
transform 1 0 129996 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1413
timestamp 1666464484
transform 1 0 131100 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1425
timestamp 1666464484
transform 1 0 132204 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1437
timestamp 1666464484
transform 1 0 133308 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_1449
timestamp 1666464484
transform 1 0 134412 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1455
timestamp 1666464484
transform 1 0 134964 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1457
timestamp 1666464484
transform 1 0 135148 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1469
timestamp 1666464484
transform 1 0 136252 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1481
timestamp 1666464484
transform 1 0 137356 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1493
timestamp 1666464484
transform 1 0 138460 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_1505
timestamp 1666464484
transform 1 0 139564 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1511
timestamp 1666464484
transform 1 0 140116 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1513
timestamp 1666464484
transform 1 0 140300 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1525
timestamp 1666464484
transform 1 0 141404 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1537
timestamp 1666464484
transform 1 0 142508 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1549
timestamp 1666464484
transform 1 0 143612 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_1561
timestamp 1666464484
transform 1 0 144716 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1567
timestamp 1666464484
transform 1 0 145268 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1569
timestamp 1666464484
transform 1 0 145452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1581
timestamp 1666464484
transform 1 0 146556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_1593
timestamp 1666464484
transform 1 0 147660 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_1601
timestamp 1666464484
transform 1 0 148396 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1666464484
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1666464484
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1666464484
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1666464484
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1666464484
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1666464484
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1666464484
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1666464484
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1666464484
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1666464484
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1666464484
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1666464484
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1666464484
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1666464484
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1666464484
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1666464484
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1666464484
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1666464484
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1666464484
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1666464484
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1666464484
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1666464484
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1666464484
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1666464484
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1666464484
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1666464484
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1666464484
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1666464484
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1666464484
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1666464484
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1666464484
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1666464484
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1666464484
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1666464484
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1666464484
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1666464484
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1666464484
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1666464484
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1666464484
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1666464484
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1666464484
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1666464484
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1666464484
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1666464484
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1666464484
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1666464484
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1666464484
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1666464484
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1666464484
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1666464484
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1666464484
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1666464484
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1666464484
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1666464484
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1666464484
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1666464484
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1666464484
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1666464484
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1666464484
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1666464484
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1666464484
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1666464484
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1666464484
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1666464484
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_601
timestamp 1666464484
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_613
timestamp 1666464484
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_625
timestamp 1666464484
transform 1 0 58604 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_637
timestamp 1666464484
transform 1 0 59708 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_643
timestamp 1666464484
transform 1 0 60260 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_645
timestamp 1666464484
transform 1 0 60444 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_657
timestamp 1666464484
transform 1 0 61548 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_669
timestamp 1666464484
transform 1 0 62652 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_681
timestamp 1666464484
transform 1 0 63756 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_693
timestamp 1666464484
transform 1 0 64860 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_699
timestamp 1666464484
transform 1 0 65412 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_701
timestamp 1666464484
transform 1 0 65596 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_713
timestamp 1666464484
transform 1 0 66700 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_725
timestamp 1666464484
transform 1 0 67804 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_737
timestamp 1666464484
transform 1 0 68908 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_749
timestamp 1666464484
transform 1 0 70012 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_755
timestamp 1666464484
transform 1 0 70564 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_757
timestamp 1666464484
transform 1 0 70748 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_769
timestamp 1666464484
transform 1 0 71852 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_781
timestamp 1666464484
transform 1 0 72956 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_793
timestamp 1666464484
transform 1 0 74060 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_805
timestamp 1666464484
transform 1 0 75164 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_811
timestamp 1666464484
transform 1 0 75716 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_813
timestamp 1666464484
transform 1 0 75900 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_825
timestamp 1666464484
transform 1 0 77004 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_837
timestamp 1666464484
transform 1 0 78108 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_849
timestamp 1666464484
transform 1 0 79212 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_861
timestamp 1666464484
transform 1 0 80316 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_867
timestamp 1666464484
transform 1 0 80868 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_869
timestamp 1666464484
transform 1 0 81052 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_881
timestamp 1666464484
transform 1 0 82156 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_893
timestamp 1666464484
transform 1 0 83260 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_905
timestamp 1666464484
transform 1 0 84364 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_917
timestamp 1666464484
transform 1 0 85468 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_923
timestamp 1666464484
transform 1 0 86020 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_925
timestamp 1666464484
transform 1 0 86204 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_937
timestamp 1666464484
transform 1 0 87308 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_949
timestamp 1666464484
transform 1 0 88412 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_961
timestamp 1666464484
transform 1 0 89516 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_973
timestamp 1666464484
transform 1 0 90620 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_979
timestamp 1666464484
transform 1 0 91172 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_981
timestamp 1666464484
transform 1 0 91356 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_993
timestamp 1666464484
transform 1 0 92460 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1005
timestamp 1666464484
transform 1 0 93564 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1017
timestamp 1666464484
transform 1 0 94668 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_1029
timestamp 1666464484
transform 1 0 95772 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1035
timestamp 1666464484
transform 1 0 96324 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1037
timestamp 1666464484
transform 1 0 96508 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1049
timestamp 1666464484
transform 1 0 97612 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1061
timestamp 1666464484
transform 1 0 98716 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1073
timestamp 1666464484
transform 1 0 99820 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_1085
timestamp 1666464484
transform 1 0 100924 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1091
timestamp 1666464484
transform 1 0 101476 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1093
timestamp 1666464484
transform 1 0 101660 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1105
timestamp 1666464484
transform 1 0 102764 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1117
timestamp 1666464484
transform 1 0 103868 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1129
timestamp 1666464484
transform 1 0 104972 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_1141
timestamp 1666464484
transform 1 0 106076 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1147
timestamp 1666464484
transform 1 0 106628 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1149
timestamp 1666464484
transform 1 0 106812 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1161
timestamp 1666464484
transform 1 0 107916 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1173
timestamp 1666464484
transform 1 0 109020 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1185
timestamp 1666464484
transform 1 0 110124 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_1197
timestamp 1666464484
transform 1 0 111228 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1203
timestamp 1666464484
transform 1 0 111780 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1205
timestamp 1666464484
transform 1 0 111964 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1217
timestamp 1666464484
transform 1 0 113068 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1229
timestamp 1666464484
transform 1 0 114172 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1241
timestamp 1666464484
transform 1 0 115276 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_1253
timestamp 1666464484
transform 1 0 116380 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1259
timestamp 1666464484
transform 1 0 116932 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1261
timestamp 1666464484
transform 1 0 117116 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1273
timestamp 1666464484
transform 1 0 118220 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1285
timestamp 1666464484
transform 1 0 119324 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1297
timestamp 1666464484
transform 1 0 120428 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_1309
timestamp 1666464484
transform 1 0 121532 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1315
timestamp 1666464484
transform 1 0 122084 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1317
timestamp 1666464484
transform 1 0 122268 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1329
timestamp 1666464484
transform 1 0 123372 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1341
timestamp 1666464484
transform 1 0 124476 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1353
timestamp 1666464484
transform 1 0 125580 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_1365
timestamp 1666464484
transform 1 0 126684 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1371
timestamp 1666464484
transform 1 0 127236 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1373
timestamp 1666464484
transform 1 0 127420 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1385
timestamp 1666464484
transform 1 0 128524 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1397
timestamp 1666464484
transform 1 0 129628 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1409
timestamp 1666464484
transform 1 0 130732 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_1421
timestamp 1666464484
transform 1 0 131836 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1427
timestamp 1666464484
transform 1 0 132388 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1429
timestamp 1666464484
transform 1 0 132572 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1441
timestamp 1666464484
transform 1 0 133676 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1453
timestamp 1666464484
transform 1 0 134780 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1465
timestamp 1666464484
transform 1 0 135884 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_1477
timestamp 1666464484
transform 1 0 136988 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1483
timestamp 1666464484
transform 1 0 137540 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1485
timestamp 1666464484
transform 1 0 137724 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1497
timestamp 1666464484
transform 1 0 138828 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1509
timestamp 1666464484
transform 1 0 139932 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1521
timestamp 1666464484
transform 1 0 141036 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_1533
timestamp 1666464484
transform 1 0 142140 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1539
timestamp 1666464484
transform 1 0 142692 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1541
timestamp 1666464484
transform 1 0 142876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1553
timestamp 1666464484
transform 1 0 143980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1565
timestamp 1666464484
transform 1 0 145084 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1577
timestamp 1666464484
transform 1 0 146188 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_1589
timestamp 1666464484
transform 1 0 147292 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1595
timestamp 1666464484
transform 1 0 147844 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_1597
timestamp 1666464484
transform 1 0 148028 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1666464484
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1666464484
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1666464484
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1666464484
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1666464484
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1666464484
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1666464484
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1666464484
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1666464484
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1666464484
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1666464484
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1666464484
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1666464484
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1666464484
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1666464484
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1666464484
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1666464484
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1666464484
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1666464484
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1666464484
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1666464484
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1666464484
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1666464484
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1666464484
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1666464484
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1666464484
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1666464484
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1666464484
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1666464484
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1666464484
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1666464484
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1666464484
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1666464484
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1666464484
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1666464484
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1666464484
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1666464484
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1666464484
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1666464484
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1666464484
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1666464484
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1666464484
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1666464484
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1666464484
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1666464484
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1666464484
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1666464484
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1666464484
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1666464484
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1666464484
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1666464484
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1666464484
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1666464484
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1666464484
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1666464484
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1666464484
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1666464484
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1666464484
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1666464484
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1666464484
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1666464484
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1666464484
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1666464484
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_597
timestamp 1666464484
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1666464484
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1666464484
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_617
timestamp 1666464484
transform 1 0 57868 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_629
timestamp 1666464484
transform 1 0 58972 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_641
timestamp 1666464484
transform 1 0 60076 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_653
timestamp 1666464484
transform 1 0 61180 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_665
timestamp 1666464484
transform 1 0 62284 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_671
timestamp 1666464484
transform 1 0 62836 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_673
timestamp 1666464484
transform 1 0 63020 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_685
timestamp 1666464484
transform 1 0 64124 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_697
timestamp 1666464484
transform 1 0 65228 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_709
timestamp 1666464484
transform 1 0 66332 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_721
timestamp 1666464484
transform 1 0 67436 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_727
timestamp 1666464484
transform 1 0 67988 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_729
timestamp 1666464484
transform 1 0 68172 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_741
timestamp 1666464484
transform 1 0 69276 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_753
timestamp 1666464484
transform 1 0 70380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_765
timestamp 1666464484
transform 1 0 71484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_777
timestamp 1666464484
transform 1 0 72588 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_783
timestamp 1666464484
transform 1 0 73140 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_785
timestamp 1666464484
transform 1 0 73324 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_797
timestamp 1666464484
transform 1 0 74428 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_809
timestamp 1666464484
transform 1 0 75532 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_821
timestamp 1666464484
transform 1 0 76636 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_833
timestamp 1666464484
transform 1 0 77740 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_839
timestamp 1666464484
transform 1 0 78292 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_841
timestamp 1666464484
transform 1 0 78476 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_853
timestamp 1666464484
transform 1 0 79580 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_865
timestamp 1666464484
transform 1 0 80684 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_877
timestamp 1666464484
transform 1 0 81788 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_889
timestamp 1666464484
transform 1 0 82892 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_895
timestamp 1666464484
transform 1 0 83444 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_897
timestamp 1666464484
transform 1 0 83628 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_909
timestamp 1666464484
transform 1 0 84732 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_921
timestamp 1666464484
transform 1 0 85836 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_933
timestamp 1666464484
transform 1 0 86940 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_945
timestamp 1666464484
transform 1 0 88044 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_951
timestamp 1666464484
transform 1 0 88596 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_953
timestamp 1666464484
transform 1 0 88780 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_965
timestamp 1666464484
transform 1 0 89884 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_977
timestamp 1666464484
transform 1 0 90988 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_989
timestamp 1666464484
transform 1 0 92092 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_1001
timestamp 1666464484
transform 1 0 93196 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_1007
timestamp 1666464484
transform 1 0 93748 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1009
timestamp 1666464484
transform 1 0 93932 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1021
timestamp 1666464484
transform 1 0 95036 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1033
timestamp 1666464484
transform 1 0 96140 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1045
timestamp 1666464484
transform 1 0 97244 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_1057
timestamp 1666464484
transform 1 0 98348 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_1063
timestamp 1666464484
transform 1 0 98900 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1065
timestamp 1666464484
transform 1 0 99084 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1077
timestamp 1666464484
transform 1 0 100188 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1089
timestamp 1666464484
transform 1 0 101292 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1101
timestamp 1666464484
transform 1 0 102396 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_1113
timestamp 1666464484
transform 1 0 103500 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_1119
timestamp 1666464484
transform 1 0 104052 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1121
timestamp 1666464484
transform 1 0 104236 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1133
timestamp 1666464484
transform 1 0 105340 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1145
timestamp 1666464484
transform 1 0 106444 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1157
timestamp 1666464484
transform 1 0 107548 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_1169
timestamp 1666464484
transform 1 0 108652 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_1175
timestamp 1666464484
transform 1 0 109204 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1177
timestamp 1666464484
transform 1 0 109388 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1189
timestamp 1666464484
transform 1 0 110492 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1201
timestamp 1666464484
transform 1 0 111596 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1213
timestamp 1666464484
transform 1 0 112700 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_1225
timestamp 1666464484
transform 1 0 113804 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_1231
timestamp 1666464484
transform 1 0 114356 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1233
timestamp 1666464484
transform 1 0 114540 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1245
timestamp 1666464484
transform 1 0 115644 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1257
timestamp 1666464484
transform 1 0 116748 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1269
timestamp 1666464484
transform 1 0 117852 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_1281
timestamp 1666464484
transform 1 0 118956 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_1287
timestamp 1666464484
transform 1 0 119508 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1289
timestamp 1666464484
transform 1 0 119692 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1301
timestamp 1666464484
transform 1 0 120796 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1313
timestamp 1666464484
transform 1 0 121900 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1325
timestamp 1666464484
transform 1 0 123004 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_1337
timestamp 1666464484
transform 1 0 124108 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_1343
timestamp 1666464484
transform 1 0 124660 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1345
timestamp 1666464484
transform 1 0 124844 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1357
timestamp 1666464484
transform 1 0 125948 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1369
timestamp 1666464484
transform 1 0 127052 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1381
timestamp 1666464484
transform 1 0 128156 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_1393
timestamp 1666464484
transform 1 0 129260 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_1399
timestamp 1666464484
transform 1 0 129812 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1401
timestamp 1666464484
transform 1 0 129996 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1413
timestamp 1666464484
transform 1 0 131100 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1425
timestamp 1666464484
transform 1 0 132204 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1437
timestamp 1666464484
transform 1 0 133308 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_1449
timestamp 1666464484
transform 1 0 134412 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_1455
timestamp 1666464484
transform 1 0 134964 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1457
timestamp 1666464484
transform 1 0 135148 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1469
timestamp 1666464484
transform 1 0 136252 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1481
timestamp 1666464484
transform 1 0 137356 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1493
timestamp 1666464484
transform 1 0 138460 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_1505
timestamp 1666464484
transform 1 0 139564 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_1511
timestamp 1666464484
transform 1 0 140116 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1513
timestamp 1666464484
transform 1 0 140300 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1525
timestamp 1666464484
transform 1 0 141404 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1537
timestamp 1666464484
transform 1 0 142508 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1549
timestamp 1666464484
transform 1 0 143612 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_1561
timestamp 1666464484
transform 1 0 144716 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_1567
timestamp 1666464484
transform 1 0 145268 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1569
timestamp 1666464484
transform 1 0 145452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1581
timestamp 1666464484
transform 1 0 146556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_1593
timestamp 1666464484
transform 1 0 147660 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_1601
timestamp 1666464484
transform 1 0 148396 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1666464484
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1666464484
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1666464484
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1666464484
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1666464484
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1666464484
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1666464484
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1666464484
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1666464484
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1666464484
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1666464484
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1666464484
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1666464484
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1666464484
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1666464484
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1666464484
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1666464484
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1666464484
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1666464484
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1666464484
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1666464484
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1666464484
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1666464484
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1666464484
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1666464484
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1666464484
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1666464484
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1666464484
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1666464484
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1666464484
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1666464484
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1666464484
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1666464484
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1666464484
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1666464484
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1666464484
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1666464484
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1666464484
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1666464484
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1666464484
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1666464484
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1666464484
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1666464484
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1666464484
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1666464484
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1666464484
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1666464484
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1666464484
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1666464484
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1666464484
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1666464484
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1666464484
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1666464484
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1666464484
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1666464484
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1666464484
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1666464484
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1666464484
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1666464484
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1666464484
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1666464484
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1666464484
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1666464484
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1666464484
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1666464484
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_613
timestamp 1666464484
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_625
timestamp 1666464484
transform 1 0 58604 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_637
timestamp 1666464484
transform 1 0 59708 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_643
timestamp 1666464484
transform 1 0 60260 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_645
timestamp 1666464484
transform 1 0 60444 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_657
timestamp 1666464484
transform 1 0 61548 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_669
timestamp 1666464484
transform 1 0 62652 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_681
timestamp 1666464484
transform 1 0 63756 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_693
timestamp 1666464484
transform 1 0 64860 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_699
timestamp 1666464484
transform 1 0 65412 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_701
timestamp 1666464484
transform 1 0 65596 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_713
timestamp 1666464484
transform 1 0 66700 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_725
timestamp 1666464484
transform 1 0 67804 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_737
timestamp 1666464484
transform 1 0 68908 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_749
timestamp 1666464484
transform 1 0 70012 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_755
timestamp 1666464484
transform 1 0 70564 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_757
timestamp 1666464484
transform 1 0 70748 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_769
timestamp 1666464484
transform 1 0 71852 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_781
timestamp 1666464484
transform 1 0 72956 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_793
timestamp 1666464484
transform 1 0 74060 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_805
timestamp 1666464484
transform 1 0 75164 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_811
timestamp 1666464484
transform 1 0 75716 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_813
timestamp 1666464484
transform 1 0 75900 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_825
timestamp 1666464484
transform 1 0 77004 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_837
timestamp 1666464484
transform 1 0 78108 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_849
timestamp 1666464484
transform 1 0 79212 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_861
timestamp 1666464484
transform 1 0 80316 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_867
timestamp 1666464484
transform 1 0 80868 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_869
timestamp 1666464484
transform 1 0 81052 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_881
timestamp 1666464484
transform 1 0 82156 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_893
timestamp 1666464484
transform 1 0 83260 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_905
timestamp 1666464484
transform 1 0 84364 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_917
timestamp 1666464484
transform 1 0 85468 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_923
timestamp 1666464484
transform 1 0 86020 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_925
timestamp 1666464484
transform 1 0 86204 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_937
timestamp 1666464484
transform 1 0 87308 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_949
timestamp 1666464484
transform 1 0 88412 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_961
timestamp 1666464484
transform 1 0 89516 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_973
timestamp 1666464484
transform 1 0 90620 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_979
timestamp 1666464484
transform 1 0 91172 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_981
timestamp 1666464484
transform 1 0 91356 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_993
timestamp 1666464484
transform 1 0 92460 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1005
timestamp 1666464484
transform 1 0 93564 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1017
timestamp 1666464484
transform 1 0 94668 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_1029
timestamp 1666464484
transform 1 0 95772 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1035
timestamp 1666464484
transform 1 0 96324 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1037
timestamp 1666464484
transform 1 0 96508 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1049
timestamp 1666464484
transform 1 0 97612 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1061
timestamp 1666464484
transform 1 0 98716 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1073
timestamp 1666464484
transform 1 0 99820 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_1085
timestamp 1666464484
transform 1 0 100924 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1091
timestamp 1666464484
transform 1 0 101476 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1093
timestamp 1666464484
transform 1 0 101660 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1105
timestamp 1666464484
transform 1 0 102764 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1117
timestamp 1666464484
transform 1 0 103868 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1129
timestamp 1666464484
transform 1 0 104972 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_1141
timestamp 1666464484
transform 1 0 106076 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1147
timestamp 1666464484
transform 1 0 106628 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1149
timestamp 1666464484
transform 1 0 106812 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1161
timestamp 1666464484
transform 1 0 107916 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1173
timestamp 1666464484
transform 1 0 109020 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1185
timestamp 1666464484
transform 1 0 110124 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_1197
timestamp 1666464484
transform 1 0 111228 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1203
timestamp 1666464484
transform 1 0 111780 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1205
timestamp 1666464484
transform 1 0 111964 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1217
timestamp 1666464484
transform 1 0 113068 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1229
timestamp 1666464484
transform 1 0 114172 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1241
timestamp 1666464484
transform 1 0 115276 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_1253
timestamp 1666464484
transform 1 0 116380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1259
timestamp 1666464484
transform 1 0 116932 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1261
timestamp 1666464484
transform 1 0 117116 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1273
timestamp 1666464484
transform 1 0 118220 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1285
timestamp 1666464484
transform 1 0 119324 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1297
timestamp 1666464484
transform 1 0 120428 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_1309
timestamp 1666464484
transform 1 0 121532 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1315
timestamp 1666464484
transform 1 0 122084 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1317
timestamp 1666464484
transform 1 0 122268 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1329
timestamp 1666464484
transform 1 0 123372 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1341
timestamp 1666464484
transform 1 0 124476 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1353
timestamp 1666464484
transform 1 0 125580 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_1365
timestamp 1666464484
transform 1 0 126684 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1371
timestamp 1666464484
transform 1 0 127236 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1373
timestamp 1666464484
transform 1 0 127420 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1385
timestamp 1666464484
transform 1 0 128524 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1397
timestamp 1666464484
transform 1 0 129628 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1409
timestamp 1666464484
transform 1 0 130732 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_1421
timestamp 1666464484
transform 1 0 131836 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1427
timestamp 1666464484
transform 1 0 132388 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1429
timestamp 1666464484
transform 1 0 132572 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1441
timestamp 1666464484
transform 1 0 133676 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1453
timestamp 1666464484
transform 1 0 134780 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1465
timestamp 1666464484
transform 1 0 135884 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_1477
timestamp 1666464484
transform 1 0 136988 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1483
timestamp 1666464484
transform 1 0 137540 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1485
timestamp 1666464484
transform 1 0 137724 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1497
timestamp 1666464484
transform 1 0 138828 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1509
timestamp 1666464484
transform 1 0 139932 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1521
timestamp 1666464484
transform 1 0 141036 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_1533
timestamp 1666464484
transform 1 0 142140 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1539
timestamp 1666464484
transform 1 0 142692 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1541
timestamp 1666464484
transform 1 0 142876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1553
timestamp 1666464484
transform 1 0 143980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1565
timestamp 1666464484
transform 1 0 145084 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1577
timestamp 1666464484
transform 1 0 146188 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_1589
timestamp 1666464484
transform 1 0 147292 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1595
timestamp 1666464484
transform 1 0 147844 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_1597
timestamp 1666464484
transform 1 0 148028 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1666464484
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1666464484
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1666464484
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1666464484
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1666464484
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1666464484
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1666464484
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1666464484
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1666464484
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1666464484
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1666464484
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1666464484
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1666464484
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1666464484
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1666464484
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1666464484
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1666464484
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1666464484
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1666464484
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1666464484
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1666464484
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1666464484
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1666464484
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1666464484
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1666464484
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1666464484
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1666464484
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1666464484
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1666464484
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1666464484
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1666464484
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1666464484
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1666464484
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1666464484
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1666464484
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1666464484
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1666464484
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1666464484
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1666464484
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1666464484
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1666464484
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1666464484
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1666464484
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1666464484
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1666464484
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1666464484
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1666464484
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1666464484
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1666464484
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1666464484
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1666464484
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1666464484
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1666464484
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1666464484
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1666464484
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1666464484
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1666464484
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1666464484
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1666464484
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1666464484
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1666464484
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1666464484
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1666464484
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_597
timestamp 1666464484
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1666464484
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1666464484
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_617
timestamp 1666464484
transform 1 0 57868 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_629
timestamp 1666464484
transform 1 0 58972 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_641
timestamp 1666464484
transform 1 0 60076 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_653
timestamp 1666464484
transform 1 0 61180 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_665
timestamp 1666464484
transform 1 0 62284 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_671
timestamp 1666464484
transform 1 0 62836 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_673
timestamp 1666464484
transform 1 0 63020 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_685
timestamp 1666464484
transform 1 0 64124 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_697
timestamp 1666464484
transform 1 0 65228 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_709
timestamp 1666464484
transform 1 0 66332 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_721
timestamp 1666464484
transform 1 0 67436 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_727
timestamp 1666464484
transform 1 0 67988 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_729
timestamp 1666464484
transform 1 0 68172 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_741
timestamp 1666464484
transform 1 0 69276 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_753
timestamp 1666464484
transform 1 0 70380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_765
timestamp 1666464484
transform 1 0 71484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_777
timestamp 1666464484
transform 1 0 72588 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_783
timestamp 1666464484
transform 1 0 73140 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_785
timestamp 1666464484
transform 1 0 73324 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_797
timestamp 1666464484
transform 1 0 74428 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_809
timestamp 1666464484
transform 1 0 75532 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_821
timestamp 1666464484
transform 1 0 76636 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_833
timestamp 1666464484
transform 1 0 77740 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_839
timestamp 1666464484
transform 1 0 78292 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_841
timestamp 1666464484
transform 1 0 78476 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_853
timestamp 1666464484
transform 1 0 79580 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_865
timestamp 1666464484
transform 1 0 80684 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_877
timestamp 1666464484
transform 1 0 81788 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_889
timestamp 1666464484
transform 1 0 82892 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_895
timestamp 1666464484
transform 1 0 83444 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_897
timestamp 1666464484
transform 1 0 83628 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_909
timestamp 1666464484
transform 1 0 84732 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_921
timestamp 1666464484
transform 1 0 85836 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_933
timestamp 1666464484
transform 1 0 86940 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_945
timestamp 1666464484
transform 1 0 88044 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_951
timestamp 1666464484
transform 1 0 88596 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_953
timestamp 1666464484
transform 1 0 88780 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_965
timestamp 1666464484
transform 1 0 89884 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_977
timestamp 1666464484
transform 1 0 90988 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_989
timestamp 1666464484
transform 1 0 92092 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_1001
timestamp 1666464484
transform 1 0 93196 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_1007
timestamp 1666464484
transform 1 0 93748 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1009
timestamp 1666464484
transform 1 0 93932 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1021
timestamp 1666464484
transform 1 0 95036 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1033
timestamp 1666464484
transform 1 0 96140 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1045
timestamp 1666464484
transform 1 0 97244 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_1057
timestamp 1666464484
transform 1 0 98348 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_1063
timestamp 1666464484
transform 1 0 98900 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1065
timestamp 1666464484
transform 1 0 99084 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1077
timestamp 1666464484
transform 1 0 100188 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1089
timestamp 1666464484
transform 1 0 101292 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1101
timestamp 1666464484
transform 1 0 102396 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_1113
timestamp 1666464484
transform 1 0 103500 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_1119
timestamp 1666464484
transform 1 0 104052 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1121
timestamp 1666464484
transform 1 0 104236 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1133
timestamp 1666464484
transform 1 0 105340 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1145
timestamp 1666464484
transform 1 0 106444 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1157
timestamp 1666464484
transform 1 0 107548 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_1169
timestamp 1666464484
transform 1 0 108652 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_1175
timestamp 1666464484
transform 1 0 109204 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1177
timestamp 1666464484
transform 1 0 109388 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1189
timestamp 1666464484
transform 1 0 110492 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1201
timestamp 1666464484
transform 1 0 111596 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1213
timestamp 1666464484
transform 1 0 112700 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_1225
timestamp 1666464484
transform 1 0 113804 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_1231
timestamp 1666464484
transform 1 0 114356 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1233
timestamp 1666464484
transform 1 0 114540 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1245
timestamp 1666464484
transform 1 0 115644 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1257
timestamp 1666464484
transform 1 0 116748 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1269
timestamp 1666464484
transform 1 0 117852 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_1281
timestamp 1666464484
transform 1 0 118956 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_1287
timestamp 1666464484
transform 1 0 119508 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1289
timestamp 1666464484
transform 1 0 119692 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1301
timestamp 1666464484
transform 1 0 120796 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1313
timestamp 1666464484
transform 1 0 121900 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1325
timestamp 1666464484
transform 1 0 123004 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_1337
timestamp 1666464484
transform 1 0 124108 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_1343
timestamp 1666464484
transform 1 0 124660 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1345
timestamp 1666464484
transform 1 0 124844 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1357
timestamp 1666464484
transform 1 0 125948 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1369
timestamp 1666464484
transform 1 0 127052 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1381
timestamp 1666464484
transform 1 0 128156 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_1393
timestamp 1666464484
transform 1 0 129260 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_1399
timestamp 1666464484
transform 1 0 129812 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1401
timestamp 1666464484
transform 1 0 129996 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1413
timestamp 1666464484
transform 1 0 131100 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1425
timestamp 1666464484
transform 1 0 132204 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1437
timestamp 1666464484
transform 1 0 133308 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_1449
timestamp 1666464484
transform 1 0 134412 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_1455
timestamp 1666464484
transform 1 0 134964 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1457
timestamp 1666464484
transform 1 0 135148 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1469
timestamp 1666464484
transform 1 0 136252 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1481
timestamp 1666464484
transform 1 0 137356 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1493
timestamp 1666464484
transform 1 0 138460 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_1505
timestamp 1666464484
transform 1 0 139564 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_1511
timestamp 1666464484
transform 1 0 140116 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1513
timestamp 1666464484
transform 1 0 140300 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1525
timestamp 1666464484
transform 1 0 141404 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1537
timestamp 1666464484
transform 1 0 142508 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1549
timestamp 1666464484
transform 1 0 143612 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_1561
timestamp 1666464484
transform 1 0 144716 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_1567
timestamp 1666464484
transform 1 0 145268 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1569
timestamp 1666464484
transform 1 0 145452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1581
timestamp 1666464484
transform 1 0 146556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_1593
timestamp 1666464484
transform 1 0 147660 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_1601
timestamp 1666464484
transform 1 0 148396 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1666464484
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1666464484
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1666464484
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1666464484
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1666464484
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1666464484
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1666464484
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1666464484
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1666464484
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1666464484
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1666464484
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1666464484
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1666464484
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1666464484
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1666464484
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1666464484
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1666464484
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1666464484
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1666464484
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1666464484
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1666464484
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1666464484
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1666464484
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1666464484
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1666464484
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1666464484
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1666464484
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1666464484
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1666464484
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1666464484
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1666464484
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1666464484
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1666464484
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1666464484
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1666464484
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1666464484
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1666464484
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1666464484
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1666464484
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1666464484
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1666464484
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1666464484
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1666464484
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1666464484
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1666464484
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1666464484
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1666464484
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1666464484
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1666464484
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1666464484
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1666464484
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1666464484
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1666464484
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1666464484
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1666464484
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1666464484
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1666464484
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1666464484
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1666464484
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1666464484
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1666464484
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1666464484
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1666464484
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1666464484
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_601
timestamp 1666464484
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_613
timestamp 1666464484
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_625
timestamp 1666464484
transform 1 0 58604 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_637
timestamp 1666464484
transform 1 0 59708 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_643
timestamp 1666464484
transform 1 0 60260 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_645
timestamp 1666464484
transform 1 0 60444 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_657
timestamp 1666464484
transform 1 0 61548 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_669
timestamp 1666464484
transform 1 0 62652 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_681
timestamp 1666464484
transform 1 0 63756 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_693
timestamp 1666464484
transform 1 0 64860 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_699
timestamp 1666464484
transform 1 0 65412 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_701
timestamp 1666464484
transform 1 0 65596 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_713
timestamp 1666464484
transform 1 0 66700 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_725
timestamp 1666464484
transform 1 0 67804 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_737
timestamp 1666464484
transform 1 0 68908 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_749
timestamp 1666464484
transform 1 0 70012 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_755
timestamp 1666464484
transform 1 0 70564 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_757
timestamp 1666464484
transform 1 0 70748 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_769
timestamp 1666464484
transform 1 0 71852 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_781
timestamp 1666464484
transform 1 0 72956 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_793
timestamp 1666464484
transform 1 0 74060 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_805
timestamp 1666464484
transform 1 0 75164 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_811
timestamp 1666464484
transform 1 0 75716 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_813
timestamp 1666464484
transform 1 0 75900 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_825
timestamp 1666464484
transform 1 0 77004 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_837
timestamp 1666464484
transform 1 0 78108 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_849
timestamp 1666464484
transform 1 0 79212 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_861
timestamp 1666464484
transform 1 0 80316 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_867
timestamp 1666464484
transform 1 0 80868 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_869
timestamp 1666464484
transform 1 0 81052 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_881
timestamp 1666464484
transform 1 0 82156 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_893
timestamp 1666464484
transform 1 0 83260 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_905
timestamp 1666464484
transform 1 0 84364 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_917
timestamp 1666464484
transform 1 0 85468 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_923
timestamp 1666464484
transform 1 0 86020 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_925
timestamp 1666464484
transform 1 0 86204 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_937
timestamp 1666464484
transform 1 0 87308 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_949
timestamp 1666464484
transform 1 0 88412 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_961
timestamp 1666464484
transform 1 0 89516 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_973
timestamp 1666464484
transform 1 0 90620 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_979
timestamp 1666464484
transform 1 0 91172 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_981
timestamp 1666464484
transform 1 0 91356 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_993
timestamp 1666464484
transform 1 0 92460 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1005
timestamp 1666464484
transform 1 0 93564 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1017
timestamp 1666464484
transform 1 0 94668 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_1029
timestamp 1666464484
transform 1 0 95772 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1035
timestamp 1666464484
transform 1 0 96324 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1037
timestamp 1666464484
transform 1 0 96508 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1049
timestamp 1666464484
transform 1 0 97612 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1061
timestamp 1666464484
transform 1 0 98716 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1073
timestamp 1666464484
transform 1 0 99820 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_1085
timestamp 1666464484
transform 1 0 100924 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1091
timestamp 1666464484
transform 1 0 101476 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1093
timestamp 1666464484
transform 1 0 101660 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1105
timestamp 1666464484
transform 1 0 102764 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1117
timestamp 1666464484
transform 1 0 103868 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1129
timestamp 1666464484
transform 1 0 104972 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_1141
timestamp 1666464484
transform 1 0 106076 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1147
timestamp 1666464484
transform 1 0 106628 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1149
timestamp 1666464484
transform 1 0 106812 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1161
timestamp 1666464484
transform 1 0 107916 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1173
timestamp 1666464484
transform 1 0 109020 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1185
timestamp 1666464484
transform 1 0 110124 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_1197
timestamp 1666464484
transform 1 0 111228 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1203
timestamp 1666464484
transform 1 0 111780 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1205
timestamp 1666464484
transform 1 0 111964 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1217
timestamp 1666464484
transform 1 0 113068 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1229
timestamp 1666464484
transform 1 0 114172 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1241
timestamp 1666464484
transform 1 0 115276 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_1253
timestamp 1666464484
transform 1 0 116380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1259
timestamp 1666464484
transform 1 0 116932 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1261
timestamp 1666464484
transform 1 0 117116 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1273
timestamp 1666464484
transform 1 0 118220 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1285
timestamp 1666464484
transform 1 0 119324 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1297
timestamp 1666464484
transform 1 0 120428 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_1309
timestamp 1666464484
transform 1 0 121532 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1315
timestamp 1666464484
transform 1 0 122084 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1317
timestamp 1666464484
transform 1 0 122268 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1329
timestamp 1666464484
transform 1 0 123372 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1341
timestamp 1666464484
transform 1 0 124476 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1353
timestamp 1666464484
transform 1 0 125580 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_1365
timestamp 1666464484
transform 1 0 126684 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1371
timestamp 1666464484
transform 1 0 127236 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1373
timestamp 1666464484
transform 1 0 127420 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1385
timestamp 1666464484
transform 1 0 128524 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1397
timestamp 1666464484
transform 1 0 129628 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1409
timestamp 1666464484
transform 1 0 130732 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_1421
timestamp 1666464484
transform 1 0 131836 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1427
timestamp 1666464484
transform 1 0 132388 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1429
timestamp 1666464484
transform 1 0 132572 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1441
timestamp 1666464484
transform 1 0 133676 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1453
timestamp 1666464484
transform 1 0 134780 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1465
timestamp 1666464484
transform 1 0 135884 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_1477
timestamp 1666464484
transform 1 0 136988 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1483
timestamp 1666464484
transform 1 0 137540 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1485
timestamp 1666464484
transform 1 0 137724 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1497
timestamp 1666464484
transform 1 0 138828 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1509
timestamp 1666464484
transform 1 0 139932 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1521
timestamp 1666464484
transform 1 0 141036 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_1533
timestamp 1666464484
transform 1 0 142140 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1539
timestamp 1666464484
transform 1 0 142692 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1541
timestamp 1666464484
transform 1 0 142876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1553
timestamp 1666464484
transform 1 0 143980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1565
timestamp 1666464484
transform 1 0 145084 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1577
timestamp 1666464484
transform 1 0 146188 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_1589
timestamp 1666464484
transform 1 0 147292 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1595
timestamp 1666464484
transform 1 0 147844 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_1597
timestamp 1666464484
transform 1 0 148028 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1666464484
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1666464484
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1666464484
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1666464484
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1666464484
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1666464484
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1666464484
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1666464484
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1666464484
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1666464484
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1666464484
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1666464484
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1666464484
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1666464484
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1666464484
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1666464484
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1666464484
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1666464484
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1666464484
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1666464484
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1666464484
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1666464484
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1666464484
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1666464484
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1666464484
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1666464484
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1666464484
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1666464484
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1666464484
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1666464484
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1666464484
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1666464484
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1666464484
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1666464484
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1666464484
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1666464484
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1666464484
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1666464484
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1666464484
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1666464484
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1666464484
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1666464484
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1666464484
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1666464484
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1666464484
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1666464484
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1666464484
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1666464484
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1666464484
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1666464484
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1666464484
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1666464484
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1666464484
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1666464484
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1666464484
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1666464484
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1666464484
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1666464484
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1666464484
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1666464484
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1666464484
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1666464484
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1666464484
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_597
timestamp 1666464484
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1666464484
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1666464484
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_617
timestamp 1666464484
transform 1 0 57868 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_629
timestamp 1666464484
transform 1 0 58972 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_641
timestamp 1666464484
transform 1 0 60076 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_653
timestamp 1666464484
transform 1 0 61180 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_665
timestamp 1666464484
transform 1 0 62284 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_671
timestamp 1666464484
transform 1 0 62836 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_673
timestamp 1666464484
transform 1 0 63020 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_685
timestamp 1666464484
transform 1 0 64124 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_697
timestamp 1666464484
transform 1 0 65228 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_709
timestamp 1666464484
transform 1 0 66332 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_721
timestamp 1666464484
transform 1 0 67436 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_727
timestamp 1666464484
transform 1 0 67988 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_729
timestamp 1666464484
transform 1 0 68172 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_741
timestamp 1666464484
transform 1 0 69276 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_753
timestamp 1666464484
transform 1 0 70380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_765
timestamp 1666464484
transform 1 0 71484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_777
timestamp 1666464484
transform 1 0 72588 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_783
timestamp 1666464484
transform 1 0 73140 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_785
timestamp 1666464484
transform 1 0 73324 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_797
timestamp 1666464484
transform 1 0 74428 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_809
timestamp 1666464484
transform 1 0 75532 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_821
timestamp 1666464484
transform 1 0 76636 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_833
timestamp 1666464484
transform 1 0 77740 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_839
timestamp 1666464484
transform 1 0 78292 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_841
timestamp 1666464484
transform 1 0 78476 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_853
timestamp 1666464484
transform 1 0 79580 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_865
timestamp 1666464484
transform 1 0 80684 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_877
timestamp 1666464484
transform 1 0 81788 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_889
timestamp 1666464484
transform 1 0 82892 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_895
timestamp 1666464484
transform 1 0 83444 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_897
timestamp 1666464484
transform 1 0 83628 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_909
timestamp 1666464484
transform 1 0 84732 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_921
timestamp 1666464484
transform 1 0 85836 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_933
timestamp 1666464484
transform 1 0 86940 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_945
timestamp 1666464484
transform 1 0 88044 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_951
timestamp 1666464484
transform 1 0 88596 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_953
timestamp 1666464484
transform 1 0 88780 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_965
timestamp 1666464484
transform 1 0 89884 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_977
timestamp 1666464484
transform 1 0 90988 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_989
timestamp 1666464484
transform 1 0 92092 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_1001
timestamp 1666464484
transform 1 0 93196 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_1007
timestamp 1666464484
transform 1 0 93748 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1009
timestamp 1666464484
transform 1 0 93932 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1021
timestamp 1666464484
transform 1 0 95036 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1033
timestamp 1666464484
transform 1 0 96140 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1045
timestamp 1666464484
transform 1 0 97244 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_1057
timestamp 1666464484
transform 1 0 98348 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_1063
timestamp 1666464484
transform 1 0 98900 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1065
timestamp 1666464484
transform 1 0 99084 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1077
timestamp 1666464484
transform 1 0 100188 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1089
timestamp 1666464484
transform 1 0 101292 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1101
timestamp 1666464484
transform 1 0 102396 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_1113
timestamp 1666464484
transform 1 0 103500 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_1119
timestamp 1666464484
transform 1 0 104052 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1121
timestamp 1666464484
transform 1 0 104236 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1133
timestamp 1666464484
transform 1 0 105340 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1145
timestamp 1666464484
transform 1 0 106444 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1157
timestamp 1666464484
transform 1 0 107548 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_1169
timestamp 1666464484
transform 1 0 108652 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_1175
timestamp 1666464484
transform 1 0 109204 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1177
timestamp 1666464484
transform 1 0 109388 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1189
timestamp 1666464484
transform 1 0 110492 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1201
timestamp 1666464484
transform 1 0 111596 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1213
timestamp 1666464484
transform 1 0 112700 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_1225
timestamp 1666464484
transform 1 0 113804 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_1231
timestamp 1666464484
transform 1 0 114356 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1233
timestamp 1666464484
transform 1 0 114540 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1245
timestamp 1666464484
transform 1 0 115644 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1257
timestamp 1666464484
transform 1 0 116748 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1269
timestamp 1666464484
transform 1 0 117852 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_1281
timestamp 1666464484
transform 1 0 118956 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_1287
timestamp 1666464484
transform 1 0 119508 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1289
timestamp 1666464484
transform 1 0 119692 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1301
timestamp 1666464484
transform 1 0 120796 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1313
timestamp 1666464484
transform 1 0 121900 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1325
timestamp 1666464484
transform 1 0 123004 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_1337
timestamp 1666464484
transform 1 0 124108 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_1343
timestamp 1666464484
transform 1 0 124660 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1345
timestamp 1666464484
transform 1 0 124844 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1357
timestamp 1666464484
transform 1 0 125948 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1369
timestamp 1666464484
transform 1 0 127052 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1381
timestamp 1666464484
transform 1 0 128156 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_1393
timestamp 1666464484
transform 1 0 129260 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_1399
timestamp 1666464484
transform 1 0 129812 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1401
timestamp 1666464484
transform 1 0 129996 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1413
timestamp 1666464484
transform 1 0 131100 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1425
timestamp 1666464484
transform 1 0 132204 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1437
timestamp 1666464484
transform 1 0 133308 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_1449
timestamp 1666464484
transform 1 0 134412 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_1455
timestamp 1666464484
transform 1 0 134964 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1457
timestamp 1666464484
transform 1 0 135148 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1469
timestamp 1666464484
transform 1 0 136252 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1481
timestamp 1666464484
transform 1 0 137356 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1493
timestamp 1666464484
transform 1 0 138460 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_1505
timestamp 1666464484
transform 1 0 139564 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_1511
timestamp 1666464484
transform 1 0 140116 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1513
timestamp 1666464484
transform 1 0 140300 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1525
timestamp 1666464484
transform 1 0 141404 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1537
timestamp 1666464484
transform 1 0 142508 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1549
timestamp 1666464484
transform 1 0 143612 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_1561
timestamp 1666464484
transform 1 0 144716 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_1567
timestamp 1666464484
transform 1 0 145268 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1569
timestamp 1666464484
transform 1 0 145452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1581
timestamp 1666464484
transform 1 0 146556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_1593
timestamp 1666464484
transform 1 0 147660 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_1601
timestamp 1666464484
transform 1 0 148396 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1666464484
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1666464484
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1666464484
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1666464484
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1666464484
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1666464484
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1666464484
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1666464484
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1666464484
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1666464484
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1666464484
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1666464484
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1666464484
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1666464484
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1666464484
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1666464484
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1666464484
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1666464484
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1666464484
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1666464484
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1666464484
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1666464484
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1666464484
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1666464484
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1666464484
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1666464484
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1666464484
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1666464484
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1666464484
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1666464484
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1666464484
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1666464484
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1666464484
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1666464484
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1666464484
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1666464484
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1666464484
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1666464484
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1666464484
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1666464484
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1666464484
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1666464484
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1666464484
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1666464484
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1666464484
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1666464484
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1666464484
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1666464484
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1666464484
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1666464484
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1666464484
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1666464484
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1666464484
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1666464484
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1666464484
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1666464484
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1666464484
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1666464484
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1666464484
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1666464484
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1666464484
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1666464484
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1666464484
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1666464484
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_601
timestamp 1666464484
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_613
timestamp 1666464484
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_625
timestamp 1666464484
transform 1 0 58604 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_637
timestamp 1666464484
transform 1 0 59708 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_643
timestamp 1666464484
transform 1 0 60260 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_645
timestamp 1666464484
transform 1 0 60444 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_657
timestamp 1666464484
transform 1 0 61548 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_669
timestamp 1666464484
transform 1 0 62652 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_681
timestamp 1666464484
transform 1 0 63756 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_693
timestamp 1666464484
transform 1 0 64860 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_699
timestamp 1666464484
transform 1 0 65412 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_701
timestamp 1666464484
transform 1 0 65596 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_713
timestamp 1666464484
transform 1 0 66700 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_725
timestamp 1666464484
transform 1 0 67804 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_737
timestamp 1666464484
transform 1 0 68908 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_749
timestamp 1666464484
transform 1 0 70012 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_755
timestamp 1666464484
transform 1 0 70564 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_757
timestamp 1666464484
transform 1 0 70748 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_769
timestamp 1666464484
transform 1 0 71852 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_781
timestamp 1666464484
transform 1 0 72956 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_793
timestamp 1666464484
transform 1 0 74060 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_805
timestamp 1666464484
transform 1 0 75164 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_811
timestamp 1666464484
transform 1 0 75716 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_813
timestamp 1666464484
transform 1 0 75900 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_825
timestamp 1666464484
transform 1 0 77004 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_837
timestamp 1666464484
transform 1 0 78108 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_849
timestamp 1666464484
transform 1 0 79212 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_861
timestamp 1666464484
transform 1 0 80316 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_867
timestamp 1666464484
transform 1 0 80868 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_869
timestamp 1666464484
transform 1 0 81052 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_881
timestamp 1666464484
transform 1 0 82156 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_893
timestamp 1666464484
transform 1 0 83260 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_905
timestamp 1666464484
transform 1 0 84364 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_917
timestamp 1666464484
transform 1 0 85468 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_923
timestamp 1666464484
transform 1 0 86020 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_925
timestamp 1666464484
transform 1 0 86204 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_937
timestamp 1666464484
transform 1 0 87308 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_949
timestamp 1666464484
transform 1 0 88412 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_961
timestamp 1666464484
transform 1 0 89516 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_973
timestamp 1666464484
transform 1 0 90620 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_979
timestamp 1666464484
transform 1 0 91172 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_981
timestamp 1666464484
transform 1 0 91356 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_993
timestamp 1666464484
transform 1 0 92460 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1005
timestamp 1666464484
transform 1 0 93564 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1017
timestamp 1666464484
transform 1 0 94668 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_1029
timestamp 1666464484
transform 1 0 95772 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1035
timestamp 1666464484
transform 1 0 96324 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1037
timestamp 1666464484
transform 1 0 96508 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1049
timestamp 1666464484
transform 1 0 97612 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1061
timestamp 1666464484
transform 1 0 98716 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1073
timestamp 1666464484
transform 1 0 99820 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_1085
timestamp 1666464484
transform 1 0 100924 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1091
timestamp 1666464484
transform 1 0 101476 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1093
timestamp 1666464484
transform 1 0 101660 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1105
timestamp 1666464484
transform 1 0 102764 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1117
timestamp 1666464484
transform 1 0 103868 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1129
timestamp 1666464484
transform 1 0 104972 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_1141
timestamp 1666464484
transform 1 0 106076 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1147
timestamp 1666464484
transform 1 0 106628 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1149
timestamp 1666464484
transform 1 0 106812 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1161
timestamp 1666464484
transform 1 0 107916 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1173
timestamp 1666464484
transform 1 0 109020 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1185
timestamp 1666464484
transform 1 0 110124 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_1197
timestamp 1666464484
transform 1 0 111228 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1203
timestamp 1666464484
transform 1 0 111780 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1205
timestamp 1666464484
transform 1 0 111964 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1217
timestamp 1666464484
transform 1 0 113068 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1229
timestamp 1666464484
transform 1 0 114172 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1241
timestamp 1666464484
transform 1 0 115276 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_1253
timestamp 1666464484
transform 1 0 116380 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1259
timestamp 1666464484
transform 1 0 116932 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1261
timestamp 1666464484
transform 1 0 117116 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1273
timestamp 1666464484
transform 1 0 118220 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1285
timestamp 1666464484
transform 1 0 119324 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1297
timestamp 1666464484
transform 1 0 120428 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_1309
timestamp 1666464484
transform 1 0 121532 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1315
timestamp 1666464484
transform 1 0 122084 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1317
timestamp 1666464484
transform 1 0 122268 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1329
timestamp 1666464484
transform 1 0 123372 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1341
timestamp 1666464484
transform 1 0 124476 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1353
timestamp 1666464484
transform 1 0 125580 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_1365
timestamp 1666464484
transform 1 0 126684 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1371
timestamp 1666464484
transform 1 0 127236 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1373
timestamp 1666464484
transform 1 0 127420 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1385
timestamp 1666464484
transform 1 0 128524 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1397
timestamp 1666464484
transform 1 0 129628 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1409
timestamp 1666464484
transform 1 0 130732 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_1421
timestamp 1666464484
transform 1 0 131836 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1427
timestamp 1666464484
transform 1 0 132388 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1429
timestamp 1666464484
transform 1 0 132572 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1441
timestamp 1666464484
transform 1 0 133676 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1453
timestamp 1666464484
transform 1 0 134780 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1465
timestamp 1666464484
transform 1 0 135884 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_1477
timestamp 1666464484
transform 1 0 136988 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1483
timestamp 1666464484
transform 1 0 137540 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1485
timestamp 1666464484
transform 1 0 137724 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1497
timestamp 1666464484
transform 1 0 138828 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1509
timestamp 1666464484
transform 1 0 139932 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1521
timestamp 1666464484
transform 1 0 141036 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_1533
timestamp 1666464484
transform 1 0 142140 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1539
timestamp 1666464484
transform 1 0 142692 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1541
timestamp 1666464484
transform 1 0 142876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1553
timestamp 1666464484
transform 1 0 143980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1565
timestamp 1666464484
transform 1 0 145084 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1577
timestamp 1666464484
transform 1 0 146188 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_1589
timestamp 1666464484
transform 1 0 147292 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1595
timestamp 1666464484
transform 1 0 147844 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_1597
timestamp 1666464484
transform 1 0 148028 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1666464484
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1666464484
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1666464484
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1666464484
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1666464484
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1666464484
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1666464484
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1666464484
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1666464484
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1666464484
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1666464484
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1666464484
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1666464484
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1666464484
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1666464484
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1666464484
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1666464484
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1666464484
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1666464484
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1666464484
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1666464484
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1666464484
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1666464484
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1666464484
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1666464484
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1666464484
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1666464484
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1666464484
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1666464484
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1666464484
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1666464484
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1666464484
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1666464484
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1666464484
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1666464484
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1666464484
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1666464484
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1666464484
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1666464484
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1666464484
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1666464484
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1666464484
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1666464484
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1666464484
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1666464484
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1666464484
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1666464484
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1666464484
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1666464484
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1666464484
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1666464484
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1666464484
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1666464484
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1666464484
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1666464484
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1666464484
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1666464484
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1666464484
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1666464484
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1666464484
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1666464484
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_573
timestamp 1666464484
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_585
timestamp 1666464484
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_597
timestamp 1666464484
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1666464484
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1666464484
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_617
timestamp 1666464484
transform 1 0 57868 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_629
timestamp 1666464484
transform 1 0 58972 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_641
timestamp 1666464484
transform 1 0 60076 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_653
timestamp 1666464484
transform 1 0 61180 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_665
timestamp 1666464484
transform 1 0 62284 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_671
timestamp 1666464484
transform 1 0 62836 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_673
timestamp 1666464484
transform 1 0 63020 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_685
timestamp 1666464484
transform 1 0 64124 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_697
timestamp 1666464484
transform 1 0 65228 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_709
timestamp 1666464484
transform 1 0 66332 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_721
timestamp 1666464484
transform 1 0 67436 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_727
timestamp 1666464484
transform 1 0 67988 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_729
timestamp 1666464484
transform 1 0 68172 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_741
timestamp 1666464484
transform 1 0 69276 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_753
timestamp 1666464484
transform 1 0 70380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_765
timestamp 1666464484
transform 1 0 71484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_777
timestamp 1666464484
transform 1 0 72588 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_783
timestamp 1666464484
transform 1 0 73140 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_785
timestamp 1666464484
transform 1 0 73324 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_797
timestamp 1666464484
transform 1 0 74428 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_809
timestamp 1666464484
transform 1 0 75532 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_821
timestamp 1666464484
transform 1 0 76636 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_833
timestamp 1666464484
transform 1 0 77740 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_839
timestamp 1666464484
transform 1 0 78292 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_841
timestamp 1666464484
transform 1 0 78476 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_853
timestamp 1666464484
transform 1 0 79580 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_865
timestamp 1666464484
transform 1 0 80684 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_877
timestamp 1666464484
transform 1 0 81788 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_889
timestamp 1666464484
transform 1 0 82892 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_895
timestamp 1666464484
transform 1 0 83444 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_897
timestamp 1666464484
transform 1 0 83628 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_909
timestamp 1666464484
transform 1 0 84732 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_921
timestamp 1666464484
transform 1 0 85836 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_933
timestamp 1666464484
transform 1 0 86940 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_945
timestamp 1666464484
transform 1 0 88044 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_951
timestamp 1666464484
transform 1 0 88596 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_953
timestamp 1666464484
transform 1 0 88780 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_965
timestamp 1666464484
transform 1 0 89884 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_977
timestamp 1666464484
transform 1 0 90988 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_989
timestamp 1666464484
transform 1 0 92092 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_1001
timestamp 1666464484
transform 1 0 93196 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_1007
timestamp 1666464484
transform 1 0 93748 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1009
timestamp 1666464484
transform 1 0 93932 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1021
timestamp 1666464484
transform 1 0 95036 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1033
timestamp 1666464484
transform 1 0 96140 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1045
timestamp 1666464484
transform 1 0 97244 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_1057
timestamp 1666464484
transform 1 0 98348 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_1063
timestamp 1666464484
transform 1 0 98900 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1065
timestamp 1666464484
transform 1 0 99084 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1077
timestamp 1666464484
transform 1 0 100188 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1089
timestamp 1666464484
transform 1 0 101292 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1101
timestamp 1666464484
transform 1 0 102396 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_1113
timestamp 1666464484
transform 1 0 103500 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_1119
timestamp 1666464484
transform 1 0 104052 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1121
timestamp 1666464484
transform 1 0 104236 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1133
timestamp 1666464484
transform 1 0 105340 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1145
timestamp 1666464484
transform 1 0 106444 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1157
timestamp 1666464484
transform 1 0 107548 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_1169
timestamp 1666464484
transform 1 0 108652 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_1175
timestamp 1666464484
transform 1 0 109204 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1177
timestamp 1666464484
transform 1 0 109388 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1189
timestamp 1666464484
transform 1 0 110492 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1201
timestamp 1666464484
transform 1 0 111596 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1213
timestamp 1666464484
transform 1 0 112700 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_1225
timestamp 1666464484
transform 1 0 113804 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_1231
timestamp 1666464484
transform 1 0 114356 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1233
timestamp 1666464484
transform 1 0 114540 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1245
timestamp 1666464484
transform 1 0 115644 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1257
timestamp 1666464484
transform 1 0 116748 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1269
timestamp 1666464484
transform 1 0 117852 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_1281
timestamp 1666464484
transform 1 0 118956 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_1287
timestamp 1666464484
transform 1 0 119508 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1289
timestamp 1666464484
transform 1 0 119692 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1301
timestamp 1666464484
transform 1 0 120796 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1313
timestamp 1666464484
transform 1 0 121900 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1325
timestamp 1666464484
transform 1 0 123004 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_1337
timestamp 1666464484
transform 1 0 124108 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_1343
timestamp 1666464484
transform 1 0 124660 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1345
timestamp 1666464484
transform 1 0 124844 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1357
timestamp 1666464484
transform 1 0 125948 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1369
timestamp 1666464484
transform 1 0 127052 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1381
timestamp 1666464484
transform 1 0 128156 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_1393
timestamp 1666464484
transform 1 0 129260 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_1399
timestamp 1666464484
transform 1 0 129812 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1401
timestamp 1666464484
transform 1 0 129996 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1413
timestamp 1666464484
transform 1 0 131100 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1425
timestamp 1666464484
transform 1 0 132204 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1437
timestamp 1666464484
transform 1 0 133308 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_1449
timestamp 1666464484
transform 1 0 134412 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_1455
timestamp 1666464484
transform 1 0 134964 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1457
timestamp 1666464484
transform 1 0 135148 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1469
timestamp 1666464484
transform 1 0 136252 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1481
timestamp 1666464484
transform 1 0 137356 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1493
timestamp 1666464484
transform 1 0 138460 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_1505
timestamp 1666464484
transform 1 0 139564 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_1511
timestamp 1666464484
transform 1 0 140116 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1513
timestamp 1666464484
transform 1 0 140300 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1525
timestamp 1666464484
transform 1 0 141404 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1537
timestamp 1666464484
transform 1 0 142508 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1549
timestamp 1666464484
transform 1 0 143612 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_1561
timestamp 1666464484
transform 1 0 144716 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_1567
timestamp 1666464484
transform 1 0 145268 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1569
timestamp 1666464484
transform 1 0 145452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1581
timestamp 1666464484
transform 1 0 146556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_1593
timestamp 1666464484
transform 1 0 147660 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_1601
timestamp 1666464484
transform 1 0 148396 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1666464484
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1666464484
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1666464484
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1666464484
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1666464484
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1666464484
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1666464484
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1666464484
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1666464484
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1666464484
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1666464484
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1666464484
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1666464484
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1666464484
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1666464484
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1666464484
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1666464484
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1666464484
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1666464484
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1666464484
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1666464484
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1666464484
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1666464484
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1666464484
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1666464484
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1666464484
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1666464484
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1666464484
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1666464484
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1666464484
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1666464484
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1666464484
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1666464484
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1666464484
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1666464484
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1666464484
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1666464484
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1666464484
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1666464484
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1666464484
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1666464484
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1666464484
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1666464484
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1666464484
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1666464484
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1666464484
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1666464484
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1666464484
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1666464484
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1666464484
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1666464484
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1666464484
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1666464484
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1666464484
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1666464484
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1666464484
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1666464484
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1666464484
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1666464484
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1666464484
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_569
timestamp 1666464484
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1666464484
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1666464484
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1666464484
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_601
timestamp 1666464484
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_613
timestamp 1666464484
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_625
timestamp 1666464484
transform 1 0 58604 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_637
timestamp 1666464484
transform 1 0 59708 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_643
timestamp 1666464484
transform 1 0 60260 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_645
timestamp 1666464484
transform 1 0 60444 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_657
timestamp 1666464484
transform 1 0 61548 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_669
timestamp 1666464484
transform 1 0 62652 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_681
timestamp 1666464484
transform 1 0 63756 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_693
timestamp 1666464484
transform 1 0 64860 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_699
timestamp 1666464484
transform 1 0 65412 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_701
timestamp 1666464484
transform 1 0 65596 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_713
timestamp 1666464484
transform 1 0 66700 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_725
timestamp 1666464484
transform 1 0 67804 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_737
timestamp 1666464484
transform 1 0 68908 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_749
timestamp 1666464484
transform 1 0 70012 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_755
timestamp 1666464484
transform 1 0 70564 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_757
timestamp 1666464484
transform 1 0 70748 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_769
timestamp 1666464484
transform 1 0 71852 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_781
timestamp 1666464484
transform 1 0 72956 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_793
timestamp 1666464484
transform 1 0 74060 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_805
timestamp 1666464484
transform 1 0 75164 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_811
timestamp 1666464484
transform 1 0 75716 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_813
timestamp 1666464484
transform 1 0 75900 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_825
timestamp 1666464484
transform 1 0 77004 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_837
timestamp 1666464484
transform 1 0 78108 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_849
timestamp 1666464484
transform 1 0 79212 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_861
timestamp 1666464484
transform 1 0 80316 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_867
timestamp 1666464484
transform 1 0 80868 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_869
timestamp 1666464484
transform 1 0 81052 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_881
timestamp 1666464484
transform 1 0 82156 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_893
timestamp 1666464484
transform 1 0 83260 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_905
timestamp 1666464484
transform 1 0 84364 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_917
timestamp 1666464484
transform 1 0 85468 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_923
timestamp 1666464484
transform 1 0 86020 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_925
timestamp 1666464484
transform 1 0 86204 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_937
timestamp 1666464484
transform 1 0 87308 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_949
timestamp 1666464484
transform 1 0 88412 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_961
timestamp 1666464484
transform 1 0 89516 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_973
timestamp 1666464484
transform 1 0 90620 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_979
timestamp 1666464484
transform 1 0 91172 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_981
timestamp 1666464484
transform 1 0 91356 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_993
timestamp 1666464484
transform 1 0 92460 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1005
timestamp 1666464484
transform 1 0 93564 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1017
timestamp 1666464484
transform 1 0 94668 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_1029
timestamp 1666464484
transform 1 0 95772 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1035
timestamp 1666464484
transform 1 0 96324 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1037
timestamp 1666464484
transform 1 0 96508 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1049
timestamp 1666464484
transform 1 0 97612 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1061
timestamp 1666464484
transform 1 0 98716 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1073
timestamp 1666464484
transform 1 0 99820 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_1085
timestamp 1666464484
transform 1 0 100924 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1091
timestamp 1666464484
transform 1 0 101476 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1093
timestamp 1666464484
transform 1 0 101660 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1105
timestamp 1666464484
transform 1 0 102764 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1117
timestamp 1666464484
transform 1 0 103868 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1129
timestamp 1666464484
transform 1 0 104972 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_1141
timestamp 1666464484
transform 1 0 106076 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1147
timestamp 1666464484
transform 1 0 106628 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1149
timestamp 1666464484
transform 1 0 106812 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1161
timestamp 1666464484
transform 1 0 107916 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1173
timestamp 1666464484
transform 1 0 109020 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1185
timestamp 1666464484
transform 1 0 110124 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_1197
timestamp 1666464484
transform 1 0 111228 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1203
timestamp 1666464484
transform 1 0 111780 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1205
timestamp 1666464484
transform 1 0 111964 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1217
timestamp 1666464484
transform 1 0 113068 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1229
timestamp 1666464484
transform 1 0 114172 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1241
timestamp 1666464484
transform 1 0 115276 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_1253
timestamp 1666464484
transform 1 0 116380 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1259
timestamp 1666464484
transform 1 0 116932 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1261
timestamp 1666464484
transform 1 0 117116 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1273
timestamp 1666464484
transform 1 0 118220 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1285
timestamp 1666464484
transform 1 0 119324 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1297
timestamp 1666464484
transform 1 0 120428 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_1309
timestamp 1666464484
transform 1 0 121532 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1315
timestamp 1666464484
transform 1 0 122084 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1317
timestamp 1666464484
transform 1 0 122268 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1329
timestamp 1666464484
transform 1 0 123372 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1341
timestamp 1666464484
transform 1 0 124476 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1353
timestamp 1666464484
transform 1 0 125580 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_1365
timestamp 1666464484
transform 1 0 126684 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1371
timestamp 1666464484
transform 1 0 127236 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1373
timestamp 1666464484
transform 1 0 127420 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1385
timestamp 1666464484
transform 1 0 128524 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1397
timestamp 1666464484
transform 1 0 129628 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1409
timestamp 1666464484
transform 1 0 130732 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_1421
timestamp 1666464484
transform 1 0 131836 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1427
timestamp 1666464484
transform 1 0 132388 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1429
timestamp 1666464484
transform 1 0 132572 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1441
timestamp 1666464484
transform 1 0 133676 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1453
timestamp 1666464484
transform 1 0 134780 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1465
timestamp 1666464484
transform 1 0 135884 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_1477
timestamp 1666464484
transform 1 0 136988 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1483
timestamp 1666464484
transform 1 0 137540 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1485
timestamp 1666464484
transform 1 0 137724 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1497
timestamp 1666464484
transform 1 0 138828 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1509
timestamp 1666464484
transform 1 0 139932 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1521
timestamp 1666464484
transform 1 0 141036 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_1533
timestamp 1666464484
transform 1 0 142140 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1539
timestamp 1666464484
transform 1 0 142692 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1541
timestamp 1666464484
transform 1 0 142876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1553
timestamp 1666464484
transform 1 0 143980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1565
timestamp 1666464484
transform 1 0 145084 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1577
timestamp 1666464484
transform 1 0 146188 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_1589
timestamp 1666464484
transform 1 0 147292 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1595
timestamp 1666464484
transform 1 0 147844 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_1597
timestamp 1666464484
transform 1 0 148028 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1666464484
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1666464484
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1666464484
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1666464484
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1666464484
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1666464484
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1666464484
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1666464484
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1666464484
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1666464484
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1666464484
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1666464484
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1666464484
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1666464484
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1666464484
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1666464484
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1666464484
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1666464484
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1666464484
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1666464484
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1666464484
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1666464484
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1666464484
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1666464484
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1666464484
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1666464484
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1666464484
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1666464484
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1666464484
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1666464484
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1666464484
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1666464484
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1666464484
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1666464484
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1666464484
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1666464484
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1666464484
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1666464484
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1666464484
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1666464484
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1666464484
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1666464484
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1666464484
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1666464484
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1666464484
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1666464484
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1666464484
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1666464484
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1666464484
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_461
timestamp 1666464484
transform 1 0 43516 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_465
timestamp 1666464484
transform 1 0 43884 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_477
timestamp 1666464484
transform 1 0 44988 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_489
timestamp 1666464484
transform 1 0 46092 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_501
timestamp 1666464484
transform 1 0 47196 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1666464484
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1666464484
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1666464484
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1666464484
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1666464484
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1666464484
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1666464484
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_573
timestamp 1666464484
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_585
timestamp 1666464484
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_597
timestamp 1666464484
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1666464484
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1666464484
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_617
timestamp 1666464484
transform 1 0 57868 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_629
timestamp 1666464484
transform 1 0 58972 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_641
timestamp 1666464484
transform 1 0 60076 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_653
timestamp 1666464484
transform 1 0 61180 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_665
timestamp 1666464484
transform 1 0 62284 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_671
timestamp 1666464484
transform 1 0 62836 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_673
timestamp 1666464484
transform 1 0 63020 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_685
timestamp 1666464484
transform 1 0 64124 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_697
timestamp 1666464484
transform 1 0 65228 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_709
timestamp 1666464484
transform 1 0 66332 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_721
timestamp 1666464484
transform 1 0 67436 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_727
timestamp 1666464484
transform 1 0 67988 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_729
timestamp 1666464484
transform 1 0 68172 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_741
timestamp 1666464484
transform 1 0 69276 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_753
timestamp 1666464484
transform 1 0 70380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_765
timestamp 1666464484
transform 1 0 71484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_777
timestamp 1666464484
transform 1 0 72588 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_783
timestamp 1666464484
transform 1 0 73140 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_785
timestamp 1666464484
transform 1 0 73324 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_797
timestamp 1666464484
transform 1 0 74428 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_809
timestamp 1666464484
transform 1 0 75532 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_821
timestamp 1666464484
transform 1 0 76636 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_833
timestamp 1666464484
transform 1 0 77740 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_839
timestamp 1666464484
transform 1 0 78292 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_841
timestamp 1666464484
transform 1 0 78476 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_853
timestamp 1666464484
transform 1 0 79580 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_865
timestamp 1666464484
transform 1 0 80684 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_877
timestamp 1666464484
transform 1 0 81788 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_889
timestamp 1666464484
transform 1 0 82892 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_895
timestamp 1666464484
transform 1 0 83444 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_897
timestamp 1666464484
transform 1 0 83628 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_909
timestamp 1666464484
transform 1 0 84732 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_921
timestamp 1666464484
transform 1 0 85836 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_933
timestamp 1666464484
transform 1 0 86940 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_945
timestamp 1666464484
transform 1 0 88044 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_951
timestamp 1666464484
transform 1 0 88596 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_953
timestamp 1666464484
transform 1 0 88780 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_965
timestamp 1666464484
transform 1 0 89884 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_977
timestamp 1666464484
transform 1 0 90988 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_989
timestamp 1666464484
transform 1 0 92092 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_1001
timestamp 1666464484
transform 1 0 93196 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_1007
timestamp 1666464484
transform 1 0 93748 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1009
timestamp 1666464484
transform 1 0 93932 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1021
timestamp 1666464484
transform 1 0 95036 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1033
timestamp 1666464484
transform 1 0 96140 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1045
timestamp 1666464484
transform 1 0 97244 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_1057
timestamp 1666464484
transform 1 0 98348 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_1063
timestamp 1666464484
transform 1 0 98900 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1065
timestamp 1666464484
transform 1 0 99084 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1077
timestamp 1666464484
transform 1 0 100188 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1089
timestamp 1666464484
transform 1 0 101292 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1101
timestamp 1666464484
transform 1 0 102396 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_1113
timestamp 1666464484
transform 1 0 103500 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_1119
timestamp 1666464484
transform 1 0 104052 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1121
timestamp 1666464484
transform 1 0 104236 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1133
timestamp 1666464484
transform 1 0 105340 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1145
timestamp 1666464484
transform 1 0 106444 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1157
timestamp 1666464484
transform 1 0 107548 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_1169
timestamp 1666464484
transform 1 0 108652 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_1175
timestamp 1666464484
transform 1 0 109204 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1177
timestamp 1666464484
transform 1 0 109388 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1189
timestamp 1666464484
transform 1 0 110492 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1201
timestamp 1666464484
transform 1 0 111596 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1213
timestamp 1666464484
transform 1 0 112700 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_1225
timestamp 1666464484
transform 1 0 113804 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_1231
timestamp 1666464484
transform 1 0 114356 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1233
timestamp 1666464484
transform 1 0 114540 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1245
timestamp 1666464484
transform 1 0 115644 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1257
timestamp 1666464484
transform 1 0 116748 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1269
timestamp 1666464484
transform 1 0 117852 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_1281
timestamp 1666464484
transform 1 0 118956 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_1287
timestamp 1666464484
transform 1 0 119508 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1289
timestamp 1666464484
transform 1 0 119692 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1301
timestamp 1666464484
transform 1 0 120796 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1313
timestamp 1666464484
transform 1 0 121900 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1325
timestamp 1666464484
transform 1 0 123004 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_1337
timestamp 1666464484
transform 1 0 124108 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_1343
timestamp 1666464484
transform 1 0 124660 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1345
timestamp 1666464484
transform 1 0 124844 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1357
timestamp 1666464484
transform 1 0 125948 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1369
timestamp 1666464484
transform 1 0 127052 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1381
timestamp 1666464484
transform 1 0 128156 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_1393
timestamp 1666464484
transform 1 0 129260 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_1399
timestamp 1666464484
transform 1 0 129812 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1401
timestamp 1666464484
transform 1 0 129996 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1413
timestamp 1666464484
transform 1 0 131100 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1425
timestamp 1666464484
transform 1 0 132204 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1437
timestamp 1666464484
transform 1 0 133308 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_1449
timestamp 1666464484
transform 1 0 134412 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_1455
timestamp 1666464484
transform 1 0 134964 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1457
timestamp 1666464484
transform 1 0 135148 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1469
timestamp 1666464484
transform 1 0 136252 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1481
timestamp 1666464484
transform 1 0 137356 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1493
timestamp 1666464484
transform 1 0 138460 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_1505
timestamp 1666464484
transform 1 0 139564 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_1511
timestamp 1666464484
transform 1 0 140116 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1513
timestamp 1666464484
transform 1 0 140300 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1525
timestamp 1666464484
transform 1 0 141404 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1537
timestamp 1666464484
transform 1 0 142508 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1549
timestamp 1666464484
transform 1 0 143612 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_1561
timestamp 1666464484
transform 1 0 144716 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_1567
timestamp 1666464484
transform 1 0 145268 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1569
timestamp 1666464484
transform 1 0 145452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1581
timestamp 1666464484
transform 1 0 146556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_1593
timestamp 1666464484
transform 1 0 147660 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_1601
timestamp 1666464484
transform 1 0 148396 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1666464484
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1666464484
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1666464484
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1666464484
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1666464484
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1666464484
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1666464484
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1666464484
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1666464484
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1666464484
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1666464484
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1666464484
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1666464484
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1666464484
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1666464484
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1666464484
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1666464484
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1666464484
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1666464484
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1666464484
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1666464484
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1666464484
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_209
timestamp 1666464484
transform 1 0 20332 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_215
timestamp 1666464484
transform 1 0 20884 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_218
timestamp 1666464484
transform 1 0 21160 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_230
timestamp 1666464484
transform 1 0 22264 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_242
timestamp 1666464484
transform 1 0 23368 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1666464484
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_253
timestamp 1666464484
transform 1 0 24380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_259
timestamp 1666464484
transform 1 0 24932 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_263
timestamp 1666464484
transform 1 0 25300 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_266
timestamp 1666464484
transform 1 0 25576 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_272
timestamp 1666464484
transform 1 0 26128 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_284
timestamp 1666464484
transform 1 0 27232 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_296
timestamp 1666464484
transform 1 0 28336 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1666464484
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1666464484
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1666464484
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1666464484
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1666464484
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1666464484
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1666464484
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1666464484
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1666464484
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_377
timestamp 1666464484
transform 1 0 35788 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_381
timestamp 1666464484
transform 1 0 36156 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_389
timestamp 1666464484
transform 1 0 36892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_392
timestamp 1666464484
transform 1 0 37168 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_398
timestamp 1666464484
transform 1 0 37720 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_406
timestamp 1666464484
transform 1 0 38456 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_411
timestamp 1666464484
transform 1 0 38916 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1666464484
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_421
timestamp 1666464484
transform 1 0 39836 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_431
timestamp 1666464484
transform 1 0 40756 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_439
timestamp 1666464484
transform 1 0 41492 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_442
timestamp 1666464484
transform 1 0 41768 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_450
timestamp 1666464484
transform 1 0 42504 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_454
timestamp 1666464484
transform 1 0 42872 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_60_462
timestamp 1666464484
transform 1 0 43608 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_60_470
timestamp 1666464484
transform 1 0 44344 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_60_477
timestamp 1666464484
transform 1 0 44988 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_485
timestamp 1666464484
transform 1 0 45724 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_497
timestamp 1666464484
transform 1 0 46828 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_505
timestamp 1666464484
transform 1 0 47564 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_508
timestamp 1666464484
transform 1 0 47840 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_518
timestamp 1666464484
transform 1 0 48760 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_530
timestamp 1666464484
transform 1 0 49864 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_533
timestamp 1666464484
transform 1 0 50140 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_537
timestamp 1666464484
transform 1 0 50508 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_547
timestamp 1666464484
transform 1 0 51428 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_559
timestamp 1666464484
transform 1 0 52532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_571
timestamp 1666464484
transform 1 0 53636 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_574
timestamp 1666464484
transform 1 0 53912 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_586
timestamp 1666464484
transform 1 0 55016 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_589
timestamp 1666464484
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_601
timestamp 1666464484
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_613
timestamp 1666464484
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_625
timestamp 1666464484
transform 1 0 58604 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_630
timestamp 1666464484
transform 1 0 59064 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_638
timestamp 1666464484
transform 1 0 59800 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_60_641
timestamp 1666464484
transform 1 0 60076 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_645
timestamp 1666464484
transform 1 0 60444 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_649
timestamp 1666464484
transform 1 0 60812 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_655
timestamp 1666464484
transform 1 0 61364 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_661
timestamp 1666464484
transform 1 0 61916 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_667
timestamp 1666464484
transform 1 0 62468 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_671
timestamp 1666464484
transform 1 0 62836 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_674
timestamp 1666464484
transform 1 0 63112 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_682
timestamp 1666464484
transform 1 0 63848 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_688
timestamp 1666464484
transform 1 0 64400 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_698
timestamp 1666464484
transform 1 0 65320 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_701
timestamp 1666464484
transform 1 0 65596 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_706
timestamp 1666464484
transform 1 0 66056 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_718
timestamp 1666464484
transform 1 0 67160 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_730
timestamp 1666464484
transform 1 0 68264 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_738
timestamp 1666464484
transform 1 0 69000 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_742
timestamp 1666464484
transform 1 0 69368 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_754
timestamp 1666464484
transform 1 0 70472 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_757
timestamp 1666464484
transform 1 0 70748 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_769
timestamp 1666464484
transform 1 0 71852 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_781
timestamp 1666464484
transform 1 0 72956 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_793
timestamp 1666464484
transform 1 0 74060 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_805
timestamp 1666464484
transform 1 0 75164 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_811
timestamp 1666464484
transform 1 0 75716 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_813
timestamp 1666464484
transform 1 0 75900 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_825
timestamp 1666464484
transform 1 0 77004 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_837
timestamp 1666464484
transform 1 0 78108 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_849
timestamp 1666464484
transform 1 0 79212 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_854
timestamp 1666464484
transform 1 0 79672 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_860
timestamp 1666464484
transform 1 0 80224 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_866
timestamp 1666464484
transform 1 0 80776 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_869
timestamp 1666464484
transform 1 0 81052 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_873
timestamp 1666464484
transform 1 0 81420 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_879
timestamp 1666464484
transform 1 0 81972 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_885
timestamp 1666464484
transform 1 0 82524 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_897
timestamp 1666464484
transform 1 0 83628 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_909
timestamp 1666464484
transform 1 0 84732 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_921
timestamp 1666464484
transform 1 0 85836 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_925
timestamp 1666464484
transform 1 0 86204 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_937
timestamp 1666464484
transform 1 0 87308 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_949
timestamp 1666464484
transform 1 0 88412 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_961
timestamp 1666464484
transform 1 0 89516 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_973
timestamp 1666464484
transform 1 0 90620 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_979
timestamp 1666464484
transform 1 0 91172 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_981
timestamp 1666464484
transform 1 0 91356 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_993
timestamp 1666464484
transform 1 0 92460 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1005
timestamp 1666464484
transform 1 0 93564 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1017
timestamp 1666464484
transform 1 0 94668 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_1029
timestamp 1666464484
transform 1 0 95772 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1035
timestamp 1666464484
transform 1 0 96324 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1037
timestamp 1666464484
transform 1 0 96508 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1049
timestamp 1666464484
transform 1 0 97612 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1061
timestamp 1666464484
transform 1 0 98716 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1073
timestamp 1666464484
transform 1 0 99820 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_1085
timestamp 1666464484
transform 1 0 100924 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1091
timestamp 1666464484
transform 1 0 101476 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1093
timestamp 1666464484
transform 1 0 101660 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1105
timestamp 1666464484
transform 1 0 102764 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1117
timestamp 1666464484
transform 1 0 103868 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1129
timestamp 1666464484
transform 1 0 104972 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_1141
timestamp 1666464484
transform 1 0 106076 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1147
timestamp 1666464484
transform 1 0 106628 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1149
timestamp 1666464484
transform 1 0 106812 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1161
timestamp 1666464484
transform 1 0 107916 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1173
timestamp 1666464484
transform 1 0 109020 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1185
timestamp 1666464484
transform 1 0 110124 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_1197
timestamp 1666464484
transform 1 0 111228 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1203
timestamp 1666464484
transform 1 0 111780 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1205
timestamp 1666464484
transform 1 0 111964 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1217
timestamp 1666464484
transform 1 0 113068 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1229
timestamp 1666464484
transform 1 0 114172 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1241
timestamp 1666464484
transform 1 0 115276 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_1253
timestamp 1666464484
transform 1 0 116380 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1259
timestamp 1666464484
transform 1 0 116932 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1261
timestamp 1666464484
transform 1 0 117116 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1273
timestamp 1666464484
transform 1 0 118220 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1285
timestamp 1666464484
transform 1 0 119324 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1297
timestamp 1666464484
transform 1 0 120428 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_1309
timestamp 1666464484
transform 1 0 121532 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1315
timestamp 1666464484
transform 1 0 122084 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1317
timestamp 1666464484
transform 1 0 122268 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1329
timestamp 1666464484
transform 1 0 123372 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1341
timestamp 1666464484
transform 1 0 124476 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1353
timestamp 1666464484
transform 1 0 125580 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_1365
timestamp 1666464484
transform 1 0 126684 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1371
timestamp 1666464484
transform 1 0 127236 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1373
timestamp 1666464484
transform 1 0 127420 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1385
timestamp 1666464484
transform 1 0 128524 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1397
timestamp 1666464484
transform 1 0 129628 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1409
timestamp 1666464484
transform 1 0 130732 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_1421
timestamp 1666464484
transform 1 0 131836 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1427
timestamp 1666464484
transform 1 0 132388 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1429
timestamp 1666464484
transform 1 0 132572 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1441
timestamp 1666464484
transform 1 0 133676 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1453
timestamp 1666464484
transform 1 0 134780 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1465
timestamp 1666464484
transform 1 0 135884 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_1477
timestamp 1666464484
transform 1 0 136988 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1483
timestamp 1666464484
transform 1 0 137540 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1485
timestamp 1666464484
transform 1 0 137724 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1497
timestamp 1666464484
transform 1 0 138828 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1509
timestamp 1666464484
transform 1 0 139932 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1521
timestamp 1666464484
transform 1 0 141036 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_1533
timestamp 1666464484
transform 1 0 142140 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1539
timestamp 1666464484
transform 1 0 142692 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1541
timestamp 1666464484
transform 1 0 142876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1553
timestamp 1666464484
transform 1 0 143980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1565
timestamp 1666464484
transform 1 0 145084 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1577
timestamp 1666464484
transform 1 0 146188 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_1589
timestamp 1666464484
transform 1 0 147292 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1595
timestamp 1666464484
transform 1 0 147844 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_1597
timestamp 1666464484
transform 1 0 148028 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1666464484
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1666464484
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1666464484
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1666464484
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1666464484
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1666464484
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1666464484
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1666464484
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1666464484
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1666464484
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1666464484
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1666464484
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1666464484
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1666464484
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1666464484
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1666464484
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1666464484
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1666464484
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1666464484
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1666464484
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_193
timestamp 1666464484
transform 1 0 18860 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_201
timestamp 1666464484
transform 1 0 19596 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_205
timestamp 1666464484
transform 1 0 19964 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_213
timestamp 1666464484
transform 1 0 20700 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_61_218
timestamp 1666464484
transform 1 0 21160 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1666464484
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1666464484
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_249
timestamp 1666464484
transform 1 0 24012 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_252
timestamp 1666464484
transform 1 0 24288 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_258
timestamp 1666464484
transform 1 0 24840 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_264
timestamp 1666464484
transform 1 0 25392 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_270
timestamp 1666464484
transform 1 0 25944 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_61_278
timestamp 1666464484
transform 1 0 26680 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_281
timestamp 1666464484
transform 1 0 26956 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_289
timestamp 1666464484
transform 1 0 27692 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_294
timestamp 1666464484
transform 1 0 28152 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_300
timestamp 1666464484
transform 1 0 28704 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_306
timestamp 1666464484
transform 1 0 29256 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_318
timestamp 1666464484
transform 1 0 30360 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_326
timestamp 1666464484
transform 1 0 31096 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_61_334
timestamp 1666464484
transform 1 0 31832 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_337
timestamp 1666464484
transform 1 0 32108 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_345
timestamp 1666464484
transform 1 0 32844 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_350
timestamp 1666464484
transform 1 0 33304 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_364
timestamp 1666464484
transform 1 0 34592 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_372
timestamp 1666464484
transform 1 0 35328 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_378
timestamp 1666464484
transform 1 0 35880 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_384
timestamp 1666464484
transform 1 0 36432 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_390
timestamp 1666464484
transform 1 0 36984 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_393
timestamp 1666464484
transform 1 0 37260 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_398
timestamp 1666464484
transform 1 0 37720 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_404
timestamp 1666464484
transform 1 0 38272 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_410
timestamp 1666464484
transform 1 0 38824 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_416
timestamp 1666464484
transform 1 0 39376 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_422
timestamp 1666464484
transform 1 0 39928 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_428
timestamp 1666464484
transform 1 0 40480 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_434
timestamp 1666464484
transform 1 0 41032 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_440
timestamp 1666464484
transform 1 0 41584 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_446
timestamp 1666464484
transform 1 0 42136 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_449
timestamp 1666464484
transform 1 0 42412 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_454
timestamp 1666464484
transform 1 0 42872 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_458
timestamp 1666464484
transform 1 0 43240 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_461
timestamp 1666464484
transform 1 0 43516 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_467
timestamp 1666464484
transform 1 0 44068 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_473
timestamp 1666464484
transform 1 0 44620 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_477
timestamp 1666464484
transform 1 0 44988 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_480
timestamp 1666464484
transform 1 0 45264 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_490
timestamp 1666464484
transform 1 0 46184 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_496
timestamp 1666464484
transform 1 0 46736 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_502
timestamp 1666464484
transform 1 0 47288 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_505
timestamp 1666464484
transform 1 0 47564 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_509
timestamp 1666464484
transform 1 0 47932 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_512
timestamp 1666464484
transform 1 0 48208 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_518
timestamp 1666464484
transform 1 0 48760 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_524
timestamp 1666464484
transform 1 0 49312 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_532
timestamp 1666464484
transform 1 0 50048 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_538
timestamp 1666464484
transform 1 0 50600 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_546
timestamp 1666464484
transform 1 0 51336 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_552
timestamp 1666464484
transform 1 0 51888 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_558
timestamp 1666464484
transform 1 0 52440 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_561
timestamp 1666464484
transform 1 0 52716 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_566
timestamp 1666464484
transform 1 0 53176 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_574
timestamp 1666464484
transform 1 0 53912 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_577
timestamp 1666464484
transform 1 0 54188 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_585
timestamp 1666464484
transform 1 0 54924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_588
timestamp 1666464484
transform 1 0 55200 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_61_598
timestamp 1666464484
transform 1 0 56120 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_608
timestamp 1666464484
transform 1 0 57040 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_614
timestamp 1666464484
transform 1 0 57592 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_617
timestamp 1666464484
transform 1 0 57868 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_621
timestamp 1666464484
transform 1 0 58236 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_627
timestamp 1666464484
transform 1 0 58788 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_631
timestamp 1666464484
transform 1 0 59156 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_634
timestamp 1666464484
transform 1 0 59432 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_640
timestamp 1666464484
transform 1 0 59984 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_646
timestamp 1666464484
transform 1 0 60536 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_652
timestamp 1666464484
transform 1 0 61088 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_658
timestamp 1666464484
transform 1 0 61640 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_664
timestamp 1666464484
transform 1 0 62192 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_670
timestamp 1666464484
transform 1 0 62744 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_673
timestamp 1666464484
transform 1 0 63020 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_679
timestamp 1666464484
transform 1 0 63572 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_682
timestamp 1666464484
transform 1 0 63848 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_688
timestamp 1666464484
transform 1 0 64400 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_694
timestamp 1666464484
transform 1 0 64952 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_701
timestamp 1666464484
transform 1 0 65596 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_707
timestamp 1666464484
transform 1 0 66148 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_711
timestamp 1666464484
transform 1 0 66516 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_714
timestamp 1666464484
transform 1 0 66792 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_720
timestamp 1666464484
transform 1 0 67344 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_729
timestamp 1666464484
transform 1 0 68172 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_61_734
timestamp 1666464484
transform 1 0 68632 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_742
timestamp 1666464484
transform 1 0 69368 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_748
timestamp 1666464484
transform 1 0 69920 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_760
timestamp 1666464484
transform 1 0 71024 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_772
timestamp 1666464484
transform 1 0 72128 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_785
timestamp 1666464484
transform 1 0 73324 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_797
timestamp 1666464484
transform 1 0 74428 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_803
timestamp 1666464484
transform 1 0 74980 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_806
timestamp 1666464484
transform 1 0 75256 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_818
timestamp 1666464484
transform 1 0 76360 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_830
timestamp 1666464484
transform 1 0 77464 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_838
timestamp 1666464484
transform 1 0 78200 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_841
timestamp 1666464484
transform 1 0 78476 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_847
timestamp 1666464484
transform 1 0 79028 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_855
timestamp 1666464484
transform 1 0 79764 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_858
timestamp 1666464484
transform 1 0 80040 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_864
timestamp 1666464484
transform 1 0 80592 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_872
timestamp 1666464484
transform 1 0 81328 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_878
timestamp 1666464484
transform 1 0 81880 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_884
timestamp 1666464484
transform 1 0 82432 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_890
timestamp 1666464484
transform 1 0 82984 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_61_897
timestamp 1666464484
transform 1 0 83628 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_901
timestamp 1666464484
transform 1 0 83996 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_907
timestamp 1666464484
transform 1 0 84548 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_915
timestamp 1666464484
transform 1 0 85284 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_927
timestamp 1666464484
transform 1 0 86388 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_939
timestamp 1666464484
transform 1 0 87492 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_951
timestamp 1666464484
transform 1 0 88596 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_953
timestamp 1666464484
transform 1 0 88780 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_965
timestamp 1666464484
transform 1 0 89884 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_977
timestamp 1666464484
transform 1 0 90988 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_989
timestamp 1666464484
transform 1 0 92092 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_1001
timestamp 1666464484
transform 1 0 93196 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_1007
timestamp 1666464484
transform 1 0 93748 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1009
timestamp 1666464484
transform 1 0 93932 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1021
timestamp 1666464484
transform 1 0 95036 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1033
timestamp 1666464484
transform 1 0 96140 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1045
timestamp 1666464484
transform 1 0 97244 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_1057
timestamp 1666464484
transform 1 0 98348 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_1063
timestamp 1666464484
transform 1 0 98900 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1065
timestamp 1666464484
transform 1 0 99084 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1077
timestamp 1666464484
transform 1 0 100188 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1089
timestamp 1666464484
transform 1 0 101292 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1101
timestamp 1666464484
transform 1 0 102396 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_1113
timestamp 1666464484
transform 1 0 103500 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_1119
timestamp 1666464484
transform 1 0 104052 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1121
timestamp 1666464484
transform 1 0 104236 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1133
timestamp 1666464484
transform 1 0 105340 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1145
timestamp 1666464484
transform 1 0 106444 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1157
timestamp 1666464484
transform 1 0 107548 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_1169
timestamp 1666464484
transform 1 0 108652 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_1175
timestamp 1666464484
transform 1 0 109204 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1177
timestamp 1666464484
transform 1 0 109388 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1189
timestamp 1666464484
transform 1 0 110492 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1201
timestamp 1666464484
transform 1 0 111596 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1213
timestamp 1666464484
transform 1 0 112700 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_1225
timestamp 1666464484
transform 1 0 113804 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_1231
timestamp 1666464484
transform 1 0 114356 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1233
timestamp 1666464484
transform 1 0 114540 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1245
timestamp 1666464484
transform 1 0 115644 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1257
timestamp 1666464484
transform 1 0 116748 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1269
timestamp 1666464484
transform 1 0 117852 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_1281
timestamp 1666464484
transform 1 0 118956 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_1287
timestamp 1666464484
transform 1 0 119508 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1289
timestamp 1666464484
transform 1 0 119692 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1301
timestamp 1666464484
transform 1 0 120796 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1313
timestamp 1666464484
transform 1 0 121900 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1325
timestamp 1666464484
transform 1 0 123004 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_1337
timestamp 1666464484
transform 1 0 124108 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_1343
timestamp 1666464484
transform 1 0 124660 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1345
timestamp 1666464484
transform 1 0 124844 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1357
timestamp 1666464484
transform 1 0 125948 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1369
timestamp 1666464484
transform 1 0 127052 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1381
timestamp 1666464484
transform 1 0 128156 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_1393
timestamp 1666464484
transform 1 0 129260 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_1399
timestamp 1666464484
transform 1 0 129812 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1401
timestamp 1666464484
transform 1 0 129996 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1413
timestamp 1666464484
transform 1 0 131100 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1425
timestamp 1666464484
transform 1 0 132204 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1437
timestamp 1666464484
transform 1 0 133308 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_1449
timestamp 1666464484
transform 1 0 134412 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_1455
timestamp 1666464484
transform 1 0 134964 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1457
timestamp 1666464484
transform 1 0 135148 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1469
timestamp 1666464484
transform 1 0 136252 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1481
timestamp 1666464484
transform 1 0 137356 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1493
timestamp 1666464484
transform 1 0 138460 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_1505
timestamp 1666464484
transform 1 0 139564 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_1511
timestamp 1666464484
transform 1 0 140116 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1513
timestamp 1666464484
transform 1 0 140300 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1525
timestamp 1666464484
transform 1 0 141404 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1537
timestamp 1666464484
transform 1 0 142508 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1549
timestamp 1666464484
transform 1 0 143612 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_1561
timestamp 1666464484
transform 1 0 144716 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_1567
timestamp 1666464484
transform 1 0 145268 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1569
timestamp 1666464484
transform 1 0 145452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1581
timestamp 1666464484
transform 1 0 146556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_1593
timestamp 1666464484
transform 1 0 147660 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_1601
timestamp 1666464484
transform 1 0 148396 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1666464484
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1666464484
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1666464484
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1666464484
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1666464484
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_53
timestamp 1666464484
transform 1 0 5980 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_61
timestamp 1666464484
transform 1 0 6716 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_64
timestamp 1666464484
transform 1 0 6992 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_76
timestamp 1666464484
transform 1 0 8096 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_85
timestamp 1666464484
transform 1 0 8924 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_89
timestamp 1666464484
transform 1 0 9292 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_95
timestamp 1666464484
transform 1 0 9844 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_98
timestamp 1666464484
transform 1 0 10120 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_110
timestamp 1666464484
transform 1 0 11224 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_122
timestamp 1666464484
transform 1 0 12328 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_134
timestamp 1666464484
transform 1 0 13432 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1666464484
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1666464484
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1666464484
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_179
timestamp 1666464484
transform 1 0 17572 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_191
timestamp 1666464484
transform 1 0 18676 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1666464484
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_197
timestamp 1666464484
transform 1 0 19228 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_202
timestamp 1666464484
transform 1 0 19688 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_208
timestamp 1666464484
transform 1 0 20240 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_214
timestamp 1666464484
transform 1 0 20792 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_221
timestamp 1666464484
transform 1 0 21436 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_227
timestamp 1666464484
transform 1 0 21988 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_231
timestamp 1666464484
transform 1 0 22356 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_234
timestamp 1666464484
transform 1 0 22632 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_244
timestamp 1666464484
transform 1 0 23552 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_250
timestamp 1666464484
transform 1 0 24104 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_253
timestamp 1666464484
transform 1 0 24380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_257
timestamp 1666464484
transform 1 0 24748 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_262
timestamp 1666464484
transform 1 0 25208 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_272
timestamp 1666464484
transform 1 0 26128 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_281
timestamp 1666464484
transform 1 0 26956 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_287
timestamp 1666464484
transform 1 0 27508 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_292
timestamp 1666464484
transform 1 0 27968 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_298
timestamp 1666464484
transform 1 0 28520 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1666464484
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1666464484
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_309
timestamp 1666464484
transform 1 0 29532 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_313
timestamp 1666464484
transform 1 0 29900 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_321
timestamp 1666464484
transform 1 0 30636 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_324
timestamp 1666464484
transform 1 0 30912 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_334
timestamp 1666464484
transform 1 0 31832 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_341
timestamp 1666464484
transform 1 0 32476 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_347
timestamp 1666464484
transform 1 0 33028 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_350
timestamp 1666464484
transform 1 0 33304 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_356
timestamp 1666464484
transform 1 0 33856 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_362
timestamp 1666464484
transform 1 0 34408 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_365
timestamp 1666464484
transform 1 0 34684 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_371
timestamp 1666464484
transform 1 0 35236 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_374
timestamp 1666464484
transform 1 0 35512 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_381
timestamp 1666464484
transform 1 0 36156 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_388
timestamp 1666464484
transform 1 0 36800 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_394
timestamp 1666464484
transform 1 0 37352 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_401
timestamp 1666464484
transform 1 0 37996 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_409
timestamp 1666464484
transform 1 0 38732 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_412
timestamp 1666464484
transform 1 0 39008 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_418
timestamp 1666464484
transform 1 0 39560 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_421
timestamp 1666464484
transform 1 0 39836 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_426
timestamp 1666464484
transform 1 0 40296 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_434
timestamp 1666464484
transform 1 0 41032 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_441
timestamp 1666464484
transform 1 0 41676 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_447
timestamp 1666464484
transform 1 0 42228 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_452
timestamp 1666464484
transform 1 0 42688 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_463
timestamp 1666464484
transform 1 0 43700 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_470
timestamp 1666464484
transform 1 0 44344 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_62_477
timestamp 1666464484
transform 1 0 44988 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_482
timestamp 1666464484
transform 1 0 45448 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_488
timestamp 1666464484
transform 1 0 46000 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_494
timestamp 1666464484
transform 1 0 46552 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_501
timestamp 1666464484
transform 1 0 47196 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_509
timestamp 1666464484
transform 1 0 47932 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_512
timestamp 1666464484
transform 1 0 48208 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_520
timestamp 1666464484
transform 1 0 48944 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_527
timestamp 1666464484
transform 1 0 49588 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1666464484
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_533
timestamp 1666464484
transform 1 0 50140 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_537
timestamp 1666464484
transform 1 0 50508 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_541
timestamp 1666464484
transform 1 0 50876 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_549
timestamp 1666464484
transform 1 0 51612 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_556
timestamp 1666464484
transform 1 0 52256 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_564
timestamp 1666464484
transform 1 0 52992 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_572
timestamp 1666464484
transform 1 0 53728 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_578
timestamp 1666464484
transform 1 0 54280 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_582
timestamp 1666464484
transform 1 0 54648 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_585
timestamp 1666464484
transform 1 0 54924 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_589
timestamp 1666464484
transform 1 0 55292 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_593
timestamp 1666464484
transform 1 0 55660 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_596
timestamp 1666464484
transform 1 0 55936 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_602
timestamp 1666464484
transform 1 0 56488 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_610
timestamp 1666464484
transform 1 0 57224 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_62_621
timestamp 1666464484
transform 1 0 58236 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_631
timestamp 1666464484
transform 1 0 59156 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_639
timestamp 1666464484
transform 1 0 59892 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_643
timestamp 1666464484
transform 1 0 60260 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_645
timestamp 1666464484
transform 1 0 60444 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_650
timestamp 1666464484
transform 1 0 60904 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_654
timestamp 1666464484
transform 1 0 61272 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_661
timestamp 1666464484
transform 1 0 61916 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_667
timestamp 1666464484
transform 1 0 62468 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_672
timestamp 1666464484
transform 1 0 62928 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_684
timestamp 1666464484
transform 1 0 64032 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_692
timestamp 1666464484
transform 1 0 64768 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_698
timestamp 1666464484
transform 1 0 65320 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_701
timestamp 1666464484
transform 1 0 65596 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_707
timestamp 1666464484
transform 1 0 66148 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_715
timestamp 1666464484
transform 1 0 66884 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_718
timestamp 1666464484
transform 1 0 67160 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_724
timestamp 1666464484
transform 1 0 67712 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_732
timestamp 1666464484
transform 1 0 68448 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_741
timestamp 1666464484
transform 1 0 69276 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_747
timestamp 1666464484
transform 1 0 69828 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_751
timestamp 1666464484
transform 1 0 70196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_754
timestamp 1666464484
transform 1 0 70472 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_757
timestamp 1666464484
transform 1 0 70748 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_761
timestamp 1666464484
transform 1 0 71116 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_773
timestamp 1666464484
transform 1 0 72220 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_778
timestamp 1666464484
transform 1 0 72680 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_790
timestamp 1666464484
transform 1 0 73784 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_794
timestamp 1666464484
transform 1 0 74152 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_801
timestamp 1666464484
transform 1 0 74796 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_807
timestamp 1666464484
transform 1 0 75348 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_811
timestamp 1666464484
transform 1 0 75716 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_813
timestamp 1666464484
transform 1 0 75900 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_818
timestamp 1666464484
transform 1 0 76360 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_826
timestamp 1666464484
transform 1 0 77096 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_830
timestamp 1666464484
transform 1 0 77464 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_836
timestamp 1666464484
transform 1 0 78016 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_844
timestamp 1666464484
transform 1 0 78752 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_850
timestamp 1666464484
transform 1 0 79304 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_62_862
timestamp 1666464484
transform 1 0 80408 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_62_869
timestamp 1666464484
transform 1 0 81052 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_880
timestamp 1666464484
transform 1 0 82064 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_886
timestamp 1666464484
transform 1 0 82616 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_892
timestamp 1666464484
transform 1 0 83168 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_898
timestamp 1666464484
transform 1 0 83720 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_904
timestamp 1666464484
transform 1 0 84272 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_910
timestamp 1666464484
transform 1 0 84824 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_914
timestamp 1666464484
transform 1 0 85192 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_917
timestamp 1666464484
transform 1 0 85468 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_923
timestamp 1666464484
transform 1 0 86020 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_925
timestamp 1666464484
transform 1 0 86204 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_929
timestamp 1666464484
transform 1 0 86572 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_941
timestamp 1666464484
transform 1 0 87676 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_953
timestamp 1666464484
transform 1 0 88780 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_958
timestamp 1666464484
transform 1 0 89240 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_964
timestamp 1666464484
transform 1 0 89792 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_970
timestamp 1666464484
transform 1 0 90344 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_976
timestamp 1666464484
transform 1 0 90896 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_981
timestamp 1666464484
transform 1 0 91356 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_993
timestamp 1666464484
transform 1 0 92460 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_999
timestamp 1666464484
transform 1 0 93012 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_1007
timestamp 1666464484
transform 1 0 93748 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_1011
timestamp 1666464484
transform 1 0 94116 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_1019
timestamp 1666464484
transform 1 0 94852 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1023
timestamp 1666464484
transform 1 0 95220 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_1026
timestamp 1666464484
transform 1 0 95496 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_1032
timestamp 1666464484
transform 1 0 96048 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1037
timestamp 1666464484
transform 1 0 96508 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_1049
timestamp 1666464484
transform 1 0 97612 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_1053
timestamp 1666464484
transform 1 0 97980 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1059
timestamp 1666464484
transform 1 0 98532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_1071
timestamp 1666464484
transform 1 0 99636 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_1079
timestamp 1666464484
transform 1 0 100372 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_1083
timestamp 1666464484
transform 1 0 100740 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1091
timestamp 1666464484
transform 1 0 101476 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1093
timestamp 1666464484
transform 1 0 101660 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1105
timestamp 1666464484
transform 1 0 102764 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_1108
timestamp 1666464484
transform 1 0 103040 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1114
timestamp 1666464484
transform 1 0 103592 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_1126
timestamp 1666464484
transform 1 0 104696 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_1131
timestamp 1666464484
transform 1 0 105156 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_1139
timestamp 1666464484
transform 1 0 105892 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_1145
timestamp 1666464484
transform 1 0 106444 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_1149
timestamp 1666464484
transform 1 0 106812 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_1153
timestamp 1666464484
transform 1 0 107180 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1159
timestamp 1666464484
transform 1 0 107732 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1171
timestamp 1666464484
transform 1 0 108836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_1183
timestamp 1666464484
transform 1 0 109940 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_1191
timestamp 1666464484
transform 1 0 110676 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_1195
timestamp 1666464484
transform 1 0 111044 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1203
timestamp 1666464484
transform 1 0 111780 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_1205
timestamp 1666464484
transform 1 0 111964 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_1209
timestamp 1666464484
transform 1 0 112332 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_1215
timestamp 1666464484
transform 1 0 112884 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_1223
timestamp 1666464484
transform 1 0 113620 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1227
timestamp 1666464484
transform 1 0 113988 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_1230
timestamp 1666464484
transform 1 0 114264 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_1236
timestamp 1666464484
transform 1 0 114816 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1240
timestamp 1666464484
transform 1 0 115184 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1243
timestamp 1666464484
transform 1 0 115460 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_1255
timestamp 1666464484
transform 1 0 116564 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1259
timestamp 1666464484
transform 1 0 116932 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_1261
timestamp 1666464484
transform 1 0 117116 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1271
timestamp 1666464484
transform 1 0 118036 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1283
timestamp 1666464484
transform 1 0 119140 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_1295
timestamp 1666464484
transform 1 0 120244 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_1305
timestamp 1666464484
transform 1 0 121164 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_1311
timestamp 1666464484
transform 1 0 121716 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1315
timestamp 1666464484
transform 1 0 122084 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_1317
timestamp 1666464484
transform 1 0 122268 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1327
timestamp 1666464484
transform 1 0 123188 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1339
timestamp 1666464484
transform 1 0 124292 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_1351
timestamp 1666464484
transform 1 0 125396 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_1359
timestamp 1666464484
transform 1 0 126132 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_1363
timestamp 1666464484
transform 1 0 126500 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1371
timestamp 1666464484
transform 1 0 127236 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1373
timestamp 1666464484
transform 1 0 127420 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1385
timestamp 1666464484
transform 1 0 128524 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1397
timestamp 1666464484
transform 1 0 129628 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1409
timestamp 1666464484
transform 1 0 130732 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_1421
timestamp 1666464484
transform 1 0 131836 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1427
timestamp 1666464484
transform 1 0 132388 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1429
timestamp 1666464484
transform 1 0 132572 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1441
timestamp 1666464484
transform 1 0 133676 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1453
timestamp 1666464484
transform 1 0 134780 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1465
timestamp 1666464484
transform 1 0 135884 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1468
timestamp 1666464484
transform 1 0 136160 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_1480
timestamp 1666464484
transform 1 0 137264 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_1485
timestamp 1666464484
transform 1 0 137724 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1489
timestamp 1666464484
transform 1 0 138092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1501
timestamp 1666464484
transform 1 0 139196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1513
timestamp 1666464484
transform 1 0 140300 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1525
timestamp 1666464484
transform 1 0 141404 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_1537
timestamp 1666464484
transform 1 0 142508 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_1541
timestamp 1666464484
transform 1 0 142876 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1551
timestamp 1666464484
transform 1 0 143796 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1563
timestamp 1666464484
transform 1 0 144900 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1575
timestamp 1666464484
transform 1 0 146004 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_1587
timestamp 1666464484
transform 1 0 147108 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1595
timestamp 1666464484
transform 1 0 147844 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_1597
timestamp 1666464484
transform 1 0 148028 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1666464484
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1666464484
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_27
timestamp 1666464484
transform 1 0 3588 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_32
timestamp 1666464484
transform 1 0 4048 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_38
timestamp 1666464484
transform 1 0 4600 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_50
timestamp 1666464484
transform 1 0 5704 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_57
timestamp 1666464484
transform 1 0 6348 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_62
timestamp 1666464484
transform 1 0 6808 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_68
timestamp 1666464484
transform 1 0 7360 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_76
timestamp 1666464484
transform 1 0 8096 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_80
timestamp 1666464484
transform 1 0 8464 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_86
timestamp 1666464484
transform 1 0 9016 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_97
timestamp 1666464484
transform 1 0 10028 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_103
timestamp 1666464484
transform 1 0 10580 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1666464484
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_113
timestamp 1666464484
transform 1 0 11500 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_121
timestamp 1666464484
transform 1 0 12236 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_124
timestamp 1666464484
transform 1 0 12512 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_136
timestamp 1666464484
transform 1 0 13616 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_141
timestamp 1666464484
transform 1 0 14076 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_147
timestamp 1666464484
transform 1 0 14628 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_159
timestamp 1666464484
transform 1 0 15732 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_164
timestamp 1666464484
transform 1 0 16192 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_169
timestamp 1666464484
transform 1 0 16652 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_175
timestamp 1666464484
transform 1 0 17204 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_179
timestamp 1666464484
transform 1 0 17572 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_185
timestamp 1666464484
transform 1 0 18124 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_191
timestamp 1666464484
transform 1 0 18676 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_198
timestamp 1666464484
transform 1 0 19320 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_205
timestamp 1666464484
transform 1 0 19964 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_211
timestamp 1666464484
transform 1 0 20516 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_215
timestamp 1666464484
transform 1 0 20884 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1666464484
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_225
timestamp 1666464484
transform 1 0 21804 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_231
timestamp 1666464484
transform 1 0 22356 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_237
timestamp 1666464484
transform 1 0 22908 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_244
timestamp 1666464484
transform 1 0 23552 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_257
timestamp 1666464484
transform 1 0 24748 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_264
timestamp 1666464484
transform 1 0 25392 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_272
timestamp 1666464484
transform 1 0 26128 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_278
timestamp 1666464484
transform 1 0 26680 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_281
timestamp 1666464484
transform 1 0 26956 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_287
timestamp 1666464484
transform 1 0 27508 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_297
timestamp 1666464484
transform 1 0 28428 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_305
timestamp 1666464484
transform 1 0 29164 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_311
timestamp 1666464484
transform 1 0 29716 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_317
timestamp 1666464484
transform 1 0 30268 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_322
timestamp 1666464484
transform 1 0 30728 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_328
timestamp 1666464484
transform 1 0 31280 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_334
timestamp 1666464484
transform 1 0 31832 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_337
timestamp 1666464484
transform 1 0 32108 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_342
timestamp 1666464484
transform 1 0 32568 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_352
timestamp 1666464484
transform 1 0 33488 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_361
timestamp 1666464484
transform 1 0 34316 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_369
timestamp 1666464484
transform 1 0 35052 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_374
timestamp 1666464484
transform 1 0 35512 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_382
timestamp 1666464484
transform 1 0 36248 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_390
timestamp 1666464484
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_393
timestamp 1666464484
transform 1 0 37260 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_403
timestamp 1666464484
transform 1 0 38180 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_411
timestamp 1666464484
transform 1 0 38916 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_422
timestamp 1666464484
transform 1 0 39928 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_426
timestamp 1666464484
transform 1 0 40296 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_430
timestamp 1666464484
transform 1 0 40664 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_438
timestamp 1666464484
transform 1 0 41400 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_446
timestamp 1666464484
transform 1 0 42136 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_449
timestamp 1666464484
transform 1 0 42412 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_460
timestamp 1666464484
transform 1 0 43424 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_468
timestamp 1666464484
transform 1 0 44160 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_476
timestamp 1666464484
transform 1 0 44896 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_483
timestamp 1666464484
transform 1 0 45540 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_487
timestamp 1666464484
transform 1 0 45908 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_492
timestamp 1666464484
transform 1 0 46368 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_498
timestamp 1666464484
transform 1 0 46920 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_502
timestamp 1666464484
transform 1 0 47288 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_505
timestamp 1666464484
transform 1 0 47564 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_516
timestamp 1666464484
transform 1 0 48576 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_524
timestamp 1666464484
transform 1 0 49312 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_532
timestamp 1666464484
transform 1 0 50048 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_537
timestamp 1666464484
transform 1 0 50508 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_543
timestamp 1666464484
transform 1 0 51060 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_550
timestamp 1666464484
transform 1 0 51704 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_558
timestamp 1666464484
transform 1 0 52440 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_561
timestamp 1666464484
transform 1 0 52716 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_565
timestamp 1666464484
transform 1 0 53084 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_573
timestamp 1666464484
transform 1 0 53820 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_581
timestamp 1666464484
transform 1 0 54556 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_588
timestamp 1666464484
transform 1 0 55200 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_596
timestamp 1666464484
transform 1 0 55936 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_603
timestamp 1666464484
transform 1 0 56580 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_611
timestamp 1666464484
transform 1 0 57316 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1666464484
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_617
timestamp 1666464484
transform 1 0 57868 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_628
timestamp 1666464484
transform 1 0 58880 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_632
timestamp 1666464484
transform 1 0 59248 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_637
timestamp 1666464484
transform 1 0 59708 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_645
timestamp 1666464484
transform 1 0 60444 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_653
timestamp 1666464484
transform 1 0 61180 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_663
timestamp 1666464484
transform 1 0 62100 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_670
timestamp 1666464484
transform 1 0 62744 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_673
timestamp 1666464484
transform 1 0 63020 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_678
timestamp 1666464484
transform 1 0 63480 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_691
timestamp 1666464484
transform 1 0 64676 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_704
timestamp 1666464484
transform 1 0 65872 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_712
timestamp 1666464484
transform 1 0 66608 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_721
timestamp 1666464484
transform 1 0 67436 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_727
timestamp 1666464484
transform 1 0 67988 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_729
timestamp 1666464484
transform 1 0 68172 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_733
timestamp 1666464484
transform 1 0 68540 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_738
timestamp 1666464484
transform 1 0 69000 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_746
timestamp 1666464484
transform 1 0 69736 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_754
timestamp 1666464484
transform 1 0 70472 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_761
timestamp 1666464484
transform 1 0 71116 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_765
timestamp 1666464484
transform 1 0 71484 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_768
timestamp 1666464484
transform 1 0 71760 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_774
timestamp 1666464484
transform 1 0 72312 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_781
timestamp 1666464484
transform 1 0 72956 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_785
timestamp 1666464484
transform 1 0 73324 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_789
timestamp 1666464484
transform 1 0 73692 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_795
timestamp 1666464484
transform 1 0 74244 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_802
timestamp 1666464484
transform 1 0 74888 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_812
timestamp 1666464484
transform 1 0 75808 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_822
timestamp 1666464484
transform 1 0 76728 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_828
timestamp 1666464484
transform 1 0 77280 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_834
timestamp 1666464484
transform 1 0 77832 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_841
timestamp 1666464484
transform 1 0 78476 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_847
timestamp 1666464484
transform 1 0 79028 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_853
timestamp 1666464484
transform 1 0 79580 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_863
timestamp 1666464484
transform 1 0 80500 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_876
timestamp 1666464484
transform 1 0 81696 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_884
timestamp 1666464484
transform 1 0 82432 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_892
timestamp 1666464484
transform 1 0 83168 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_897
timestamp 1666464484
transform 1 0 83628 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_903
timestamp 1666464484
transform 1 0 84180 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_915
timestamp 1666464484
transform 1 0 85284 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_921
timestamp 1666464484
transform 1 0 85836 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_929
timestamp 1666464484
transform 1 0 86572 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_935
timestamp 1666464484
transform 1 0 87124 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_941
timestamp 1666464484
transform 1 0 87676 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_947
timestamp 1666464484
transform 1 0 88228 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_951
timestamp 1666464484
transform 1 0 88596 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_953
timestamp 1666464484
transform 1 0 88780 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_957
timestamp 1666464484
transform 1 0 89148 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_962
timestamp 1666464484
transform 1 0 89608 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_968
timestamp 1666464484
transform 1 0 90160 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_973
timestamp 1666464484
transform 1 0 90620 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_979
timestamp 1666464484
transform 1 0 91172 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_985
timestamp 1666464484
transform 1 0 91724 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_991
timestamp 1666464484
transform 1 0 92276 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1003
timestamp 1666464484
transform 1 0 93380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1007
timestamp 1666464484
transform 1 0 93748 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_1009
timestamp 1666464484
transform 1 0 93932 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_1013
timestamp 1666464484
transform 1 0 94300 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1024
timestamp 1666464484
transform 1 0 95312 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1032
timestamp 1666464484
transform 1 0 96048 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1038
timestamp 1666464484
transform 1 0 96600 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_1044
timestamp 1666464484
transform 1 0 97152 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1054
timestamp 1666464484
transform 1 0 98072 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_1062
timestamp 1666464484
transform 1 0 98808 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_1065
timestamp 1666464484
transform 1 0 99084 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1069
timestamp 1666464484
transform 1 0 99452 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_1075
timestamp 1666464484
transform 1 0 100004 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1081
timestamp 1666464484
transform 1 0 100556 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1084
timestamp 1666464484
transform 1 0 100832 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_1092
timestamp 1666464484
transform 1 0 101568 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1098
timestamp 1666464484
transform 1 0 102120 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_1101
timestamp 1666464484
transform 1 0 102396 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1107
timestamp 1666464484
transform 1 0 102948 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1112
timestamp 1666464484
transform 1 0 103408 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_1118
timestamp 1666464484
transform 1 0 103960 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_1121
timestamp 1666464484
transform 1 0 104236 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_1125
timestamp 1666464484
transform 1 0 104604 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1137
timestamp 1666464484
transform 1 0 105708 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1145
timestamp 1666464484
transform 1 0 106444 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1152
timestamp 1666464484
transform 1 0 107088 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1158
timestamp 1666464484
transform 1 0 107640 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1164
timestamp 1666464484
transform 1 0 108192 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_1170
timestamp 1666464484
transform 1 0 108744 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_1177
timestamp 1666464484
transform 1 0 109388 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1181
timestamp 1666464484
transform 1 0 109756 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1185
timestamp 1666464484
transform 1 0 110124 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1188
timestamp 1666464484
transform 1 0 110400 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1195
timestamp 1666464484
transform 1 0 111044 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_1201
timestamp 1666464484
transform 1 0 111596 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1209
timestamp 1666464484
transform 1 0 112332 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1214
timestamp 1666464484
transform 1 0 112792 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1220
timestamp 1666464484
transform 1 0 113344 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1228
timestamp 1666464484
transform 1 0 114080 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1233
timestamp 1666464484
transform 1 0 114540 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1237
timestamp 1666464484
transform 1 0 114908 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1241
timestamp 1666464484
transform 1 0 115276 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1247
timestamp 1666464484
transform 1 0 115828 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_1253
timestamp 1666464484
transform 1 0 116380 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_63_1263
timestamp 1666464484
transform 1 0 117300 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1273
timestamp 1666464484
transform 1 0 118220 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1279
timestamp 1666464484
transform 1 0 118772 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_1285
timestamp 1666464484
transform 1 0 119324 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_1289
timestamp 1666464484
transform 1 0 119692 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_1293
timestamp 1666464484
transform 1 0 120060 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1301
timestamp 1666464484
transform 1 0 120796 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1304
timestamp 1666464484
transform 1 0 121072 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_1312
timestamp 1666464484
transform 1 0 121808 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1320
timestamp 1666464484
transform 1 0 122544 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1323
timestamp 1666464484
transform 1 0 122820 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1330
timestamp 1666464484
transform 1 0 123464 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1336
timestamp 1666464484
transform 1 0 124016 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_1342
timestamp 1666464484
transform 1 0 124568 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_1345
timestamp 1666464484
transform 1 0 124844 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1349
timestamp 1666464484
transform 1 0 125212 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_1355
timestamp 1666464484
transform 1 0 125764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1361
timestamp 1666464484
transform 1 0 126316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1366
timestamp 1666464484
transform 1 0 126776 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1372
timestamp 1666464484
transform 1 0 127328 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1378
timestamp 1666464484
transform 1 0 127880 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1384
timestamp 1666464484
transform 1 0 128432 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1388
timestamp 1666464484
transform 1 0 128800 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1391
timestamp 1666464484
transform 1 0 129076 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1395
timestamp 1666464484
transform 1 0 129444 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_1398
timestamp 1666464484
transform 1 0 129720 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_1401
timestamp 1666464484
transform 1 0 129996 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1407
timestamp 1666464484
transform 1 0 130548 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1413
timestamp 1666464484
transform 1 0 131100 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1419
timestamp 1666464484
transform 1 0 131652 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1426
timestamp 1666464484
transform 1 0 132296 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1432
timestamp 1666464484
transform 1 0 132848 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_1438
timestamp 1666464484
transform 1 0 133400 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_63_1448
timestamp 1666464484
transform 1 0 134320 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_63_1457
timestamp 1666464484
transform 1 0 135148 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1463
timestamp 1666464484
transform 1 0 135700 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1467
timestamp 1666464484
transform 1 0 136068 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_1473
timestamp 1666464484
transform 1 0 136620 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_1481
timestamp 1666464484
transform 1 0 137356 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1487
timestamp 1666464484
transform 1 0 137908 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_1493
timestamp 1666464484
transform 1 0 138460 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_1501
timestamp 1666464484
transform 1 0 139196 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_1506
timestamp 1666464484
transform 1 0 139656 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_1513
timestamp 1666464484
transform 1 0 140300 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_1517
timestamp 1666464484
transform 1 0 140668 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1528
timestamp 1666464484
transform 1 0 141680 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1534
timestamp 1666464484
transform 1 0 142232 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_1540
timestamp 1666464484
transform 1 0 142784 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1548
timestamp 1666464484
transform 1 0 143520 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1552
timestamp 1666464484
transform 1 0 143888 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_1558
timestamp 1666464484
transform 1 0 144440 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_1566
timestamp 1666464484
transform 1 0 145176 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_1569
timestamp 1666464484
transform 1 0 145452 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1575
timestamp 1666464484
transform 1 0 146004 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1579
timestamp 1666464484
transform 1 0 146372 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1585
timestamp 1666464484
transform 1 0 146924 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_1591
timestamp 1666464484
transform 1 0 147476 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1666464484
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_15
timestamp 1666464484
transform 1 0 2484 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_21
timestamp 1666464484
transform 1 0 3036 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1666464484
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_29
timestamp 1666464484
transform 1 0 3772 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_37
timestamp 1666464484
transform 1 0 4508 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_42
timestamp 1666464484
transform 1 0 4968 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_52
timestamp 1666464484
transform 1 0 5888 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_57
timestamp 1666464484
transform 1 0 6348 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_62
timestamp 1666464484
transform 1 0 6808 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_64_72
timestamp 1666464484
transform 1 0 7728 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_82
timestamp 1666464484
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_85
timestamp 1666464484
transform 1 0 8924 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_92
timestamp 1666464484
transform 1 0 9568 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_101
timestamp 1666464484
transform 1 0 10396 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_105
timestamp 1666464484
transform 1 0 10764 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_110
timestamp 1666464484
transform 1 0 11224 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_113
timestamp 1666464484
transform 1 0 11500 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_117
timestamp 1666464484
transform 1 0 11868 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_122
timestamp 1666464484
transform 1 0 12328 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_64_132
timestamp 1666464484
transform 1 0 13248 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_64_141
timestamp 1666464484
transform 1 0 14076 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_147
timestamp 1666464484
transform 1 0 14628 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_152
timestamp 1666464484
transform 1 0 15088 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_64_162
timestamp 1666464484
transform 1 0 16008 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1666464484
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_175
timestamp 1666464484
transform 1 0 17204 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_182
timestamp 1666464484
transform 1 0 17848 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_192
timestamp 1666464484
transform 1 0 18768 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1666464484
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_203
timestamp 1666464484
transform 1 0 19780 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_207
timestamp 1666464484
transform 1 0 20148 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_212
timestamp 1666464484
transform 1 0 20608 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_222
timestamp 1666464484
transform 1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_225
timestamp 1666464484
transform 1 0 21804 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_232
timestamp 1666464484
transform 1 0 22448 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_242
timestamp 1666464484
transform 1 0 23368 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_246
timestamp 1666464484
transform 1 0 23736 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_250
timestamp 1666464484
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1666464484
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_264
timestamp 1666464484
transform 1 0 25392 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_270
timestamp 1666464484
transform 1 0 25944 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_278
timestamp 1666464484
transform 1 0 26680 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1666464484
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_286
timestamp 1666464484
transform 1 0 27416 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_299
timestamp 1666464484
transform 1 0 28612 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_306
timestamp 1666464484
transform 1 0 29256 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1666464484
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_315
timestamp 1666464484
transform 1 0 30084 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_319
timestamp 1666464484
transform 1 0 30452 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_324
timestamp 1666464484
transform 1 0 30912 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_332
timestamp 1666464484
transform 1 0 31648 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1666464484
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_343
timestamp 1666464484
transform 1 0 32660 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_349
timestamp 1666464484
transform 1 0 33212 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_354
timestamp 1666464484
transform 1 0 33672 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_362
timestamp 1666464484
transform 1 0 34408 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_365
timestamp 1666464484
transform 1 0 34684 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_377
timestamp 1666464484
transform 1 0 35788 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_390
timestamp 1666464484
transform 1 0 36984 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_393
timestamp 1666464484
transform 1 0 37260 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_399
timestamp 1666464484
transform 1 0 37812 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_409
timestamp 1666464484
transform 1 0 38732 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_417
timestamp 1666464484
transform 1 0 39468 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_421
timestamp 1666464484
transform 1 0 39836 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_427
timestamp 1666464484
transform 1 0 40388 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_440
timestamp 1666464484
transform 1 0 41584 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_446
timestamp 1666464484
transform 1 0 42136 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_449
timestamp 1666464484
transform 1 0 42412 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_453
timestamp 1666464484
transform 1 0 42780 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_463
timestamp 1666464484
transform 1 0 43700 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_469
timestamp 1666464484
transform 1 0 44252 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_474
timestamp 1666464484
transform 1 0 44712 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_477
timestamp 1666464484
transform 1 0 44988 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_483
timestamp 1666464484
transform 1 0 45540 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_491
timestamp 1666464484
transform 1 0 46276 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_497
timestamp 1666464484
transform 1 0 46828 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_502
timestamp 1666464484
transform 1 0 47288 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_505
timestamp 1666464484
transform 1 0 47564 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_517
timestamp 1666464484
transform 1 0 48668 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_525
timestamp 1666464484
transform 1 0 49404 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_530
timestamp 1666464484
transform 1 0 49864 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_533
timestamp 1666464484
transform 1 0 50140 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_537
timestamp 1666464484
transform 1 0 50508 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_545
timestamp 1666464484
transform 1 0 51244 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_558
timestamp 1666464484
transform 1 0 52440 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_561
timestamp 1666464484
transform 1 0 52716 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_572
timestamp 1666464484
transform 1 0 53728 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_578
timestamp 1666464484
transform 1 0 54280 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_586
timestamp 1666464484
transform 1 0 55016 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_589
timestamp 1666464484
transform 1 0 55292 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_593
timestamp 1666464484
transform 1 0 55660 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_601
timestamp 1666464484
transform 1 0 56396 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_614
timestamp 1666464484
transform 1 0 57592 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_617
timestamp 1666464484
transform 1 0 57868 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_628
timestamp 1666464484
transform 1 0 58880 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_634
timestamp 1666464484
transform 1 0 59432 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_642
timestamp 1666464484
transform 1 0 60168 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_645
timestamp 1666464484
transform 1 0 60444 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_658
timestamp 1666464484
transform 1 0 61640 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_667
timestamp 1666464484
transform 1 0 62468 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_671
timestamp 1666464484
transform 1 0 62836 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_673
timestamp 1666464484
transform 1 0 63020 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_684
timestamp 1666464484
transform 1 0 64032 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_697
timestamp 1666464484
transform 1 0 65228 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_701
timestamp 1666464484
transform 1 0 65596 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_64_716
timestamp 1666464484
transform 1 0 66976 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_726
timestamp 1666464484
transform 1 0 67896 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_729
timestamp 1666464484
transform 1 0 68172 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_740
timestamp 1666464484
transform 1 0 69184 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_752
timestamp 1666464484
transform 1 0 70288 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_757
timestamp 1666464484
transform 1 0 70748 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_768
timestamp 1666464484
transform 1 0 71760 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_776
timestamp 1666464484
transform 1 0 72496 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_782
timestamp 1666464484
transform 1 0 73048 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_785
timestamp 1666464484
transform 1 0 73324 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_792
timestamp 1666464484
transform 1 0 73968 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_800
timestamp 1666464484
transform 1 0 74704 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_810
timestamp 1666464484
transform 1 0 75624 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_813
timestamp 1666464484
transform 1 0 75900 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_817
timestamp 1666464484
transform 1 0 76268 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_827
timestamp 1666464484
transform 1 0 77188 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_835
timestamp 1666464484
transform 1 0 77924 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_839
timestamp 1666464484
transform 1 0 78292 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_841
timestamp 1666464484
transform 1 0 78476 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_856
timestamp 1666464484
transform 1 0 79856 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_864
timestamp 1666464484
transform 1 0 80592 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_869
timestamp 1666464484
transform 1 0 81052 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_880
timestamp 1666464484
transform 1 0 82064 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_893
timestamp 1666464484
transform 1 0 83260 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_897
timestamp 1666464484
transform 1 0 83628 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_903
timestamp 1666464484
transform 1 0 84180 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_911
timestamp 1666464484
transform 1 0 84916 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_919
timestamp 1666464484
transform 1 0 85652 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_923
timestamp 1666464484
transform 1 0 86020 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_925
timestamp 1666464484
transform 1 0 86204 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_931
timestamp 1666464484
transform 1 0 86756 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_939
timestamp 1666464484
transform 1 0 87492 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_947
timestamp 1666464484
transform 1 0 88228 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_951
timestamp 1666464484
transform 1 0 88596 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_953
timestamp 1666464484
transform 1 0 88780 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_959
timestamp 1666464484
transform 1 0 89332 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_967
timestamp 1666464484
transform 1 0 90068 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_975
timestamp 1666464484
transform 1 0 90804 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_979
timestamp 1666464484
transform 1 0 91172 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_981
timestamp 1666464484
transform 1 0 91356 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_987
timestamp 1666464484
transform 1 0 91908 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_995
timestamp 1666464484
transform 1 0 92644 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1003
timestamp 1666464484
transform 1 0 93380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1007
timestamp 1666464484
transform 1 0 93748 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_1009
timestamp 1666464484
transform 1 0 93932 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1015
timestamp 1666464484
transform 1 0 94484 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1023
timestamp 1666464484
transform 1 0 95220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1031
timestamp 1666464484
transform 1 0 95956 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1035
timestamp 1666464484
transform 1 0 96324 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_1037
timestamp 1666464484
transform 1 0 96508 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1043
timestamp 1666464484
transform 1 0 97060 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1051
timestamp 1666464484
transform 1 0 97796 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1059
timestamp 1666464484
transform 1 0 98532 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1063
timestamp 1666464484
transform 1 0 98900 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_1065
timestamp 1666464484
transform 1 0 99084 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1071
timestamp 1666464484
transform 1 0 99636 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1079
timestamp 1666464484
transform 1 0 100372 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1087
timestamp 1666464484
transform 1 0 101108 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1091
timestamp 1666464484
transform 1 0 101476 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_1093
timestamp 1666464484
transform 1 0 101660 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1099
timestamp 1666464484
transform 1 0 102212 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1107
timestamp 1666464484
transform 1 0 102948 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1115
timestamp 1666464484
transform 1 0 103684 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1119
timestamp 1666464484
transform 1 0 104052 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_1121
timestamp 1666464484
transform 1 0 104236 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1127
timestamp 1666464484
transform 1 0 104788 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1135
timestamp 1666464484
transform 1 0 105524 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1143
timestamp 1666464484
transform 1 0 106260 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1147
timestamp 1666464484
transform 1 0 106628 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_1149
timestamp 1666464484
transform 1 0 106812 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1155
timestamp 1666464484
transform 1 0 107364 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1163
timestamp 1666464484
transform 1 0 108100 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1167
timestamp 1666464484
transform 1 0 108468 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1172
timestamp 1666464484
transform 1 0 108928 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_1177
timestamp 1666464484
transform 1 0 109388 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1183
timestamp 1666464484
transform 1 0 109940 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1191
timestamp 1666464484
transform 1 0 110676 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1199
timestamp 1666464484
transform 1 0 111412 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1203
timestamp 1666464484
transform 1 0 111780 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_1205
timestamp 1666464484
transform 1 0 111964 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1211
timestamp 1666464484
transform 1 0 112516 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1219
timestamp 1666464484
transform 1 0 113252 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1227
timestamp 1666464484
transform 1 0 113988 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1231
timestamp 1666464484
transform 1 0 114356 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_1233
timestamp 1666464484
transform 1 0 114540 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1239
timestamp 1666464484
transform 1 0 115092 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1247
timestamp 1666464484
transform 1 0 115828 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1255
timestamp 1666464484
transform 1 0 116564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1259
timestamp 1666464484
transform 1 0 116932 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_1261
timestamp 1666464484
transform 1 0 117116 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1267
timestamp 1666464484
transform 1 0 117668 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1275
timestamp 1666464484
transform 1 0 118404 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1283
timestamp 1666464484
transform 1 0 119140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1287
timestamp 1666464484
transform 1 0 119508 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_1289
timestamp 1666464484
transform 1 0 119692 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1295
timestamp 1666464484
transform 1 0 120244 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1303
timestamp 1666464484
transform 1 0 120980 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1311
timestamp 1666464484
transform 1 0 121716 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1315
timestamp 1666464484
transform 1 0 122084 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_1317
timestamp 1666464484
transform 1 0 122268 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1323
timestamp 1666464484
transform 1 0 122820 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1331
timestamp 1666464484
transform 1 0 123556 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1339
timestamp 1666464484
transform 1 0 124292 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1343
timestamp 1666464484
transform 1 0 124660 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_1345
timestamp 1666464484
transform 1 0 124844 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1351
timestamp 1666464484
transform 1 0 125396 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1359
timestamp 1666464484
transform 1 0 126132 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1367
timestamp 1666464484
transform 1 0 126868 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1371
timestamp 1666464484
transform 1 0 127236 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_1373
timestamp 1666464484
transform 1 0 127420 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1379
timestamp 1666464484
transform 1 0 127972 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1387
timestamp 1666464484
transform 1 0 128708 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1395
timestamp 1666464484
transform 1 0 129444 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1399
timestamp 1666464484
transform 1 0 129812 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_1401
timestamp 1666464484
transform 1 0 129996 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1407
timestamp 1666464484
transform 1 0 130548 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1415
timestamp 1666464484
transform 1 0 131284 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1423
timestamp 1666464484
transform 1 0 132020 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1427
timestamp 1666464484
transform 1 0 132388 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_1429
timestamp 1666464484
transform 1 0 132572 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1435
timestamp 1666464484
transform 1 0 133124 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1443
timestamp 1666464484
transform 1 0 133860 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1447
timestamp 1666464484
transform 1 0 134228 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1452
timestamp 1666464484
transform 1 0 134688 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_1457
timestamp 1666464484
transform 1 0 135148 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1463
timestamp 1666464484
transform 1 0 135700 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1467
timestamp 1666464484
transform 1 0 136068 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_1472
timestamp 1666464484
transform 1 0 136528 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_1482
timestamp 1666464484
transform 1 0 137448 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_1485
timestamp 1666464484
transform 1 0 137724 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_1492
timestamp 1666464484
transform 1 0 138368 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1502
timestamp 1666464484
transform 1 0 139288 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_1509
timestamp 1666464484
transform 1 0 139932 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_1513
timestamp 1666464484
transform 1 0 140300 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1519
timestamp 1666464484
transform 1 0 140852 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1527
timestamp 1666464484
transform 1 0 141588 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1535
timestamp 1666464484
transform 1 0 142324 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1539
timestamp 1666464484
transform 1 0 142692 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_1541
timestamp 1666464484
transform 1 0 142876 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1547
timestamp 1666464484
transform 1 0 143428 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1555
timestamp 1666464484
transform 1 0 144164 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1563
timestamp 1666464484
transform 1 0 144900 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1567
timestamp 1666464484
transform 1 0 145268 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_1569
timestamp 1666464484
transform 1 0 145452 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1575
timestamp 1666464484
transform 1 0 146004 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1583
timestamp 1666464484
transform 1 0 146740 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1587
timestamp 1666464484
transform 1 0 147108 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1592
timestamp 1666464484
transform 1 0 147568 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_1597
timestamp 1666464484
transform 1 0 148028 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 148856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 148856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 148856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 148856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 148856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 148856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 148856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 148856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 148856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 148856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 148856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 148856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 148856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 148856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 148856 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 148856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 148856 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 148856 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 148856 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 148856 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 148856 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 148856 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 148856 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 148856 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 148856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 148856 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 148856 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 148856 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666464484
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666464484
transform -1 0 148856 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666464484
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666464484
transform -1 0 148856 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666464484
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666464484
transform -1 0 148856 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666464484
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666464484
transform -1 0 148856 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666464484
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666464484
transform -1 0 148856 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666464484
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666464484
transform -1 0 148856 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666464484
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666464484
transform -1 0 148856 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666464484
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666464484
transform -1 0 148856 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666464484
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666464484
transform -1 0 148856 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666464484
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666464484
transform -1 0 148856 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666464484
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666464484
transform -1 0 148856 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666464484
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666464484
transform -1 0 148856 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666464484
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666464484
transform -1 0 148856 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666464484
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666464484
transform -1 0 148856 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666464484
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666464484
transform -1 0 148856 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666464484
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666464484
transform -1 0 148856 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666464484
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666464484
transform -1 0 148856 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1666464484
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1666464484
transform -1 0 148856 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1666464484
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1666464484
transform -1 0 148856 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1666464484
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1666464484
transform -1 0 148856 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1666464484
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1666464484
transform -1 0 148856 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1666464484
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1666464484
transform -1 0 148856 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1666464484
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1666464484
transform -1 0 148856 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1666464484
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1666464484
transform -1 0 148856 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1666464484
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1666464484
transform -1 0 148856 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1666464484
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1666464484
transform -1 0 148856 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1666464484
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1666464484
transform -1 0 148856 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1666464484
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1666464484
transform -1 0 148856 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1666464484
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1666464484
transform -1 0 148856 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1666464484
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1666464484
transform -1 0 148856 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1666464484
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1666464484
transform -1 0 148856 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1666464484
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1666464484
transform -1 0 148856 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1666464484
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1666464484
transform -1 0 148856 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1666464484
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1666464484
transform -1 0 148856 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1666464484
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1666464484
transform -1 0 148856 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1666464484
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1666464484
transform -1 0 148856 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1666464484
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1666464484
transform -1 0 148856 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1666464484
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1666464484
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1666464484
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1666464484
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1666464484
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1666464484
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1666464484
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1666464484
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1666464484
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1666464484
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1666464484
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1666464484
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1666464484
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1666464484
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1666464484
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1666464484
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1666464484
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1666464484
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1666464484
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1666464484
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1666464484
transform 1 0 70656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1666464484
transform 1 0 73232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1666464484
transform 1 0 75808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1666464484
transform 1 0 78384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1666464484
transform 1 0 80960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1666464484
transform 1 0 83536 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1666464484
transform 1 0 86112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1666464484
transform 1 0 88688 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1666464484
transform 1 0 91264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1666464484
transform 1 0 93840 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1666464484
transform 1 0 96416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1666464484
transform 1 0 98992 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1666464484
transform 1 0 101568 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1666464484
transform 1 0 104144 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1666464484
transform 1 0 106720 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1666464484
transform 1 0 109296 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1666464484
transform 1 0 111872 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1666464484
transform 1 0 114448 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1666464484
transform 1 0 117024 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1666464484
transform 1 0 119600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1666464484
transform 1 0 122176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1666464484
transform 1 0 124752 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1666464484
transform 1 0 127328 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1666464484
transform 1 0 129904 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1666464484
transform 1 0 132480 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1666464484
transform 1 0 135056 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1666464484
transform 1 0 137632 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1666464484
transform 1 0 140208 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1666464484
transform 1 0 142784 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1666464484
transform 1 0 145360 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1666464484
transform 1 0 147936 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1666464484
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1666464484
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1666464484
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1666464484
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1666464484
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1666464484
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1666464484
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1666464484
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1666464484
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1666464484
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1666464484
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1666464484
transform 1 0 78384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1666464484
transform 1 0 83536 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1666464484
transform 1 0 88688 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1666464484
transform 1 0 93840 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666464484
transform 1 0 98992 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666464484
transform 1 0 104144 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666464484
transform 1 0 109296 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666464484
transform 1 0 114448 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666464484
transform 1 0 119600 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666464484
transform 1 0 124752 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666464484
transform 1 0 129904 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666464484
transform 1 0 135056 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666464484
transform 1 0 140208 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666464484
transform 1 0 145360 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666464484
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666464484
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666464484
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666464484
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666464484
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666464484
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666464484
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666464484
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666464484
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666464484
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666464484
transform 1 0 70656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666464484
transform 1 0 75808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666464484
transform 1 0 80960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666464484
transform 1 0 86112 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666464484
transform 1 0 91264 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666464484
transform 1 0 96416 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666464484
transform 1 0 101568 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666464484
transform 1 0 106720 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666464484
transform 1 0 111872 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666464484
transform 1 0 117024 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666464484
transform 1 0 122176 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666464484
transform 1 0 127328 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666464484
transform 1 0 132480 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666464484
transform 1 0 137632 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666464484
transform 1 0 142784 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666464484
transform 1 0 147936 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666464484
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666464484
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666464484
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666464484
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666464484
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666464484
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666464484
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666464484
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666464484
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666464484
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666464484
transform 1 0 73232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666464484
transform 1 0 78384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666464484
transform 1 0 83536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666464484
transform 1 0 88688 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666464484
transform 1 0 93840 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666464484
transform 1 0 98992 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666464484
transform 1 0 104144 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666464484
transform 1 0 109296 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666464484
transform 1 0 114448 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666464484
transform 1 0 119600 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666464484
transform 1 0 124752 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666464484
transform 1 0 129904 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666464484
transform 1 0 135056 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666464484
transform 1 0 140208 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666464484
transform 1 0 145360 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666464484
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666464484
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666464484
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666464484
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666464484
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666464484
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666464484
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666464484
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666464484
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666464484
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666464484
transform 1 0 70656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666464484
transform 1 0 75808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666464484
transform 1 0 80960 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666464484
transform 1 0 86112 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666464484
transform 1 0 91264 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1666464484
transform 1 0 96416 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1666464484
transform 1 0 101568 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1666464484
transform 1 0 106720 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1666464484
transform 1 0 111872 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1666464484
transform 1 0 117024 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1666464484
transform 1 0 122176 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1666464484
transform 1 0 127328 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1666464484
transform 1 0 132480 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1666464484
transform 1 0 137632 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1666464484
transform 1 0 142784 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1666464484
transform 1 0 147936 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1666464484
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1666464484
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1666464484
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1666464484
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1666464484
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1666464484
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1666464484
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1666464484
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1666464484
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1666464484
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1666464484
transform 1 0 73232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1666464484
transform 1 0 78384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1666464484
transform 1 0 83536 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1666464484
transform 1 0 88688 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1666464484
transform 1 0 93840 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1666464484
transform 1 0 98992 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1666464484
transform 1 0 104144 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1666464484
transform 1 0 109296 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1666464484
transform 1 0 114448 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1666464484
transform 1 0 119600 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1666464484
transform 1 0 124752 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1666464484
transform 1 0 129904 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1666464484
transform 1 0 135056 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1666464484
transform 1 0 140208 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1666464484
transform 1 0 145360 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1666464484
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1666464484
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1666464484
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1666464484
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1666464484
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1666464484
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1666464484
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1666464484
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1666464484
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1666464484
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1666464484
transform 1 0 70656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1666464484
transform 1 0 75808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1666464484
transform 1 0 80960 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1666464484
transform 1 0 86112 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1666464484
transform 1 0 91264 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1666464484
transform 1 0 96416 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1666464484
transform 1 0 101568 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1666464484
transform 1 0 106720 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1666464484
transform 1 0 111872 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1666464484
transform 1 0 117024 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1666464484
transform 1 0 122176 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1666464484
transform 1 0 127328 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1666464484
transform 1 0 132480 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1666464484
transform 1 0 137632 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1666464484
transform 1 0 142784 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1666464484
transform 1 0 147936 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1666464484
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1666464484
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1666464484
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1666464484
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1666464484
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1666464484
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1666464484
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1666464484
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1666464484
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1666464484
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1666464484
transform 1 0 73232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1666464484
transform 1 0 78384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1666464484
transform 1 0 83536 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1666464484
transform 1 0 88688 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1666464484
transform 1 0 93840 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1666464484
transform 1 0 98992 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1666464484
transform 1 0 104144 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1666464484
transform 1 0 109296 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1666464484
transform 1 0 114448 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1666464484
transform 1 0 119600 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1666464484
transform 1 0 124752 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1666464484
transform 1 0 129904 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1666464484
transform 1 0 135056 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1666464484
transform 1 0 140208 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1666464484
transform 1 0 145360 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1666464484
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1666464484
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1666464484
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1666464484
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1666464484
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1666464484
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1666464484
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1666464484
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1666464484
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1666464484
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1666464484
transform 1 0 70656 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1666464484
transform 1 0 75808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1666464484
transform 1 0 80960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1666464484
transform 1 0 86112 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1666464484
transform 1 0 91264 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1666464484
transform 1 0 96416 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1666464484
transform 1 0 101568 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1666464484
transform 1 0 106720 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1666464484
transform 1 0 111872 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1666464484
transform 1 0 117024 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1666464484
transform 1 0 122176 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1666464484
transform 1 0 127328 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1666464484
transform 1 0 132480 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1666464484
transform 1 0 137632 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1666464484
transform 1 0 142784 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1666464484
transform 1 0 147936 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1666464484
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1666464484
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1666464484
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1666464484
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1666464484
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1666464484
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1666464484
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1666464484
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1666464484
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1666464484
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1666464484
transform 1 0 73232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1666464484
transform 1 0 78384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1666464484
transform 1 0 83536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1666464484
transform 1 0 88688 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1666464484
transform 1 0 93840 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1666464484
transform 1 0 98992 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1666464484
transform 1 0 104144 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1666464484
transform 1 0 109296 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1666464484
transform 1 0 114448 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1666464484
transform 1 0 119600 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1666464484
transform 1 0 124752 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1666464484
transform 1 0 129904 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1666464484
transform 1 0 135056 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1666464484
transform 1 0 140208 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1666464484
transform 1 0 145360 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1666464484
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1666464484
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1666464484
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1666464484
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1666464484
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1666464484
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1666464484
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1666464484
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1666464484
transform 1 0 60352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1666464484
transform 1 0 65504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1666464484
transform 1 0 70656 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1666464484
transform 1 0 75808 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1666464484
transform 1 0 80960 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1666464484
transform 1 0 86112 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1666464484
transform 1 0 91264 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1666464484
transform 1 0 96416 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1666464484
transform 1 0 101568 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1666464484
transform 1 0 106720 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1666464484
transform 1 0 111872 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1666464484
transform 1 0 117024 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1666464484
transform 1 0 122176 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1666464484
transform 1 0 127328 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1666464484
transform 1 0 132480 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1666464484
transform 1 0 137632 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1666464484
transform 1 0 142784 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1666464484
transform 1 0 147936 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1666464484
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1666464484
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1666464484
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1666464484
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1666464484
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1666464484
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1666464484
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1666464484
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1666464484
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1666464484
transform 1 0 62928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1666464484
transform 1 0 68080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1666464484
transform 1 0 73232 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1666464484
transform 1 0 78384 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1666464484
transform 1 0 83536 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1666464484
transform 1 0 88688 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1666464484
transform 1 0 93840 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1666464484
transform 1 0 98992 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1666464484
transform 1 0 104144 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1666464484
transform 1 0 109296 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1666464484
transform 1 0 114448 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1666464484
transform 1 0 119600 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1666464484
transform 1 0 124752 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1666464484
transform 1 0 129904 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1666464484
transform 1 0 135056 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1666464484
transform 1 0 140208 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1666464484
transform 1 0 145360 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1666464484
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1666464484
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1666464484
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1666464484
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1666464484
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1666464484
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1666464484
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1666464484
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1666464484
transform 1 0 60352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1666464484
transform 1 0 65504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1666464484
transform 1 0 70656 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1666464484
transform 1 0 75808 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1666464484
transform 1 0 80960 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1666464484
transform 1 0 86112 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1666464484
transform 1 0 91264 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1666464484
transform 1 0 96416 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1666464484
transform 1 0 101568 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1666464484
transform 1 0 106720 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1666464484
transform 1 0 111872 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1666464484
transform 1 0 117024 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1666464484
transform 1 0 122176 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1666464484
transform 1 0 127328 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1666464484
transform 1 0 132480 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1666464484
transform 1 0 137632 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1666464484
transform 1 0 142784 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1666464484
transform 1 0 147936 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1666464484
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1666464484
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1666464484
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1666464484
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1666464484
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1666464484
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1666464484
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1666464484
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1666464484
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1666464484
transform 1 0 62928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1666464484
transform 1 0 68080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1666464484
transform 1 0 73232 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1666464484
transform 1 0 78384 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1666464484
transform 1 0 83536 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1666464484
transform 1 0 88688 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1666464484
transform 1 0 93840 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1666464484
transform 1 0 98992 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1666464484
transform 1 0 104144 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1666464484
transform 1 0 109296 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1666464484
transform 1 0 114448 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1666464484
transform 1 0 119600 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1666464484
transform 1 0 124752 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1666464484
transform 1 0 129904 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1666464484
transform 1 0 135056 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1666464484
transform 1 0 140208 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1666464484
transform 1 0 145360 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1666464484
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1666464484
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1666464484
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1666464484
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1666464484
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1666464484
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1666464484
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1666464484
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1666464484
transform 1 0 60352 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1666464484
transform 1 0 65504 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1666464484
transform 1 0 70656 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1666464484
transform 1 0 75808 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1666464484
transform 1 0 80960 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1666464484
transform 1 0 86112 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1666464484
transform 1 0 91264 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1666464484
transform 1 0 96416 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1666464484
transform 1 0 101568 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1666464484
transform 1 0 106720 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1666464484
transform 1 0 111872 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1666464484
transform 1 0 117024 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1666464484
transform 1 0 122176 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1666464484
transform 1 0 127328 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1666464484
transform 1 0 132480 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1666464484
transform 1 0 137632 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1666464484
transform 1 0 142784 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1666464484
transform 1 0 147936 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1666464484
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1666464484
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1666464484
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1666464484
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1666464484
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1666464484
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1666464484
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1666464484
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1666464484
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1666464484
transform 1 0 62928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1666464484
transform 1 0 68080 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1666464484
transform 1 0 73232 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1666464484
transform 1 0 78384 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1666464484
transform 1 0 83536 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1666464484
transform 1 0 88688 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1666464484
transform 1 0 93840 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1666464484
transform 1 0 98992 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1666464484
transform 1 0 104144 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1666464484
transform 1 0 109296 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1666464484
transform 1 0 114448 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1666464484
transform 1 0 119600 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1666464484
transform 1 0 124752 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1666464484
transform 1 0 129904 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1666464484
transform 1 0 135056 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1666464484
transform 1 0 140208 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1666464484
transform 1 0 145360 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1666464484
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1666464484
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1666464484
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1666464484
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1666464484
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1666464484
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1666464484
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1666464484
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1666464484
transform 1 0 60352 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1666464484
transform 1 0 65504 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1666464484
transform 1 0 70656 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1666464484
transform 1 0 75808 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1666464484
transform 1 0 80960 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1666464484
transform 1 0 86112 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1666464484
transform 1 0 91264 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1666464484
transform 1 0 96416 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1666464484
transform 1 0 101568 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1666464484
transform 1 0 106720 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1666464484
transform 1 0 111872 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1666464484
transform 1 0 117024 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1666464484
transform 1 0 122176 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1666464484
transform 1 0 127328 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1666464484
transform 1 0 132480 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1666464484
transform 1 0 137632 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1666464484
transform 1 0 142784 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1666464484
transform 1 0 147936 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1666464484
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1666464484
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1666464484
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1666464484
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1666464484
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1666464484
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1666464484
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1666464484
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1666464484
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1666464484
transform 1 0 62928 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1666464484
transform 1 0 68080 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1666464484
transform 1 0 73232 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1666464484
transform 1 0 78384 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1666464484
transform 1 0 83536 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1666464484
transform 1 0 88688 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1666464484
transform 1 0 93840 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1666464484
transform 1 0 98992 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1666464484
transform 1 0 104144 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1666464484
transform 1 0 109296 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1666464484
transform 1 0 114448 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1666464484
transform 1 0 119600 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1666464484
transform 1 0 124752 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1666464484
transform 1 0 129904 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1666464484
transform 1 0 135056 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1666464484
transform 1 0 140208 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1666464484
transform 1 0 145360 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1666464484
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1666464484
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1666464484
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1666464484
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1666464484
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1666464484
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1666464484
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1666464484
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1666464484
transform 1 0 60352 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1666464484
transform 1 0 65504 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1666464484
transform 1 0 70656 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1666464484
transform 1 0 75808 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1666464484
transform 1 0 80960 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1666464484
transform 1 0 86112 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1666464484
transform 1 0 91264 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1666464484
transform 1 0 96416 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1666464484
transform 1 0 101568 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1666464484
transform 1 0 106720 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1666464484
transform 1 0 111872 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1666464484
transform 1 0 117024 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1666464484
transform 1 0 122176 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1666464484
transform 1 0 127328 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1666464484
transform 1 0 132480 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1666464484
transform 1 0 137632 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1666464484
transform 1 0 142784 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1666464484
transform 1 0 147936 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1666464484
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1666464484
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1666464484
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1666464484
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1666464484
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1666464484
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1666464484
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1666464484
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1666464484
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1666464484
transform 1 0 62928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1666464484
transform 1 0 68080 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1666464484
transform 1 0 73232 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1666464484
transform 1 0 78384 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1666464484
transform 1 0 83536 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1666464484
transform 1 0 88688 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1666464484
transform 1 0 93840 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1666464484
transform 1 0 98992 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1666464484
transform 1 0 104144 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1666464484
transform 1 0 109296 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1666464484
transform 1 0 114448 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1666464484
transform 1 0 119600 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1666464484
transform 1 0 124752 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1666464484
transform 1 0 129904 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1666464484
transform 1 0 135056 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1666464484
transform 1 0 140208 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1666464484
transform 1 0 145360 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1666464484
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1666464484
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1666464484
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1666464484
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1666464484
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1666464484
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1666464484
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1666464484
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1666464484
transform 1 0 60352 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1666464484
transform 1 0 65504 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1666464484
transform 1 0 70656 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1666464484
transform 1 0 75808 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1666464484
transform 1 0 80960 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1666464484
transform 1 0 86112 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1666464484
transform 1 0 91264 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1666464484
transform 1 0 96416 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1666464484
transform 1 0 101568 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1666464484
transform 1 0 106720 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1666464484
transform 1 0 111872 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1666464484
transform 1 0 117024 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1666464484
transform 1 0 122176 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1666464484
transform 1 0 127328 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1666464484
transform 1 0 132480 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1666464484
transform 1 0 137632 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1666464484
transform 1 0 142784 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1666464484
transform 1 0 147936 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1666464484
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1666464484
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1666464484
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1666464484
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1666464484
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1666464484
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1666464484
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1666464484
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1666464484
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1666464484
transform 1 0 62928 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1666464484
transform 1 0 68080 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1666464484
transform 1 0 73232 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1666464484
transform 1 0 78384 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1666464484
transform 1 0 83536 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1666464484
transform 1 0 88688 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1666464484
transform 1 0 93840 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1666464484
transform 1 0 98992 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1666464484
transform 1 0 104144 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1666464484
transform 1 0 109296 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1666464484
transform 1 0 114448 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1666464484
transform 1 0 119600 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1666464484
transform 1 0 124752 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1666464484
transform 1 0 129904 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1666464484
transform 1 0 135056 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1666464484
transform 1 0 140208 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1666464484
transform 1 0 145360 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1666464484
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1666464484
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1666464484
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1666464484
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1666464484
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1666464484
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1666464484
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1666464484
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1666464484
transform 1 0 60352 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1666464484
transform 1 0 65504 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1666464484
transform 1 0 70656 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1666464484
transform 1 0 75808 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1666464484
transform 1 0 80960 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1666464484
transform 1 0 86112 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1666464484
transform 1 0 91264 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1666464484
transform 1 0 96416 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1666464484
transform 1 0 101568 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1666464484
transform 1 0 106720 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1666464484
transform 1 0 111872 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1666464484
transform 1 0 117024 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1666464484
transform 1 0 122176 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1666464484
transform 1 0 127328 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1666464484
transform 1 0 132480 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1666464484
transform 1 0 137632 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1666464484
transform 1 0 142784 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1666464484
transform 1 0 147936 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1666464484
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1666464484
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1666464484
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1666464484
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1666464484
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1666464484
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1666464484
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1666464484
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1666464484
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1666464484
transform 1 0 62928 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1666464484
transform 1 0 68080 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1666464484
transform 1 0 73232 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1666464484
transform 1 0 78384 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1666464484
transform 1 0 83536 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1666464484
transform 1 0 88688 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1666464484
transform 1 0 93840 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1666464484
transform 1 0 98992 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1666464484
transform 1 0 104144 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1666464484
transform 1 0 109296 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1666464484
transform 1 0 114448 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1666464484
transform 1 0 119600 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1666464484
transform 1 0 124752 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1666464484
transform 1 0 129904 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1666464484
transform 1 0 135056 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1666464484
transform 1 0 140208 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1666464484
transform 1 0 145360 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1666464484
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1666464484
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1666464484
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1666464484
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1666464484
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1666464484
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1666464484
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1666464484
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1666464484
transform 1 0 60352 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1666464484
transform 1 0 65504 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1666464484
transform 1 0 70656 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1666464484
transform 1 0 75808 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1666464484
transform 1 0 80960 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1666464484
transform 1 0 86112 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1666464484
transform 1 0 91264 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1666464484
transform 1 0 96416 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1666464484
transform 1 0 101568 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1666464484
transform 1 0 106720 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1666464484
transform 1 0 111872 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1666464484
transform 1 0 117024 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1666464484
transform 1 0 122176 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1666464484
transform 1 0 127328 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1666464484
transform 1 0 132480 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1666464484
transform 1 0 137632 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1666464484
transform 1 0 142784 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1666464484
transform 1 0 147936 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1666464484
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1666464484
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1666464484
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1666464484
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1666464484
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1666464484
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1666464484
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1666464484
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1666464484
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1666464484
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1666464484
transform 1 0 62928 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1666464484
transform 1 0 68080 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1666464484
transform 1 0 73232 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1666464484
transform 1 0 78384 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1666464484
transform 1 0 83536 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1666464484
transform 1 0 88688 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1666464484
transform 1 0 93840 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1666464484
transform 1 0 98992 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1666464484
transform 1 0 104144 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1666464484
transform 1 0 109296 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1666464484
transform 1 0 114448 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1666464484
transform 1 0 119600 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1666464484
transform 1 0 124752 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1666464484
transform 1 0 129904 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1666464484
transform 1 0 135056 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1666464484
transform 1 0 140208 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1666464484
transform 1 0 145360 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1666464484
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1666464484
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1666464484
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1666464484
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1666464484
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1666464484
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1666464484
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1666464484
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1666464484
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1666464484
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1666464484
transform 1 0 60352 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1666464484
transform 1 0 65504 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1666464484
transform 1 0 70656 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1666464484
transform 1 0 75808 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1666464484
transform 1 0 80960 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1666464484
transform 1 0 86112 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1666464484
transform 1 0 91264 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1666464484
transform 1 0 96416 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1666464484
transform 1 0 101568 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1666464484
transform 1 0 106720 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1666464484
transform 1 0 111872 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1666464484
transform 1 0 117024 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1666464484
transform 1 0 122176 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1666464484
transform 1 0 127328 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1666464484
transform 1 0 132480 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1666464484
transform 1 0 137632 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1666464484
transform 1 0 142784 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1666464484
transform 1 0 147936 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1666464484
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1666464484
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1666464484
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1666464484
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1666464484
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1666464484
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1666464484
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1666464484
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1666464484
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1666464484
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1666464484
transform 1 0 62928 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1666464484
transform 1 0 68080 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1666464484
transform 1 0 73232 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1666464484
transform 1 0 78384 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1666464484
transform 1 0 83536 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1666464484
transform 1 0 88688 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1666464484
transform 1 0 93840 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1666464484
transform 1 0 98992 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1666464484
transform 1 0 104144 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1666464484
transform 1 0 109296 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1666464484
transform 1 0 114448 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1666464484
transform 1 0 119600 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1666464484
transform 1 0 124752 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1666464484
transform 1 0 129904 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1666464484
transform 1 0 135056 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1666464484
transform 1 0 140208 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1666464484
transform 1 0 145360 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1666464484
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1666464484
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1666464484
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1666464484
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1666464484
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1666464484
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1666464484
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1666464484
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1666464484
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1666464484
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1666464484
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1666464484
transform 1 0 60352 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1666464484
transform 1 0 65504 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1666464484
transform 1 0 70656 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1666464484
transform 1 0 75808 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1666464484
transform 1 0 80960 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1666464484
transform 1 0 86112 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1666464484
transform 1 0 91264 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1666464484
transform 1 0 96416 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1666464484
transform 1 0 101568 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1666464484
transform 1 0 106720 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1666464484
transform 1 0 111872 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1666464484
transform 1 0 117024 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1666464484
transform 1 0 122176 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1666464484
transform 1 0 127328 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1666464484
transform 1 0 132480 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1666464484
transform 1 0 137632 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1666464484
transform 1 0 142784 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1666464484
transform 1 0 147936 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1666464484
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1666464484
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1666464484
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1666464484
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1666464484
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1666464484
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1666464484
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1666464484
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1666464484
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1666464484
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1666464484
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1666464484
transform 1 0 62928 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1666464484
transform 1 0 68080 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1666464484
transform 1 0 73232 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1666464484
transform 1 0 78384 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1666464484
transform 1 0 83536 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1666464484
transform 1 0 88688 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1666464484
transform 1 0 93840 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1666464484
transform 1 0 98992 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1666464484
transform 1 0 104144 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1666464484
transform 1 0 109296 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1666464484
transform 1 0 114448 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1666464484
transform 1 0 119600 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1666464484
transform 1 0 124752 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1666464484
transform 1 0 129904 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1666464484
transform 1 0 135056 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1666464484
transform 1 0 140208 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1666464484
transform 1 0 145360 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1666464484
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1666464484
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1666464484
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1666464484
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1666464484
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1666464484
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1666464484
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1666464484
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1666464484
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1666464484
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1666464484
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1666464484
transform 1 0 60352 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1666464484
transform 1 0 65504 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1666464484
transform 1 0 70656 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1666464484
transform 1 0 75808 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1666464484
transform 1 0 80960 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1666464484
transform 1 0 86112 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1666464484
transform 1 0 91264 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1666464484
transform 1 0 96416 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1666464484
transform 1 0 101568 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1666464484
transform 1 0 106720 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1666464484
transform 1 0 111872 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1666464484
transform 1 0 117024 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1666464484
transform 1 0 122176 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1666464484
transform 1 0 127328 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1666464484
transform 1 0 132480 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1666464484
transform 1 0 137632 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1666464484
transform 1 0 142784 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1666464484
transform 1 0 147936 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1666464484
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1666464484
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1666464484
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1666464484
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1666464484
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1666464484
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1666464484
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1666464484
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1666464484
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1666464484
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1666464484
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1666464484
transform 1 0 62928 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1666464484
transform 1 0 68080 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1666464484
transform 1 0 73232 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1666464484
transform 1 0 78384 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1666464484
transform 1 0 83536 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1666464484
transform 1 0 88688 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1666464484
transform 1 0 93840 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1666464484
transform 1 0 98992 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1666464484
transform 1 0 104144 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1666464484
transform 1 0 109296 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1666464484
transform 1 0 114448 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1666464484
transform 1 0 119600 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1666464484
transform 1 0 124752 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1666464484
transform 1 0 129904 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1666464484
transform 1 0 135056 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1666464484
transform 1 0 140208 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1666464484
transform 1 0 145360 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1666464484
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1666464484
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1666464484
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1666464484
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1666464484
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1666464484
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1666464484
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1666464484
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1666464484
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1666464484
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1666464484
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1666464484
transform 1 0 60352 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1666464484
transform 1 0 65504 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1666464484
transform 1 0 70656 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1666464484
transform 1 0 75808 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1666464484
transform 1 0 80960 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1666464484
transform 1 0 86112 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1666464484
transform 1 0 91264 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1666464484
transform 1 0 96416 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1666464484
transform 1 0 101568 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1666464484
transform 1 0 106720 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1666464484
transform 1 0 111872 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1666464484
transform 1 0 117024 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1666464484
transform 1 0 122176 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1666464484
transform 1 0 127328 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1666464484
transform 1 0 132480 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1666464484
transform 1 0 137632 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1666464484
transform 1 0 142784 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1666464484
transform 1 0 147936 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1666464484
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1666464484
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1666464484
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1666464484
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1666464484
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1666464484
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1666464484
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1666464484
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1666464484
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1666464484
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1666464484
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1666464484
transform 1 0 62928 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1666464484
transform 1 0 68080 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1666464484
transform 1 0 73232 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1666464484
transform 1 0 78384 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1666464484
transform 1 0 83536 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1666464484
transform 1 0 88688 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1666464484
transform 1 0 93840 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1666464484
transform 1 0 98992 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1666464484
transform 1 0 104144 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1666464484
transform 1 0 109296 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1666464484
transform 1 0 114448 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1666464484
transform 1 0 119600 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1666464484
transform 1 0 124752 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1666464484
transform 1 0 129904 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1666464484
transform 1 0 135056 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1666464484
transform 1 0 140208 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1666464484
transform 1 0 145360 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1666464484
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1666464484
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1666464484
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1666464484
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1666464484
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1666464484
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1666464484
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1666464484
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1666464484
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1666464484
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1666464484
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1666464484
transform 1 0 60352 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1666464484
transform 1 0 65504 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1666464484
transform 1 0 70656 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1666464484
transform 1 0 75808 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1666464484
transform 1 0 80960 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1666464484
transform 1 0 86112 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1666464484
transform 1 0 91264 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1666464484
transform 1 0 96416 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1666464484
transform 1 0 101568 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1666464484
transform 1 0 106720 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1666464484
transform 1 0 111872 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1666464484
transform 1 0 117024 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1666464484
transform 1 0 122176 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1666464484
transform 1 0 127328 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1666464484
transform 1 0 132480 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1666464484
transform 1 0 137632 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1666464484
transform 1 0 142784 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1666464484
transform 1 0 147936 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1666464484
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1666464484
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1666464484
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1666464484
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1666464484
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1666464484
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1666464484
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1666464484
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1666464484
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1666464484
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1666464484
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1666464484
transform 1 0 62928 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1666464484
transform 1 0 68080 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1666464484
transform 1 0 73232 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1666464484
transform 1 0 78384 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1666464484
transform 1 0 83536 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1666464484
transform 1 0 88688 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1666464484
transform 1 0 93840 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1666464484
transform 1 0 98992 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1666464484
transform 1 0 104144 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1666464484
transform 1 0 109296 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1666464484
transform 1 0 114448 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1666464484
transform 1 0 119600 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1666464484
transform 1 0 124752 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1666464484
transform 1 0 129904 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1666464484
transform 1 0 135056 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1666464484
transform 1 0 140208 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1666464484
transform 1 0 145360 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1666464484
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1666464484
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1666464484
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1666464484
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1666464484
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1666464484
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1666464484
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1666464484
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1666464484
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1666464484
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1666464484
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1666464484
transform 1 0 60352 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1666464484
transform 1 0 65504 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1666464484
transform 1 0 70656 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1666464484
transform 1 0 75808 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1666464484
transform 1 0 80960 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1666464484
transform 1 0 86112 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1666464484
transform 1 0 91264 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1666464484
transform 1 0 96416 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1666464484
transform 1 0 101568 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1666464484
transform 1 0 106720 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1666464484
transform 1 0 111872 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1666464484
transform 1 0 117024 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1666464484
transform 1 0 122176 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1666464484
transform 1 0 127328 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1666464484
transform 1 0 132480 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1666464484
transform 1 0 137632 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1666464484
transform 1 0 142784 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1666464484
transform 1 0 147936 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1666464484
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1666464484
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1666464484
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1666464484
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1666464484
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1666464484
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1666464484
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1666464484
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1666464484
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1666464484
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1666464484
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1666464484
transform 1 0 62928 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1666464484
transform 1 0 68080 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1666464484
transform 1 0 73232 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1666464484
transform 1 0 78384 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1666464484
transform 1 0 83536 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1666464484
transform 1 0 88688 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1666464484
transform 1 0 93840 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1666464484
transform 1 0 98992 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1666464484
transform 1 0 104144 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1666464484
transform 1 0 109296 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1666464484
transform 1 0 114448 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1666464484
transform 1 0 119600 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1666464484
transform 1 0 124752 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1666464484
transform 1 0 129904 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1666464484
transform 1 0 135056 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1666464484
transform 1 0 140208 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1666464484
transform 1 0 145360 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1666464484
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1666464484
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1666464484
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1666464484
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1666464484
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1666464484
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1666464484
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1666464484
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1666464484
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1666464484
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1666464484
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1666464484
transform 1 0 60352 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1666464484
transform 1 0 65504 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1666464484
transform 1 0 70656 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1666464484
transform 1 0 75808 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1666464484
transform 1 0 80960 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1666464484
transform 1 0 86112 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1666464484
transform 1 0 91264 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1666464484
transform 1 0 96416 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1666464484
transform 1 0 101568 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1666464484
transform 1 0 106720 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1666464484
transform 1 0 111872 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1666464484
transform 1 0 117024 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1666464484
transform 1 0 122176 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1666464484
transform 1 0 127328 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1666464484
transform 1 0 132480 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1666464484
transform 1 0 137632 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1666464484
transform 1 0 142784 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1666464484
transform 1 0 147936 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1666464484
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1666464484
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1666464484
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1666464484
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1666464484
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1666464484
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1666464484
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1666464484
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1666464484
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1666464484
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1666464484
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1666464484
transform 1 0 62928 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1666464484
transform 1 0 68080 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1666464484
transform 1 0 73232 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1666464484
transform 1 0 78384 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1666464484
transform 1 0 83536 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1666464484
transform 1 0 88688 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1666464484
transform 1 0 93840 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1666464484
transform 1 0 98992 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1666464484
transform 1 0 104144 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1666464484
transform 1 0 109296 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1666464484
transform 1 0 114448 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1666464484
transform 1 0 119600 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1666464484
transform 1 0 124752 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1666464484
transform 1 0 129904 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1666464484
transform 1 0 135056 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1666464484
transform 1 0 140208 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1666464484
transform 1 0 145360 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1666464484
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1666464484
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1666464484
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1666464484
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1666464484
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1666464484
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1666464484
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1666464484
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1666464484
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1666464484
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1666464484
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1666464484
transform 1 0 60352 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1666464484
transform 1 0 65504 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1666464484
transform 1 0 70656 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1666464484
transform 1 0 75808 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1666464484
transform 1 0 80960 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1666464484
transform 1 0 86112 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1666464484
transform 1 0 91264 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1666464484
transform 1 0 96416 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1666464484
transform 1 0 101568 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1666464484
transform 1 0 106720 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1666464484
transform 1 0 111872 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1666464484
transform 1 0 117024 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1666464484
transform 1 0 122176 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1666464484
transform 1 0 127328 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1666464484
transform 1 0 132480 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1666464484
transform 1 0 137632 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1666464484
transform 1 0 142784 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1666464484
transform 1 0 147936 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1666464484
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1666464484
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1666464484
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1666464484
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1666464484
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1666464484
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1666464484
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1666464484
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1666464484
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1666464484
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1666464484
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1666464484
transform 1 0 62928 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1666464484
transform 1 0 68080 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1666464484
transform 1 0 73232 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1666464484
transform 1 0 78384 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1666464484
transform 1 0 83536 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1666464484
transform 1 0 88688 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1666464484
transform 1 0 93840 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1666464484
transform 1 0 98992 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1666464484
transform 1 0 104144 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1666464484
transform 1 0 109296 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1666464484
transform 1 0 114448 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1666464484
transform 1 0 119600 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1666464484
transform 1 0 124752 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1666464484
transform 1 0 129904 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1666464484
transform 1 0 135056 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1666464484
transform 1 0 140208 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1666464484
transform 1 0 145360 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1666464484
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1666464484
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1666464484
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1666464484
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1666464484
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1666464484
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1666464484
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1666464484
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1666464484
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1666464484
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1666464484
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1666464484
transform 1 0 60352 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1666464484
transform 1 0 65504 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1666464484
transform 1 0 70656 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1666464484
transform 1 0 75808 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1666464484
transform 1 0 80960 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1666464484
transform 1 0 86112 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1666464484
transform 1 0 91264 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1666464484
transform 1 0 96416 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1666464484
transform 1 0 101568 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1666464484
transform 1 0 106720 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1666464484
transform 1 0 111872 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1666464484
transform 1 0 117024 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1666464484
transform 1 0 122176 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1666464484
transform 1 0 127328 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1666464484
transform 1 0 132480 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1666464484
transform 1 0 137632 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1666464484
transform 1 0 142784 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1666464484
transform 1 0 147936 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1666464484
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1666464484
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1666464484
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1666464484
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1666464484
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1666464484
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1666464484
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1666464484
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1666464484
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1666464484
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1666464484
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1666464484
transform 1 0 62928 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1666464484
transform 1 0 68080 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1666464484
transform 1 0 73232 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1666464484
transform 1 0 78384 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1399
timestamp 1666464484
transform 1 0 83536 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1400
timestamp 1666464484
transform 1 0 88688 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1401
timestamp 1666464484
transform 1 0 93840 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1402
timestamp 1666464484
transform 1 0 98992 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1403
timestamp 1666464484
transform 1 0 104144 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1404
timestamp 1666464484
transform 1 0 109296 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1405
timestamp 1666464484
transform 1 0 114448 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1406
timestamp 1666464484
transform 1 0 119600 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1407
timestamp 1666464484
transform 1 0 124752 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1408
timestamp 1666464484
transform 1 0 129904 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1409
timestamp 1666464484
transform 1 0 135056 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1410
timestamp 1666464484
transform 1 0 140208 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1411
timestamp 1666464484
transform 1 0 145360 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1412
timestamp 1666464484
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1413
timestamp 1666464484
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1414
timestamp 1666464484
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1415
timestamp 1666464484
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1416
timestamp 1666464484
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1417
timestamp 1666464484
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1418
timestamp 1666464484
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1419
timestamp 1666464484
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1420
timestamp 1666464484
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1421
timestamp 1666464484
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1422
timestamp 1666464484
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1423
timestamp 1666464484
transform 1 0 60352 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1424
timestamp 1666464484
transform 1 0 65504 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1425
timestamp 1666464484
transform 1 0 70656 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1426
timestamp 1666464484
transform 1 0 75808 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1427
timestamp 1666464484
transform 1 0 80960 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1428
timestamp 1666464484
transform 1 0 86112 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1429
timestamp 1666464484
transform 1 0 91264 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1430
timestamp 1666464484
transform 1 0 96416 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1431
timestamp 1666464484
transform 1 0 101568 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1432
timestamp 1666464484
transform 1 0 106720 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1433
timestamp 1666464484
transform 1 0 111872 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1434
timestamp 1666464484
transform 1 0 117024 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1435
timestamp 1666464484
transform 1 0 122176 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1436
timestamp 1666464484
transform 1 0 127328 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1437
timestamp 1666464484
transform 1 0 132480 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1438
timestamp 1666464484
transform 1 0 137632 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1439
timestamp 1666464484
transform 1 0 142784 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1440
timestamp 1666464484
transform 1 0 147936 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1441
timestamp 1666464484
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1442
timestamp 1666464484
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1443
timestamp 1666464484
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1444
timestamp 1666464484
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1445
timestamp 1666464484
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1446
timestamp 1666464484
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1447
timestamp 1666464484
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1448
timestamp 1666464484
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1449
timestamp 1666464484
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1450
timestamp 1666464484
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1451
timestamp 1666464484
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1452
timestamp 1666464484
transform 1 0 62928 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1453
timestamp 1666464484
transform 1 0 68080 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1454
timestamp 1666464484
transform 1 0 73232 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1455
timestamp 1666464484
transform 1 0 78384 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1456
timestamp 1666464484
transform 1 0 83536 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1457
timestamp 1666464484
transform 1 0 88688 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1458
timestamp 1666464484
transform 1 0 93840 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1459
timestamp 1666464484
transform 1 0 98992 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1460
timestamp 1666464484
transform 1 0 104144 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1461
timestamp 1666464484
transform 1 0 109296 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1462
timestamp 1666464484
transform 1 0 114448 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1463
timestamp 1666464484
transform 1 0 119600 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1464
timestamp 1666464484
transform 1 0 124752 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1465
timestamp 1666464484
transform 1 0 129904 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1466
timestamp 1666464484
transform 1 0 135056 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1467
timestamp 1666464484
transform 1 0 140208 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1468
timestamp 1666464484
transform 1 0 145360 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1469
timestamp 1666464484
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1470
timestamp 1666464484
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1471
timestamp 1666464484
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1472
timestamp 1666464484
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1473
timestamp 1666464484
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1474
timestamp 1666464484
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1475
timestamp 1666464484
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1476
timestamp 1666464484
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1477
timestamp 1666464484
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1478
timestamp 1666464484
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1479
timestamp 1666464484
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1480
timestamp 1666464484
transform 1 0 60352 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1481
timestamp 1666464484
transform 1 0 65504 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1482
timestamp 1666464484
transform 1 0 70656 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1483
timestamp 1666464484
transform 1 0 75808 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1484
timestamp 1666464484
transform 1 0 80960 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1485
timestamp 1666464484
transform 1 0 86112 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1486
timestamp 1666464484
transform 1 0 91264 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1487
timestamp 1666464484
transform 1 0 96416 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1488
timestamp 1666464484
transform 1 0 101568 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1489
timestamp 1666464484
transform 1 0 106720 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1490
timestamp 1666464484
transform 1 0 111872 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1491
timestamp 1666464484
transform 1 0 117024 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1492
timestamp 1666464484
transform 1 0 122176 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1493
timestamp 1666464484
transform 1 0 127328 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1494
timestamp 1666464484
transform 1 0 132480 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1495
timestamp 1666464484
transform 1 0 137632 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1496
timestamp 1666464484
transform 1 0 142784 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1497
timestamp 1666464484
transform 1 0 147936 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1498
timestamp 1666464484
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1499
timestamp 1666464484
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1500
timestamp 1666464484
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1501
timestamp 1666464484
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1502
timestamp 1666464484
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1503
timestamp 1666464484
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1504
timestamp 1666464484
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1505
timestamp 1666464484
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1506
timestamp 1666464484
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1507
timestamp 1666464484
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1508
timestamp 1666464484
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1509
timestamp 1666464484
transform 1 0 62928 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1510
timestamp 1666464484
transform 1 0 68080 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1511
timestamp 1666464484
transform 1 0 73232 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1512
timestamp 1666464484
transform 1 0 78384 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1513
timestamp 1666464484
transform 1 0 83536 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1514
timestamp 1666464484
transform 1 0 88688 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1515
timestamp 1666464484
transform 1 0 93840 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1516
timestamp 1666464484
transform 1 0 98992 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1517
timestamp 1666464484
transform 1 0 104144 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1518
timestamp 1666464484
transform 1 0 109296 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1519
timestamp 1666464484
transform 1 0 114448 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1520
timestamp 1666464484
transform 1 0 119600 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1521
timestamp 1666464484
transform 1 0 124752 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1522
timestamp 1666464484
transform 1 0 129904 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1523
timestamp 1666464484
transform 1 0 135056 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1524
timestamp 1666464484
transform 1 0 140208 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1525
timestamp 1666464484
transform 1 0 145360 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1526
timestamp 1666464484
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1527
timestamp 1666464484
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1528
timestamp 1666464484
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1529
timestamp 1666464484
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1530
timestamp 1666464484
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1531
timestamp 1666464484
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1532
timestamp 1666464484
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1533
timestamp 1666464484
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1534
timestamp 1666464484
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1535
timestamp 1666464484
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1536
timestamp 1666464484
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1537
timestamp 1666464484
transform 1 0 60352 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1538
timestamp 1666464484
transform 1 0 65504 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1539
timestamp 1666464484
transform 1 0 70656 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1540
timestamp 1666464484
transform 1 0 75808 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1541
timestamp 1666464484
transform 1 0 80960 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1542
timestamp 1666464484
transform 1 0 86112 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1543
timestamp 1666464484
transform 1 0 91264 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1544
timestamp 1666464484
transform 1 0 96416 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1545
timestamp 1666464484
transform 1 0 101568 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1546
timestamp 1666464484
transform 1 0 106720 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1547
timestamp 1666464484
transform 1 0 111872 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1548
timestamp 1666464484
transform 1 0 117024 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1549
timestamp 1666464484
transform 1 0 122176 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1550
timestamp 1666464484
transform 1 0 127328 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1551
timestamp 1666464484
transform 1 0 132480 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1552
timestamp 1666464484
transform 1 0 137632 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1553
timestamp 1666464484
transform 1 0 142784 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1554
timestamp 1666464484
transform 1 0 147936 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1555
timestamp 1666464484
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1556
timestamp 1666464484
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1557
timestamp 1666464484
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1558
timestamp 1666464484
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1559
timestamp 1666464484
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1560
timestamp 1666464484
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1561
timestamp 1666464484
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1562
timestamp 1666464484
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1563
timestamp 1666464484
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1564
timestamp 1666464484
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1565
timestamp 1666464484
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1566
timestamp 1666464484
transform 1 0 62928 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1567
timestamp 1666464484
transform 1 0 68080 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1568
timestamp 1666464484
transform 1 0 73232 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1569
timestamp 1666464484
transform 1 0 78384 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1570
timestamp 1666464484
transform 1 0 83536 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1571
timestamp 1666464484
transform 1 0 88688 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1572
timestamp 1666464484
transform 1 0 93840 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1573
timestamp 1666464484
transform 1 0 98992 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1574
timestamp 1666464484
transform 1 0 104144 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1575
timestamp 1666464484
transform 1 0 109296 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1576
timestamp 1666464484
transform 1 0 114448 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1577
timestamp 1666464484
transform 1 0 119600 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1578
timestamp 1666464484
transform 1 0 124752 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1579
timestamp 1666464484
transform 1 0 129904 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1580
timestamp 1666464484
transform 1 0 135056 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1581
timestamp 1666464484
transform 1 0 140208 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1582
timestamp 1666464484
transform 1 0 145360 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1583
timestamp 1666464484
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1584
timestamp 1666464484
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1585
timestamp 1666464484
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1586
timestamp 1666464484
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1587
timestamp 1666464484
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1588
timestamp 1666464484
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1589
timestamp 1666464484
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1590
timestamp 1666464484
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1591
timestamp 1666464484
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1592
timestamp 1666464484
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1593
timestamp 1666464484
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1594
timestamp 1666464484
transform 1 0 60352 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1595
timestamp 1666464484
transform 1 0 65504 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1596
timestamp 1666464484
transform 1 0 70656 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1597
timestamp 1666464484
transform 1 0 75808 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1598
timestamp 1666464484
transform 1 0 80960 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1599
timestamp 1666464484
transform 1 0 86112 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1600
timestamp 1666464484
transform 1 0 91264 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1601
timestamp 1666464484
transform 1 0 96416 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1602
timestamp 1666464484
transform 1 0 101568 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1603
timestamp 1666464484
transform 1 0 106720 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1604
timestamp 1666464484
transform 1 0 111872 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1605
timestamp 1666464484
transform 1 0 117024 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1606
timestamp 1666464484
transform 1 0 122176 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1607
timestamp 1666464484
transform 1 0 127328 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1608
timestamp 1666464484
transform 1 0 132480 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1609
timestamp 1666464484
transform 1 0 137632 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1610
timestamp 1666464484
transform 1 0 142784 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1611
timestamp 1666464484
transform 1 0 147936 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1612
timestamp 1666464484
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1613
timestamp 1666464484
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1614
timestamp 1666464484
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1615
timestamp 1666464484
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1616
timestamp 1666464484
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1617
timestamp 1666464484
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1618
timestamp 1666464484
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1619
timestamp 1666464484
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1620
timestamp 1666464484
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1621
timestamp 1666464484
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1622
timestamp 1666464484
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1623
timestamp 1666464484
transform 1 0 62928 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1624
timestamp 1666464484
transform 1 0 68080 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1625
timestamp 1666464484
transform 1 0 73232 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1626
timestamp 1666464484
transform 1 0 78384 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1627
timestamp 1666464484
transform 1 0 83536 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1628
timestamp 1666464484
transform 1 0 88688 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1629
timestamp 1666464484
transform 1 0 93840 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1630
timestamp 1666464484
transform 1 0 98992 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1631
timestamp 1666464484
transform 1 0 104144 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1632
timestamp 1666464484
transform 1 0 109296 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1633
timestamp 1666464484
transform 1 0 114448 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1634
timestamp 1666464484
transform 1 0 119600 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1635
timestamp 1666464484
transform 1 0 124752 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1636
timestamp 1666464484
transform 1 0 129904 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1637
timestamp 1666464484
transform 1 0 135056 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1638
timestamp 1666464484
transform 1 0 140208 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1639
timestamp 1666464484
transform 1 0 145360 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1640
timestamp 1666464484
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1641
timestamp 1666464484
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1642
timestamp 1666464484
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1643
timestamp 1666464484
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1644
timestamp 1666464484
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1645
timestamp 1666464484
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1646
timestamp 1666464484
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1647
timestamp 1666464484
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1648
timestamp 1666464484
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1649
timestamp 1666464484
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1650
timestamp 1666464484
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1651
timestamp 1666464484
transform 1 0 60352 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1652
timestamp 1666464484
transform 1 0 65504 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1653
timestamp 1666464484
transform 1 0 70656 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1654
timestamp 1666464484
transform 1 0 75808 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1655
timestamp 1666464484
transform 1 0 80960 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1656
timestamp 1666464484
transform 1 0 86112 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1657
timestamp 1666464484
transform 1 0 91264 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1658
timestamp 1666464484
transform 1 0 96416 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1659
timestamp 1666464484
transform 1 0 101568 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1660
timestamp 1666464484
transform 1 0 106720 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1661
timestamp 1666464484
transform 1 0 111872 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1662
timestamp 1666464484
transform 1 0 117024 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1663
timestamp 1666464484
transform 1 0 122176 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1664
timestamp 1666464484
transform 1 0 127328 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1665
timestamp 1666464484
transform 1 0 132480 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1666
timestamp 1666464484
transform 1 0 137632 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1667
timestamp 1666464484
transform 1 0 142784 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1668
timestamp 1666464484
transform 1 0 147936 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1669
timestamp 1666464484
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1670
timestamp 1666464484
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1671
timestamp 1666464484
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1672
timestamp 1666464484
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1673
timestamp 1666464484
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1674
timestamp 1666464484
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1675
timestamp 1666464484
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1676
timestamp 1666464484
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1677
timestamp 1666464484
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1678
timestamp 1666464484
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1679
timestamp 1666464484
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1680
timestamp 1666464484
transform 1 0 62928 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1681
timestamp 1666464484
transform 1 0 68080 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1682
timestamp 1666464484
transform 1 0 73232 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1683
timestamp 1666464484
transform 1 0 78384 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1684
timestamp 1666464484
transform 1 0 83536 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1685
timestamp 1666464484
transform 1 0 88688 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1686
timestamp 1666464484
transform 1 0 93840 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1687
timestamp 1666464484
transform 1 0 98992 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1688
timestamp 1666464484
transform 1 0 104144 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1689
timestamp 1666464484
transform 1 0 109296 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1690
timestamp 1666464484
transform 1 0 114448 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1691
timestamp 1666464484
transform 1 0 119600 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1692
timestamp 1666464484
transform 1 0 124752 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1693
timestamp 1666464484
transform 1 0 129904 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1694
timestamp 1666464484
transform 1 0 135056 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1695
timestamp 1666464484
transform 1 0 140208 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1696
timestamp 1666464484
transform 1 0 145360 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1697
timestamp 1666464484
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1698
timestamp 1666464484
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1699
timestamp 1666464484
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1700
timestamp 1666464484
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1701
timestamp 1666464484
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1702
timestamp 1666464484
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1703
timestamp 1666464484
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1704
timestamp 1666464484
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1705
timestamp 1666464484
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1706
timestamp 1666464484
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1707
timestamp 1666464484
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1708
timestamp 1666464484
transform 1 0 60352 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1709
timestamp 1666464484
transform 1 0 65504 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1710
timestamp 1666464484
transform 1 0 70656 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1711
timestamp 1666464484
transform 1 0 75808 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1712
timestamp 1666464484
transform 1 0 80960 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1713
timestamp 1666464484
transform 1 0 86112 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1714
timestamp 1666464484
transform 1 0 91264 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1715
timestamp 1666464484
transform 1 0 96416 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1716
timestamp 1666464484
transform 1 0 101568 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1717
timestamp 1666464484
transform 1 0 106720 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1718
timestamp 1666464484
transform 1 0 111872 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1719
timestamp 1666464484
transform 1 0 117024 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1720
timestamp 1666464484
transform 1 0 122176 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1721
timestamp 1666464484
transform 1 0 127328 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1722
timestamp 1666464484
transform 1 0 132480 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1723
timestamp 1666464484
transform 1 0 137632 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1724
timestamp 1666464484
transform 1 0 142784 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1725
timestamp 1666464484
transform 1 0 147936 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1726
timestamp 1666464484
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1727
timestamp 1666464484
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1728
timestamp 1666464484
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1729
timestamp 1666464484
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1730
timestamp 1666464484
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1731
timestamp 1666464484
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1732
timestamp 1666464484
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1733
timestamp 1666464484
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1734
timestamp 1666464484
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1735
timestamp 1666464484
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1736
timestamp 1666464484
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1737
timestamp 1666464484
transform 1 0 62928 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1738
timestamp 1666464484
transform 1 0 68080 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1739
timestamp 1666464484
transform 1 0 73232 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1740
timestamp 1666464484
transform 1 0 78384 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1741
timestamp 1666464484
transform 1 0 83536 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1742
timestamp 1666464484
transform 1 0 88688 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1743
timestamp 1666464484
transform 1 0 93840 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1744
timestamp 1666464484
transform 1 0 98992 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1745
timestamp 1666464484
transform 1 0 104144 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1746
timestamp 1666464484
transform 1 0 109296 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1747
timestamp 1666464484
transform 1 0 114448 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1748
timestamp 1666464484
transform 1 0 119600 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1749
timestamp 1666464484
transform 1 0 124752 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1750
timestamp 1666464484
transform 1 0 129904 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1751
timestamp 1666464484
transform 1 0 135056 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1752
timestamp 1666464484
transform 1 0 140208 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1753
timestamp 1666464484
transform 1 0 145360 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1754
timestamp 1666464484
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1755
timestamp 1666464484
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1756
timestamp 1666464484
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1757
timestamp 1666464484
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1758
timestamp 1666464484
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1759
timestamp 1666464484
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1760
timestamp 1666464484
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1761
timestamp 1666464484
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1762
timestamp 1666464484
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1763
timestamp 1666464484
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1764
timestamp 1666464484
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1765
timestamp 1666464484
transform 1 0 60352 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1766
timestamp 1666464484
transform 1 0 65504 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1767
timestamp 1666464484
transform 1 0 70656 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1768
timestamp 1666464484
transform 1 0 75808 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1769
timestamp 1666464484
transform 1 0 80960 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1770
timestamp 1666464484
transform 1 0 86112 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1771
timestamp 1666464484
transform 1 0 91264 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1772
timestamp 1666464484
transform 1 0 96416 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1773
timestamp 1666464484
transform 1 0 101568 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1774
timestamp 1666464484
transform 1 0 106720 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1775
timestamp 1666464484
transform 1 0 111872 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1776
timestamp 1666464484
transform 1 0 117024 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1777
timestamp 1666464484
transform 1 0 122176 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1778
timestamp 1666464484
transform 1 0 127328 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1779
timestamp 1666464484
transform 1 0 132480 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1780
timestamp 1666464484
transform 1 0 137632 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1781
timestamp 1666464484
transform 1 0 142784 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1782
timestamp 1666464484
transform 1 0 147936 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1783
timestamp 1666464484
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1784
timestamp 1666464484
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1785
timestamp 1666464484
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1786
timestamp 1666464484
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1787
timestamp 1666464484
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1788
timestamp 1666464484
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1789
timestamp 1666464484
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1790
timestamp 1666464484
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1791
timestamp 1666464484
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1792
timestamp 1666464484
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1793
timestamp 1666464484
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1794
timestamp 1666464484
transform 1 0 62928 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1795
timestamp 1666464484
transform 1 0 68080 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1796
timestamp 1666464484
transform 1 0 73232 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1797
timestamp 1666464484
transform 1 0 78384 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1798
timestamp 1666464484
transform 1 0 83536 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1799
timestamp 1666464484
transform 1 0 88688 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1800
timestamp 1666464484
transform 1 0 93840 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1801
timestamp 1666464484
transform 1 0 98992 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1802
timestamp 1666464484
transform 1 0 104144 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1803
timestamp 1666464484
transform 1 0 109296 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1804
timestamp 1666464484
transform 1 0 114448 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1805
timestamp 1666464484
transform 1 0 119600 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1806
timestamp 1666464484
transform 1 0 124752 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1807
timestamp 1666464484
transform 1 0 129904 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1808
timestamp 1666464484
transform 1 0 135056 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1809
timestamp 1666464484
transform 1 0 140208 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1810
timestamp 1666464484
transform 1 0 145360 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1811
timestamp 1666464484
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1812
timestamp 1666464484
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1813
timestamp 1666464484
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1814
timestamp 1666464484
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1815
timestamp 1666464484
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1816
timestamp 1666464484
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1817
timestamp 1666464484
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1818
timestamp 1666464484
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1819
timestamp 1666464484
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1820
timestamp 1666464484
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1821
timestamp 1666464484
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1822
timestamp 1666464484
transform 1 0 60352 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1823
timestamp 1666464484
transform 1 0 65504 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1824
timestamp 1666464484
transform 1 0 70656 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1825
timestamp 1666464484
transform 1 0 75808 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1826
timestamp 1666464484
transform 1 0 80960 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1827
timestamp 1666464484
transform 1 0 86112 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1828
timestamp 1666464484
transform 1 0 91264 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1829
timestamp 1666464484
transform 1 0 96416 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1830
timestamp 1666464484
transform 1 0 101568 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1831
timestamp 1666464484
transform 1 0 106720 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1832
timestamp 1666464484
transform 1 0 111872 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1833
timestamp 1666464484
transform 1 0 117024 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1834
timestamp 1666464484
transform 1 0 122176 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1835
timestamp 1666464484
transform 1 0 127328 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1836
timestamp 1666464484
transform 1 0 132480 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1837
timestamp 1666464484
transform 1 0 137632 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1838
timestamp 1666464484
transform 1 0 142784 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1839
timestamp 1666464484
transform 1 0 147936 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1840
timestamp 1666464484
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1841
timestamp 1666464484
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1842
timestamp 1666464484
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1843
timestamp 1666464484
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1844
timestamp 1666464484
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1845
timestamp 1666464484
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1846
timestamp 1666464484
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1847
timestamp 1666464484
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1848
timestamp 1666464484
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1849
timestamp 1666464484
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1850
timestamp 1666464484
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1851
timestamp 1666464484
transform 1 0 62928 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1852
timestamp 1666464484
transform 1 0 68080 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1853
timestamp 1666464484
transform 1 0 73232 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1854
timestamp 1666464484
transform 1 0 78384 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1855
timestamp 1666464484
transform 1 0 83536 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1856
timestamp 1666464484
transform 1 0 88688 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1857
timestamp 1666464484
transform 1 0 93840 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1858
timestamp 1666464484
transform 1 0 98992 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1859
timestamp 1666464484
transform 1 0 104144 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1860
timestamp 1666464484
transform 1 0 109296 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1861
timestamp 1666464484
transform 1 0 114448 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1862
timestamp 1666464484
transform 1 0 119600 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1863
timestamp 1666464484
transform 1 0 124752 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1864
timestamp 1666464484
transform 1 0 129904 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1865
timestamp 1666464484
transform 1 0 135056 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1866
timestamp 1666464484
transform 1 0 140208 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1867
timestamp 1666464484
transform 1 0 145360 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1868
timestamp 1666464484
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1869
timestamp 1666464484
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1870
timestamp 1666464484
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1871
timestamp 1666464484
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1872
timestamp 1666464484
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1873
timestamp 1666464484
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1874
timestamp 1666464484
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1875
timestamp 1666464484
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1876
timestamp 1666464484
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1877
timestamp 1666464484
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1878
timestamp 1666464484
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1879
timestamp 1666464484
transform 1 0 60352 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1880
timestamp 1666464484
transform 1 0 65504 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1881
timestamp 1666464484
transform 1 0 70656 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1882
timestamp 1666464484
transform 1 0 75808 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1883
timestamp 1666464484
transform 1 0 80960 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1884
timestamp 1666464484
transform 1 0 86112 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1885
timestamp 1666464484
transform 1 0 91264 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1886
timestamp 1666464484
transform 1 0 96416 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1887
timestamp 1666464484
transform 1 0 101568 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1888
timestamp 1666464484
transform 1 0 106720 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1889
timestamp 1666464484
transform 1 0 111872 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1890
timestamp 1666464484
transform 1 0 117024 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1891
timestamp 1666464484
transform 1 0 122176 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1892
timestamp 1666464484
transform 1 0 127328 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1893
timestamp 1666464484
transform 1 0 132480 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1894
timestamp 1666464484
transform 1 0 137632 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1895
timestamp 1666464484
transform 1 0 142784 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1896
timestamp 1666464484
transform 1 0 147936 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1897
timestamp 1666464484
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1898
timestamp 1666464484
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1899
timestamp 1666464484
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1900
timestamp 1666464484
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1901
timestamp 1666464484
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1902
timestamp 1666464484
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1903
timestamp 1666464484
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1904
timestamp 1666464484
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1905
timestamp 1666464484
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1906
timestamp 1666464484
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1907
timestamp 1666464484
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1908
timestamp 1666464484
transform 1 0 62928 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1909
timestamp 1666464484
transform 1 0 68080 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1910
timestamp 1666464484
transform 1 0 73232 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1911
timestamp 1666464484
transform 1 0 78384 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1912
timestamp 1666464484
transform 1 0 83536 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1913
timestamp 1666464484
transform 1 0 88688 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1914
timestamp 1666464484
transform 1 0 93840 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1915
timestamp 1666464484
transform 1 0 98992 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1916
timestamp 1666464484
transform 1 0 104144 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1917
timestamp 1666464484
transform 1 0 109296 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1918
timestamp 1666464484
transform 1 0 114448 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1919
timestamp 1666464484
transform 1 0 119600 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1920
timestamp 1666464484
transform 1 0 124752 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1921
timestamp 1666464484
transform 1 0 129904 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1922
timestamp 1666464484
transform 1 0 135056 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1923
timestamp 1666464484
transform 1 0 140208 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1924
timestamp 1666464484
transform 1 0 145360 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1925
timestamp 1666464484
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1926
timestamp 1666464484
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1927
timestamp 1666464484
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1928
timestamp 1666464484
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1929
timestamp 1666464484
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1930
timestamp 1666464484
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1931
timestamp 1666464484
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1932
timestamp 1666464484
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1933
timestamp 1666464484
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1934
timestamp 1666464484
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1935
timestamp 1666464484
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1936
timestamp 1666464484
transform 1 0 60352 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1937
timestamp 1666464484
transform 1 0 65504 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1938
timestamp 1666464484
transform 1 0 70656 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1939
timestamp 1666464484
transform 1 0 75808 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1940
timestamp 1666464484
transform 1 0 80960 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1941
timestamp 1666464484
transform 1 0 86112 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1942
timestamp 1666464484
transform 1 0 91264 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1943
timestamp 1666464484
transform 1 0 96416 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1944
timestamp 1666464484
transform 1 0 101568 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1945
timestamp 1666464484
transform 1 0 106720 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1946
timestamp 1666464484
transform 1 0 111872 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1947
timestamp 1666464484
transform 1 0 117024 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1948
timestamp 1666464484
transform 1 0 122176 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1949
timestamp 1666464484
transform 1 0 127328 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1950
timestamp 1666464484
transform 1 0 132480 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1951
timestamp 1666464484
transform 1 0 137632 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1952
timestamp 1666464484
transform 1 0 142784 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1953
timestamp 1666464484
transform 1 0 147936 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1954
timestamp 1666464484
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1955
timestamp 1666464484
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1956
timestamp 1666464484
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1957
timestamp 1666464484
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1958
timestamp 1666464484
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1959
timestamp 1666464484
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1960
timestamp 1666464484
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1961
timestamp 1666464484
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1962
timestamp 1666464484
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1963
timestamp 1666464484
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1964
timestamp 1666464484
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1965
timestamp 1666464484
transform 1 0 62928 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1966
timestamp 1666464484
transform 1 0 68080 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1967
timestamp 1666464484
transform 1 0 73232 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1968
timestamp 1666464484
transform 1 0 78384 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1969
timestamp 1666464484
transform 1 0 83536 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1970
timestamp 1666464484
transform 1 0 88688 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1971
timestamp 1666464484
transform 1 0 93840 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1972
timestamp 1666464484
transform 1 0 98992 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1973
timestamp 1666464484
transform 1 0 104144 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1974
timestamp 1666464484
transform 1 0 109296 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1975
timestamp 1666464484
transform 1 0 114448 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1976
timestamp 1666464484
transform 1 0 119600 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1977
timestamp 1666464484
transform 1 0 124752 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1978
timestamp 1666464484
transform 1 0 129904 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1979
timestamp 1666464484
transform 1 0 135056 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1980
timestamp 1666464484
transform 1 0 140208 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1981
timestamp 1666464484
transform 1 0 145360 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1982
timestamp 1666464484
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1983
timestamp 1666464484
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1984
timestamp 1666464484
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1985
timestamp 1666464484
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1986
timestamp 1666464484
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1987
timestamp 1666464484
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1988
timestamp 1666464484
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1989
timestamp 1666464484
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1990
timestamp 1666464484
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1991
timestamp 1666464484
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1992
timestamp 1666464484
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1993
timestamp 1666464484
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1994
timestamp 1666464484
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1995
timestamp 1666464484
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1996
timestamp 1666464484
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1997
timestamp 1666464484
transform 1 0 42320 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1998
timestamp 1666464484
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1999
timestamp 1666464484
transform 1 0 47472 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2000
timestamp 1666464484
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2001
timestamp 1666464484
transform 1 0 52624 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2002
timestamp 1666464484
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2003
timestamp 1666464484
transform 1 0 57776 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2004
timestamp 1666464484
transform 1 0 60352 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2005
timestamp 1666464484
transform 1 0 62928 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2006
timestamp 1666464484
transform 1 0 65504 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2007
timestamp 1666464484
transform 1 0 68080 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2008
timestamp 1666464484
transform 1 0 70656 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2009
timestamp 1666464484
transform 1 0 73232 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2010
timestamp 1666464484
transform 1 0 75808 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2011
timestamp 1666464484
transform 1 0 78384 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2012
timestamp 1666464484
transform 1 0 80960 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2013
timestamp 1666464484
transform 1 0 83536 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2014
timestamp 1666464484
transform 1 0 86112 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2015
timestamp 1666464484
transform 1 0 88688 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2016
timestamp 1666464484
transform 1 0 91264 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2017
timestamp 1666464484
transform 1 0 93840 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2018
timestamp 1666464484
transform 1 0 96416 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2019
timestamp 1666464484
transform 1 0 98992 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2020
timestamp 1666464484
transform 1 0 101568 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2021
timestamp 1666464484
transform 1 0 104144 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2022
timestamp 1666464484
transform 1 0 106720 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2023
timestamp 1666464484
transform 1 0 109296 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2024
timestamp 1666464484
transform 1 0 111872 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2025
timestamp 1666464484
transform 1 0 114448 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2026
timestamp 1666464484
transform 1 0 117024 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2027
timestamp 1666464484
transform 1 0 119600 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2028
timestamp 1666464484
transform 1 0 122176 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2029
timestamp 1666464484
transform 1 0 124752 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2030
timestamp 1666464484
transform 1 0 127328 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2031
timestamp 1666464484
transform 1 0 129904 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2032
timestamp 1666464484
transform 1 0 132480 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2033
timestamp 1666464484
transform 1 0 135056 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2034
timestamp 1666464484
transform 1 0 137632 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2035
timestamp 1666464484
transform 1 0 140208 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2036
timestamp 1666464484
transform 1 0 142784 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2037
timestamp 1666464484
transform 1 0 145360 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2038
timestamp 1666464484
transform 1 0 147936 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  _146_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 61548 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _147_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 76360 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _148_
timestamp 1666464484
transform 1 0 64032 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _149_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 74796 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _150_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 74244 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _151_
timestamp 1666464484
transform 1 0 79028 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _152_
timestamp 1666464484
transform 1 0 77280 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _153_
timestamp 1666464484
transform 1 0 76636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _154_
timestamp 1666464484
transform -1 0 81696 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _155_
timestamp 1666464484
transform 1 0 81696 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _156_
timestamp 1666464484
transform 1 0 80592 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _157_
timestamp 1666464484
transform -1 0 82064 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _158_
timestamp 1666464484
transform 1 0 82432 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _159_
timestamp 1666464484
transform 1 0 81880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _160_
timestamp 1666464484
transform 1 0 82432 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _161_
timestamp 1666464484
transform 1 0 81420 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1666464484
transform 1 0 79948 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _163_
timestamp 1666464484
transform -1 0 82064 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _164_
timestamp 1666464484
transform 1 0 81236 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1666464484
transform -1 0 80684 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _166_
timestamp 1666464484
transform 1 0 79672 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _167_
timestamp 1666464484
transform 1 0 79212 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1666464484
transform -1 0 78200 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _169_
timestamp 1666464484
transform -1 0 71760 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _170_
timestamp 1666464484
transform 1 0 70932 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _171_
timestamp 1666464484
transform -1 0 69736 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _172_
timestamp 1666464484
transform -1 0 61916 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _173_
timestamp 1666464484
transform -1 0 69184 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _174_
timestamp 1666464484
transform -1 0 70104 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _175_
timestamp 1666464484
transform -1 0 70104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _176_
timestamp 1666464484
transform -1 0 66976 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _177_
timestamp 1666464484
transform -1 0 68908 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _178_
timestamp 1666464484
transform -1 0 69000 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _179_
timestamp 1666464484
transform -1 0 65228 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _180_
timestamp 1666464484
transform -1 0 54648 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _181_
timestamp 1666464484
transform -1 0 65136 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _182_
timestamp 1666464484
transform 1 0 65504 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _183_
timestamp 1666464484
transform -1 0 65872 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _184_
timestamp 1666464484
transform -1 0 65320 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _185_
timestamp 1666464484
transform -1 0 65320 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _186_
timestamp 1666464484
transform 1 0 58052 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _187_
timestamp 1666464484
transform 1 0 57408 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _188_
timestamp 1666464484
transform 1 0 57132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _189_
timestamp 1666464484
transform 1 0 56764 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _190_
timestamp 1666464484
transform 1 0 55936 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _191_
timestamp 1666464484
transform 1 0 54740 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _192_
timestamp 1666464484
transform -1 0 58880 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _193_
timestamp 1666464484
transform 1 0 58052 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _194_
timestamp 1666464484
transform -1 0 57316 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _195_
timestamp 1666464484
transform 1 0 60812 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _196_
timestamp 1666464484
transform 1 0 60628 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1666464484
transform 1 0 59892 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _198_
timestamp 1666464484
transform -1 0 64032 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _199_
timestamp 1666464484
transform 1 0 63204 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _200_
timestamp 1666464484
transform 1 0 61824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _201_
timestamp 1666464484
transform 1 0 63848 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _202_
timestamp 1666464484
transform 1 0 63296 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _203_
timestamp 1666464484
transform -1 0 62744 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _204_
timestamp 1666464484
transform 1 0 37628 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _205_
timestamp 1666464484
transform -1 0 52440 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _206_
timestamp 1666464484
transform 1 0 51888 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _207_
timestamp 1666464484
transform 1 0 50876 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _208_
timestamp 1666464484
transform -1 0 53728 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _209_
timestamp 1666464484
transform 1 0 52900 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _210_
timestamp 1666464484
transform 1 0 51520 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _211_
timestamp 1666464484
transform -1 0 48576 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _212_
timestamp 1666464484
transform 1 0 29716 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _213_
timestamp 1666464484
transform 1 0 47012 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _214_
timestamp 1666464484
transform 1 0 46828 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _215_
timestamp 1666464484
transform -1 0 48668 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _216_
timestamp 1666464484
transform 1 0 47748 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _217_
timestamp 1666464484
transform -1 0 46460 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _218_
timestamp 1666464484
transform 1 0 42596 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _219_
timestamp 1666464484
transform -1 0 42136 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _220_
timestamp 1666464484
transform 1 0 41860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _221_
timestamp 1666464484
transform -1 0 43700 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _222_
timestamp 1666464484
transform 1 0 43792 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _223_
timestamp 1666464484
transform 1 0 42780 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _224_
timestamp 1666464484
transform 1 0 40756 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _225_
timestamp 1666464484
transform 1 0 40020 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _226_
timestamp 1666464484
transform 1 0 39192 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _227_
timestamp 1666464484
transform 1 0 37904 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _228_
timestamp 1666464484
transform 1 0 37444 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _229_
timestamp 1666464484
transform -1 0 36708 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _230_
timestamp 1666464484
transform 1 0 36156 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _231_
timestamp 1666464484
transform 1 0 35236 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _232_
timestamp 1666464484
transform -1 0 34408 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _233_
timestamp 1666464484
transform 1 0 34960 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _234_
timestamp 1666464484
transform 1 0 33764 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _235_
timestamp 1666464484
transform 1 0 33856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _236_
timestamp 1666464484
transform -1 0 28428 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _237_
timestamp 1666464484
transform 1 0 27324 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _238_
timestamp 1666464484
transform 1 0 27140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _239_
timestamp 1666464484
transform -1 0 28612 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _240_
timestamp 1666464484
transform 1 0 28520 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _241_
timestamp 1666464484
transform -1 0 26036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _242_
timestamp 1666464484
transform 1 0 23920 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _243_
timestamp 1666464484
transform 1 0 24196 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _244_
timestamp 1666464484
transform -1 0 21712 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _245_
timestamp 1666464484
transform 1 0 24564 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _246_
timestamp 1666464484
transform 1 0 22724 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _247_
timestamp 1666464484
transform 1 0 22264 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _248_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5152 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _249_
timestamp 1666464484
transform -1 0 6808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _250_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9200 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _251_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 75256 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _252_
timestamp 1666464484
transform -1 0 76360 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _253_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 62468 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _254_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 60168 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _255_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6716 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _256_
timestamp 1666464484
transform 1 0 32844 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _257_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 22080 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1666464484
transform 1 0 21252 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1666464484
transform 1 0 26404 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1666464484
transform -1 0 28060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp 1666464484
transform 1 0 33212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1666464484
transform 1 0 35788 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1666464484
transform 1 0 38180 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1666464484
transform 1 0 39836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1666464484
transform 1 0 45172 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1666464484
transform 1 0 42412 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _267_
timestamp 1666464484
transform 1 0 49036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1666464484
transform -1 0 50232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _269_
timestamp 1666464484
transform -1 0 46368 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1666464484
transform -1 0 52440 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1666464484
transform 1 0 51612 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _272_
timestamp 1666464484
transform 1 0 62284 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1666464484
transform 1 0 62192 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _274_
timestamp 1666464484
transform -1 0 61548 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _275_
timestamp 1666464484
transform 1 0 58052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _276_
timestamp 1666464484
transform 1 0 55108 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1666464484
transform 1 0 56580 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _278_
timestamp 1666464484
transform 1 0 66240 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _279_
timestamp 1666464484
transform -1 0 66608 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1666464484
transform -1 0 67436 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _281_
timestamp 1666464484
transform 1 0 68816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _282_
timestamp 1666464484
transform 1 0 69552 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _283_
timestamp 1666464484
transform 1 0 70196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _284_
timestamp 1666464484
transform 1 0 79304 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _285_
timestamp 1666464484
transform -1 0 84088 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _286_
timestamp 1666464484
transform -1 0 81512 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _287_
timestamp 1666464484
transform -1 0 81512 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _288_
timestamp 1666464484
transform -1 0 85008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _289_
timestamp 1666464484
transform 1 0 75072 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _290_
timestamp 1666464484
transform 1 0 74060 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _291_
timestamp 1666464484
transform -1 0 6348 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _292_
timestamp 1666464484
transform 1 0 30728 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _293_
timestamp 1666464484
transform -1 0 8096 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _294_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 21988 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _295_
timestamp 1666464484
transform -1 0 23828 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _296_
timestamp 1666464484
transform 1 0 27140 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _297_
timestamp 1666464484
transform 1 0 26220 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _298_
timestamp 1666464484
transform 1 0 32292 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _299_
timestamp 1666464484
transform 1 0 34868 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _300_
timestamp 1666464484
transform 1 0 37444 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _301_
timestamp 1666464484
transform 1 0 38916 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _302_
timestamp 1666464484
transform 1 0 42596 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _303_
timestamp 1666464484
transform 1 0 41584 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _304_
timestamp 1666464484
transform 1 0 47748 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _305_
timestamp 1666464484
transform 1 0 45448 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _306_
timestamp 1666464484
transform 1 0 50600 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _307_
timestamp 1666464484
transform 1 0 50600 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _308_
timestamp 1666464484
transform 1 0 63204 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _309_
timestamp 1666464484
transform 1 0 60904 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _310_
timestamp 1666464484
transform 1 0 59708 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _311_
timestamp 1666464484
transform 1 0 58052 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _312_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 54280 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _313_
timestamp 1666464484
transform 1 0 55660 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _314_
timestamp 1666464484
transform 1 0 65780 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _315_
timestamp 1666464484
transform 1 0 65228 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _316_
timestamp 1666464484
transform 1 0 69368 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _317_
timestamp 1666464484
transform 1 0 70104 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _318_
timestamp 1666464484
transform 1 0 70932 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _319_
timestamp 1666464484
transform 1 0 78476 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _320_
timestamp 1666464484
transform 1 0 81236 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _321_
timestamp 1666464484
transform 1 0 79120 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _322_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 78660 0 1 2176
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _323_
timestamp 1666464484
transform 1 0 79212 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _324_
timestamp 1666464484
transform 1 0 76084 0 1 2176
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _325_
timestamp 1666464484
transform 1 0 73508 0 1 2176
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _326_
timestamp 1666464484
transform -1 0 6072 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_2  _327_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29900 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _328_
timestamp 1666464484
transform 1 0 6532 0 1 2176
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_1  _331_
timestamp 1666464484
transform 1 0 21252 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _332_
timestamp 1666464484
transform 1 0 27140 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _333_
timestamp 1666464484
transform 1 0 32292 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _334_
timestamp 1666464484
transform 1 0 36524 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _335_
timestamp 1666464484
transform 1 0 40388 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _336_
timestamp 1666464484
transform -1 0 44712 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _337_
timestamp 1666464484
transform -1 0 48944 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _338_
timestamp 1666464484
transform -1 0 52440 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _339_
timestamp 1666464484
transform -1 0 57316 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _340_
timestamp 1666464484
transform 1 0 53452 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _341_
timestamp 1666464484
transform 1 0 29716 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _342_
timestamp 1666464484
transform 1 0 33304 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _343_
timestamp 1666464484
transform 1 0 38548 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _344_
timestamp 1666464484
transform 1 0 41768 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _345_
timestamp 1666464484
transform 1 0 45172 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _346_
timestamp 1666464484
transform 1 0 50140 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _347_
timestamp 1666464484
transform 1 0 54188 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _348_
timestamp 1666464484
transform 1 0 58788 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _349_
timestamp 1666464484
transform 1 0 6532 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _350_
timestamp 1666464484
transform 1 0 9752 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _351_
timestamp 1666464484
transform 1 0 23828 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _352_
timestamp 1666464484
transform 1 0 17296 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _353_
timestamp 1666464484
transform 1 0 20608 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _354_
timestamp 1666464484
transform 1 0 39652 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _355_
timestamp 1666464484
transform 1 0 43424 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _356_
timestamp 1666464484
transform 1 0 47012 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _357_
timestamp 1666464484
transform 1 0 51428 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _358_
timestamp 1666464484
transform -1 0 55936 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _359_
timestamp 1666464484
transform -1 0 59708 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _360_
timestamp 1666464484
transform -1 0 64032 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _361_
timestamp 1666464484
transform -1 0 69000 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _362_
timestamp 1666464484
transform -1 0 67896 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _363_
timestamp 1666464484
transform -1 0 73968 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _364_
timestamp 1666464484
transform -1 0 82432 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _365_
timestamp 1666464484
transform -1 0 85284 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _366_
timestamp 1666464484
transform -1 0 90068 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _367_
timestamp 1666464484
transform -1 0 93380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _368_
timestamp 1666464484
transform -1 0 97796 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _369_
timestamp 1666464484
transform -1 0 102212 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _370_
timestamp 1666464484
transform -1 0 105708 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _371_
timestamp 1666464484
transform -1 0 110676 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _372_
timestamp 1666464484
transform -1 0 114080 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _373_
timestamp 1666464484
transform -1 0 118220 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _374_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 122820 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _375_
timestamp 1666464484
transform -1 0 126776 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _376_
timestamp 1666464484
transform -1 0 130548 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _377_
timestamp 1666464484
transform -1 0 120980 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _378_
timestamp 1666464484
transform -1 0 112792 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _379_
timestamp 1666464484
transform -1 0 106260 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _380_
timestamp 1666464484
transform 1 0 95036 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _381_
timestamp 1666464484
transform 1 0 45908 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _382_
timestamp 1666464484
transform 1 0 21160 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _383_
timestamp 1666464484
transform 1 0 25760 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _384_
timestamp 1666464484
transform 1 0 30544 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _385_
timestamp 1666464484
transform 1 0 35880 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _386_
timestamp 1666464484
transform 1 0 41032 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _387_
timestamp 1666464484
transform 1 0 44528 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _388_
timestamp 1666464484
transform 1 0 48944 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _389_
timestamp 1666464484
transform 1 0 52624 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _390_
timestamp 1666464484
transform 1 0 56856 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _391_
timestamp 1666464484
transform 1 0 60812 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _392_
timestamp 1666464484
transform 1 0 65780 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _393_
timestamp 1666464484
transform 1 0 69368 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _394_
timestamp 1666464484
transform 1 0 75256 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _395_
timestamp 1666464484
transform 1 0 78384 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _396_
timestamp 1666464484
transform 1 0 83812 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _397_
timestamp 1666464484
transform 1 0 86204 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _398_
timestamp 1666464484
transform 1 0 90252 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _399_
timestamp 1666464484
transform 1 0 94852 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _400_
timestamp 1666464484
transform 1 0 99268 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _401_
timestamp 1666464484
transform 1 0 103316 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _402_
timestamp 1666464484
transform -1 0 107088 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _403_
timestamp 1666464484
transform -1 0 111044 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _404_
timestamp 1666464484
transform -1 0 115276 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _405_
timestamp 1666464484
transform -1 0 132296 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _406_
timestamp 1666464484
transform -1 0 123464 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _407_
timestamp 1666464484
transform -1 0 136068 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _408_
timestamp 1666464484
transform -1 0 137908 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _409_
timestamp 1666464484
transform -1 0 139932 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _410_
timestamp 1666464484
transform -1 0 141680 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _411_
timestamp 1666464484
transform -1 0 143888 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _412_
timestamp 1666464484
transform -1 0 146372 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _413_
timestamp 1666464484
transform 1 0 8188 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _414_
timestamp 1666464484
transform 1 0 19688 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _415_
timestamp 1666464484
transform 1 0 25116 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _416_
timestamp 1666464484
transform 1 0 19044 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _417_
timestamp 1666464484
transform 1 0 35144 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _418_
timestamp 1666464484
transform 1 0 21988 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _419_
timestamp 1666464484
transform 1 0 26312 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _420_
timestamp 1666464484
transform 1 0 32292 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_io_wbs_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 43700 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_io_wbs_clk
timestamp 1666464484
transform -1 0 38272 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_io_wbs_clk
timestamp 1666464484
transform -1 0 36984 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_io_wbs_clk
timestamp 1666464484
transform 1 0 46828 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_io_wbs_clk
timestamp 1666464484
transform 1 0 47748 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1666464484
transform -1 0 6808 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1666464484
transform -1 0 36156 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1666464484
transform -1 0 37996 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1666464484
transform -1 0 40296 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1666464484
transform -1 0 41676 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1666464484
transform -1 0 44344 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1666464484
transform -1 0 45540 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1666464484
transform -1 0 47196 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1666464484
transform -1 0 49588 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1666464484
transform -1 0 50876 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1666464484
transform -1 0 52256 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1666464484
transform -1 0 10396 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1666464484
transform -1 0 55200 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1666464484
transform -1 0 56580 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1666464484
transform -1 0 58236 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1666464484
transform -1 0 60904 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1666464484
transform -1 0 62744 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1666464484
transform -1 0 63480 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1666464484
transform -1 0 65596 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1666464484
transform -1 0 67436 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1666464484
transform -1 0 69276 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1666464484
transform -1 0 71116 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1666464484
transform -1 0 14076 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1666464484
transform -1 0 72956 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1666464484
transform -1 0 74796 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1666464484
transform -1 0 17848 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1666464484
transform -1 0 21436 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1666464484
transform -1 0 23552 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1666464484
transform -1 0 26956 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1666464484
transform -1 0 29256 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1666464484
transform -1 0 32476 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1666464484
transform -1 0 34316 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1666464484
transform -1 0 80592 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input34
timestamp 1666464484
transform 1 0 108560 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1666464484
transform 1 0 111044 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input36
timestamp 1666464484
transform 1 0 112884 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input37
timestamp 1666464484
transform 1 0 114724 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1666464484
transform -1 0 116564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1666464484
transform -1 0 118404 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input40
timestamp 1666464484
transform 1 0 119876 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input41
timestamp 1666464484
transform 1 0 121440 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input42
timestamp 1666464484
transform -1 0 124292 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input43
timestamp 1666464484
transform 1 0 125764 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input44
timestamp 1666464484
transform -1 0 84916 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input45
timestamp 1666464484
transform 1 0 127604 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 1666464484
transform 1 0 129076 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1666464484
transform -1 0 131284 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input48
timestamp 1666464484
transform -1 0 133124 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input49
timestamp 1666464484
transform 1 0 134320 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1666464484
transform -1 0 136528 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1666464484
transform -1 0 138368 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input52
timestamp 1666464484
transform 1 0 140484 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input53
timestamp 1666464484
transform -1 0 142324 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input54
timestamp 1666464484
transform 1 0 143796 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input55
timestamp 1666464484
transform -1 0 87492 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 1666464484
transform 1 0 145636 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input57
timestamp 1666464484
transform 1 0 147200 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input58
timestamp 1666464484
transform -1 0 90804 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1666464484
transform -1 0 94484 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input60
timestamp 1666464484
transform -1 0 97060 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input61
timestamp 1666464484
transform 1 0 100004 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input62
timestamp 1666464484
transform -1 0 102948 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input63
timestamp 1666464484
transform 1 0 105156 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input64
timestamp 1666464484
transform -1 0 107364 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1666464484
transform -1 0 57592 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input66
timestamp 1666464484
transform 1 0 61916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input67
timestamp 1666464484
transform -1 0 21528 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1666464484
transform 1 0 26312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1666464484
transform 1 0 32936 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1666464484
transform 1 0 37444 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input71
timestamp 1666464484
transform -1 0 41216 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input72
timestamp 1666464484
transform -1 0 46276 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1666464484
transform 1 0 49496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1666464484
transform 1 0 53636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1666464484
transform -1 0 5612 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input76
timestamp 1666464484
transform 1 0 14260 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input77
timestamp 1666464484
transform 1 0 60536 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input78
timestamp 1666464484
transform 1 0 64492 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input79
timestamp 1666464484
transform 1 0 68816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input80
timestamp 1666464484
transform 1 0 73508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input81
timestamp 1666464484
transform -1 0 77464 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input82
timestamp 1666464484
transform -1 0 83260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input83
timestamp 1666464484
transform -1 0 85744 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input84
timestamp 1666464484
transform 1 0 89516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1666464484
transform 1 0 94116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input86
timestamp 1666464484
transform 1 0 97796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input87
timestamp 1666464484
transform 1 0 19412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input88
timestamp 1666464484
transform 1 0 101936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input89
timestamp 1666464484
transform 1 0 106076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input90
timestamp 1666464484
transform 1 0 110308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input91
timestamp 1666464484
transform 1 0 114724 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input92
timestamp 1666464484
transform 1 0 118496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input93
timestamp 1666464484
transform 1 0 122636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input94
timestamp 1666464484
transform 1 0 126776 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input95
timestamp 1666464484
transform 1 0 130916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input96
timestamp 1666464484
transform 1 0 135332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input97
timestamp 1666464484
transform 1 0 139196 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input98
timestamp 1666464484
transform -1 0 25024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input99
timestamp 1666464484
transform 1 0 143336 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input100
timestamp 1666464484
transform -1 0 147752 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input101
timestamp 1666464484
transform 1 0 30636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input102
timestamp 1666464484
transform 1 0 35696 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input103
timestamp 1666464484
transform 1 0 40020 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input104
timestamp 1666464484
transform 1 0 44160 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input105
timestamp 1666464484
transform -1 0 48576 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input106
timestamp 1666464484
transform 1 0 52900 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input107
timestamp 1666464484
transform 1 0 56396 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input108
timestamp 1666464484
transform 1 0 6716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input109
timestamp 1666464484
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input110
timestamp 1666464484
transform 1 0 20424 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input111
timestamp 1666464484
transform -1 0 25944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input112
timestamp 1666464484
transform -1 0 31832 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input113
timestamp 1666464484
transform 1 0 8096 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input114
timestamp 1666464484
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1666464484
transform -1 0 4968 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1666464484
transform -1 0 8648 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1666464484
transform -1 0 12328 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1666464484
transform -1 0 16008 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1666464484
transform -1 0 19780 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1666464484
transform -1 0 22448 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1666464484
transform -1 0 25208 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1666464484
transform -1 0 27968 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1666464484
transform -1 0 30728 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1666464484
transform 1 0 77556 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1666464484
transform 1 0 80960 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1666464484
transform 1 0 85284 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1666464484
transform -1 0 89332 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1666464484
transform 1 0 92276 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1666464484
transform -1 0 95956 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1666464484
transform -1 0 98532 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1666464484
transform 1 0 100740 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1666464484
transform 1 0 103040 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1666464484
transform -1 0 5888 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1666464484
transform -1 0 34408 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1666464484
transform -1 0 36984 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1666464484
transform -1 0 39468 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1666464484
transform 1 0 40020 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1666464484
transform -1 0 42688 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1666464484
transform -1 0 44160 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1666464484
transform -1 0 46368 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1666464484
transform 1 0 46920 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1666464484
transform -1 0 49864 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1666464484
transform -1 0 51244 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1666464484
transform -1 0 9568 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1666464484
transform -1 0 53728 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1666464484
transform -1 0 55016 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1666464484
transform 1 0 56028 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1666464484
transform -1 0 59892 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1666464484
transform 1 0 60076 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 1666464484
transform -1 0 62928 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 1666464484
transform -1 0 64768 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 1666464484
transform -1 0 66608 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 1666464484
transform -1 0 68448 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 1666464484
transform -1 0 70288 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 1666464484
transform -1 0 13248 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 1666464484
transform -1 0 72496 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 1666464484
transform -1 0 74704 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 1666464484
transform -1 0 17204 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 1666464484
transform -1 0 20608 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 1666464484
transform -1 0 23368 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 1666464484
transform -1 0 26128 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 1666464484
transform -1 0 29164 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 1666464484
transform -1 0 31648 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1666464484
transform -1 0 33488 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1666464484
transform -1 0 79028 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1666464484
transform 1 0 107732 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1666464484
transform 1 0 109572 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1666464484
transform 1 0 112148 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1666464484
transform 1 0 113620 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1666464484
transform 1 0 115460 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1666464484
transform 1 0 117300 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1666464484
transform -1 0 119140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1666464484
transform -1 0 121716 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1666464484
transform 1 0 123188 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1666464484
transform 1 0 125028 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 1666464484
transform -1 0 83168 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 1666464484
transform 1 0 126500 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1666464484
transform 1 0 128340 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 1666464484
transform 1 0 130180 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 1666464484
transform 1 0 131652 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 1666464484
transform 1 0 133492 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 1666464484
transform 1 0 135332 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 1666464484
transform 1 0 137080 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 1666464484
transform 1 0 138920 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 1666464484
transform 1 0 141220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 1666464484
transform 1 0 143060 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 1666464484
transform -1 0 86756 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 1666464484
transform 1 0 144532 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 1666464484
transform 1 0 146372 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 1666464484
transform 1 0 89240 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 1666464484
transform 1 0 93012 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 1666464484
transform -1 0 96048 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1666464484
transform 1 0 98440 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 1666464484
transform 1 0 101200 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 1666464484
transform 1 0 104420 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1666464484
transform -1 0 106444 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 1666464484
transform -1 0 2944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1666464484
transform -1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 1666464484
transform 1 0 59156 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 1666464484
transform 1 0 63296 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 1666464484
transform 1 0 67528 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1666464484
transform 1 0 72404 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 1666464484
transform 1 0 75716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1666464484
transform 1 0 77832 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output205
timestamp 1666464484
transform -1 0 84364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 1666464484
transform 1 0 88136 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 1666464484
transform 1 0 92276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 1666464484
transform 1 0 96692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 1666464484
transform -1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1666464484
transform 1 0 100556 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 1666464484
transform 1 0 104696 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1666464484
transform 1 0 109572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 1666464484
transform 1 0 112976 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 1666464484
transform 1 0 117300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 1666464484
transform 1 0 121256 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output216
timestamp 1666464484
transform 1 0 125396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output217
timestamp 1666464484
transform 1 0 130180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 1666464484
transform 1 0 133676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output219
timestamp 1666464484
transform 1 0 137908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 1666464484
transform -1 0 23644 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 1666464484
transform 1 0 141956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 1666464484
transform 1 0 146096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 1666464484
transform 1 0 28796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output224
timestamp 1666464484
transform 1 0 34960 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 1666464484
transform 1 0 38640 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output226
timestamp 1666464484
transform 1 0 41768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 1666464484
transform 1 0 46736 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output228
timestamp 1666464484
transform 1 0 50876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output229
timestamp 1666464484
transform 1 0 53360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 1666464484
transform -1 0 4048 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output231
timestamp 1666464484
transform 1 0 76360 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output232
timestamp 1666464484
transform -1 0 7728 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output233
timestamp 1666464484
transform -1 0 11224 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output234
timestamp 1666464484
transform -1 0 15088 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output235
timestamp 1666464484
transform -1 0 18768 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output236
timestamp 1666464484
transform 1 0 80040 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output237
timestamp 1666464484
transform 1 0 83812 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output238
timestamp 1666464484
transform -1 0 88228 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output239
timestamp 1666464484
transform 1 0 91540 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  wb_memory_240 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 3036 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wb_memory_241
timestamp 1666464484
transform 1 0 74612 0 -1 36992
box -38 -48 314 592
<< labels >>
flabel metal2 s 4526 39200 4582 40000 0 FreeSans 224 90 0 0 addr_mem0[0]
port 0 nsew signal tristate
flabel metal2 s 8206 39200 8262 40000 0 FreeSans 224 90 0 0 addr_mem0[1]
port 1 nsew signal tristate
flabel metal2 s 11886 39200 11942 40000 0 FreeSans 224 90 0 0 addr_mem0[2]
port 2 nsew signal tristate
flabel metal2 s 15566 39200 15622 40000 0 FreeSans 224 90 0 0 addr_mem0[3]
port 3 nsew signal tristate
flabel metal2 s 19246 39200 19302 40000 0 FreeSans 224 90 0 0 addr_mem0[4]
port 4 nsew signal tristate
flabel metal2 s 22006 39200 22062 40000 0 FreeSans 224 90 0 0 addr_mem0[5]
port 5 nsew signal tristate
flabel metal2 s 24766 39200 24822 40000 0 FreeSans 224 90 0 0 addr_mem0[6]
port 6 nsew signal tristate
flabel metal2 s 27526 39200 27582 40000 0 FreeSans 224 90 0 0 addr_mem0[7]
port 7 nsew signal tristate
flabel metal2 s 30286 39200 30342 40000 0 FreeSans 224 90 0 0 addr_mem0[8]
port 8 nsew signal tristate
flabel metal2 s 77206 39200 77262 40000 0 FreeSans 224 90 0 0 addr_mem1[0]
port 9 nsew signal tristate
flabel metal2 s 80886 39200 80942 40000 0 FreeSans 224 90 0 0 addr_mem1[1]
port 10 nsew signal tristate
flabel metal2 s 84566 39200 84622 40000 0 FreeSans 224 90 0 0 addr_mem1[2]
port 11 nsew signal tristate
flabel metal2 s 88246 39200 88302 40000 0 FreeSans 224 90 0 0 addr_mem1[3]
port 12 nsew signal tristate
flabel metal2 s 91926 39200 91982 40000 0 FreeSans 224 90 0 0 addr_mem1[4]
port 13 nsew signal tristate
flabel metal2 s 94686 39200 94742 40000 0 FreeSans 224 90 0 0 addr_mem1[5]
port 14 nsew signal tristate
flabel metal2 s 97446 39200 97502 40000 0 FreeSans 224 90 0 0 addr_mem1[6]
port 15 nsew signal tristate
flabel metal2 s 100206 39200 100262 40000 0 FreeSans 224 90 0 0 addr_mem1[7]
port 16 nsew signal tristate
flabel metal2 s 102966 39200 103022 40000 0 FreeSans 224 90 0 0 addr_mem1[8]
port 17 nsew signal tristate
flabel metal2 s 2686 39200 2742 40000 0 FreeSans 224 90 0 0 csb_mem0
port 18 nsew signal tristate
flabel metal2 s 75366 39200 75422 40000 0 FreeSans 224 90 0 0 csb_mem1
port 19 nsew signal tristate
flabel metal2 s 5446 39200 5502 40000 0 FreeSans 224 90 0 0 din_mem0[0]
port 20 nsew signal tristate
flabel metal2 s 34886 39200 34942 40000 0 FreeSans 224 90 0 0 din_mem0[10]
port 21 nsew signal tristate
flabel metal2 s 36726 39200 36782 40000 0 FreeSans 224 90 0 0 din_mem0[11]
port 22 nsew signal tristate
flabel metal2 s 38566 39200 38622 40000 0 FreeSans 224 90 0 0 din_mem0[12]
port 23 nsew signal tristate
flabel metal2 s 40406 39200 40462 40000 0 FreeSans 224 90 0 0 din_mem0[13]
port 24 nsew signal tristate
flabel metal2 s 42246 39200 42302 40000 0 FreeSans 224 90 0 0 din_mem0[14]
port 25 nsew signal tristate
flabel metal2 s 44086 39200 44142 40000 0 FreeSans 224 90 0 0 din_mem0[15]
port 26 nsew signal tristate
flabel metal2 s 45926 39200 45982 40000 0 FreeSans 224 90 0 0 din_mem0[16]
port 27 nsew signal tristate
flabel metal2 s 47766 39200 47822 40000 0 FreeSans 224 90 0 0 din_mem0[17]
port 28 nsew signal tristate
flabel metal2 s 49606 39200 49662 40000 0 FreeSans 224 90 0 0 din_mem0[18]
port 29 nsew signal tristate
flabel metal2 s 51446 39200 51502 40000 0 FreeSans 224 90 0 0 din_mem0[19]
port 30 nsew signal tristate
flabel metal2 s 9126 39200 9182 40000 0 FreeSans 224 90 0 0 din_mem0[1]
port 31 nsew signal tristate
flabel metal2 s 53286 39200 53342 40000 0 FreeSans 224 90 0 0 din_mem0[20]
port 32 nsew signal tristate
flabel metal2 s 55126 39200 55182 40000 0 FreeSans 224 90 0 0 din_mem0[21]
port 33 nsew signal tristate
flabel metal2 s 56966 39200 57022 40000 0 FreeSans 224 90 0 0 din_mem0[22]
port 34 nsew signal tristate
flabel metal2 s 58806 39200 58862 40000 0 FreeSans 224 90 0 0 din_mem0[23]
port 35 nsew signal tristate
flabel metal2 s 60646 39200 60702 40000 0 FreeSans 224 90 0 0 din_mem0[24]
port 36 nsew signal tristate
flabel metal2 s 62486 39200 62542 40000 0 FreeSans 224 90 0 0 din_mem0[25]
port 37 nsew signal tristate
flabel metal2 s 64326 39200 64382 40000 0 FreeSans 224 90 0 0 din_mem0[26]
port 38 nsew signal tristate
flabel metal2 s 66166 39200 66222 40000 0 FreeSans 224 90 0 0 din_mem0[27]
port 39 nsew signal tristate
flabel metal2 s 68006 39200 68062 40000 0 FreeSans 224 90 0 0 din_mem0[28]
port 40 nsew signal tristate
flabel metal2 s 69846 39200 69902 40000 0 FreeSans 224 90 0 0 din_mem0[29]
port 41 nsew signal tristate
flabel metal2 s 12806 39200 12862 40000 0 FreeSans 224 90 0 0 din_mem0[2]
port 42 nsew signal tristate
flabel metal2 s 71686 39200 71742 40000 0 FreeSans 224 90 0 0 din_mem0[30]
port 43 nsew signal tristate
flabel metal2 s 73526 39200 73582 40000 0 FreeSans 224 90 0 0 din_mem0[31]
port 44 nsew signal tristate
flabel metal2 s 16486 39200 16542 40000 0 FreeSans 224 90 0 0 din_mem0[3]
port 45 nsew signal tristate
flabel metal2 s 20166 39200 20222 40000 0 FreeSans 224 90 0 0 din_mem0[4]
port 46 nsew signal tristate
flabel metal2 s 22926 39200 22982 40000 0 FreeSans 224 90 0 0 din_mem0[5]
port 47 nsew signal tristate
flabel metal2 s 25686 39200 25742 40000 0 FreeSans 224 90 0 0 din_mem0[6]
port 48 nsew signal tristate
flabel metal2 s 28446 39200 28502 40000 0 FreeSans 224 90 0 0 din_mem0[7]
port 49 nsew signal tristate
flabel metal2 s 31206 39200 31262 40000 0 FreeSans 224 90 0 0 din_mem0[8]
port 50 nsew signal tristate
flabel metal2 s 33046 39200 33102 40000 0 FreeSans 224 90 0 0 din_mem0[9]
port 51 nsew signal tristate
flabel metal2 s 78126 39200 78182 40000 0 FreeSans 224 90 0 0 din_mem1[0]
port 52 nsew signal tristate
flabel metal2 s 107566 39200 107622 40000 0 FreeSans 224 90 0 0 din_mem1[10]
port 53 nsew signal tristate
flabel metal2 s 109406 39200 109462 40000 0 FreeSans 224 90 0 0 din_mem1[11]
port 54 nsew signal tristate
flabel metal2 s 111246 39200 111302 40000 0 FreeSans 224 90 0 0 din_mem1[12]
port 55 nsew signal tristate
flabel metal2 s 113086 39200 113142 40000 0 FreeSans 224 90 0 0 din_mem1[13]
port 56 nsew signal tristate
flabel metal2 s 114926 39200 114982 40000 0 FreeSans 224 90 0 0 din_mem1[14]
port 57 nsew signal tristate
flabel metal2 s 116766 39200 116822 40000 0 FreeSans 224 90 0 0 din_mem1[15]
port 58 nsew signal tristate
flabel metal2 s 118606 39200 118662 40000 0 FreeSans 224 90 0 0 din_mem1[16]
port 59 nsew signal tristate
flabel metal2 s 120446 39200 120502 40000 0 FreeSans 224 90 0 0 din_mem1[17]
port 60 nsew signal tristate
flabel metal2 s 122286 39200 122342 40000 0 FreeSans 224 90 0 0 din_mem1[18]
port 61 nsew signal tristate
flabel metal2 s 124126 39200 124182 40000 0 FreeSans 224 90 0 0 din_mem1[19]
port 62 nsew signal tristate
flabel metal2 s 81806 39200 81862 40000 0 FreeSans 224 90 0 0 din_mem1[1]
port 63 nsew signal tristate
flabel metal2 s 125966 39200 126022 40000 0 FreeSans 224 90 0 0 din_mem1[20]
port 64 nsew signal tristate
flabel metal2 s 127806 39200 127862 40000 0 FreeSans 224 90 0 0 din_mem1[21]
port 65 nsew signal tristate
flabel metal2 s 129646 39200 129702 40000 0 FreeSans 224 90 0 0 din_mem1[22]
port 66 nsew signal tristate
flabel metal2 s 131486 39200 131542 40000 0 FreeSans 224 90 0 0 din_mem1[23]
port 67 nsew signal tristate
flabel metal2 s 133326 39200 133382 40000 0 FreeSans 224 90 0 0 din_mem1[24]
port 68 nsew signal tristate
flabel metal2 s 135166 39200 135222 40000 0 FreeSans 224 90 0 0 din_mem1[25]
port 69 nsew signal tristate
flabel metal2 s 137006 39200 137062 40000 0 FreeSans 224 90 0 0 din_mem1[26]
port 70 nsew signal tristate
flabel metal2 s 138846 39200 138902 40000 0 FreeSans 224 90 0 0 din_mem1[27]
port 71 nsew signal tristate
flabel metal2 s 140686 39200 140742 40000 0 FreeSans 224 90 0 0 din_mem1[28]
port 72 nsew signal tristate
flabel metal2 s 142526 39200 142582 40000 0 FreeSans 224 90 0 0 din_mem1[29]
port 73 nsew signal tristate
flabel metal2 s 85486 39200 85542 40000 0 FreeSans 224 90 0 0 din_mem1[2]
port 74 nsew signal tristate
flabel metal2 s 144366 39200 144422 40000 0 FreeSans 224 90 0 0 din_mem1[30]
port 75 nsew signal tristate
flabel metal2 s 146206 39200 146262 40000 0 FreeSans 224 90 0 0 din_mem1[31]
port 76 nsew signal tristate
flabel metal2 s 89166 39200 89222 40000 0 FreeSans 224 90 0 0 din_mem1[3]
port 77 nsew signal tristate
flabel metal2 s 92846 39200 92902 40000 0 FreeSans 224 90 0 0 din_mem1[4]
port 78 nsew signal tristate
flabel metal2 s 95606 39200 95662 40000 0 FreeSans 224 90 0 0 din_mem1[5]
port 79 nsew signal tristate
flabel metal2 s 98366 39200 98422 40000 0 FreeSans 224 90 0 0 din_mem1[6]
port 80 nsew signal tristate
flabel metal2 s 101126 39200 101182 40000 0 FreeSans 224 90 0 0 din_mem1[7]
port 81 nsew signal tristate
flabel metal2 s 103886 39200 103942 40000 0 FreeSans 224 90 0 0 din_mem1[8]
port 82 nsew signal tristate
flabel metal2 s 105726 39200 105782 40000 0 FreeSans 224 90 0 0 din_mem1[9]
port 83 nsew signal tristate
flabel metal2 s 6366 39200 6422 40000 0 FreeSans 224 90 0 0 dout_mem0[0]
port 84 nsew signal input
flabel metal2 s 35806 39200 35862 40000 0 FreeSans 224 90 0 0 dout_mem0[10]
port 85 nsew signal input
flabel metal2 s 37646 39200 37702 40000 0 FreeSans 224 90 0 0 dout_mem0[11]
port 86 nsew signal input
flabel metal2 s 39486 39200 39542 40000 0 FreeSans 224 90 0 0 dout_mem0[12]
port 87 nsew signal input
flabel metal2 s 41326 39200 41382 40000 0 FreeSans 224 90 0 0 dout_mem0[13]
port 88 nsew signal input
flabel metal2 s 43166 39200 43222 40000 0 FreeSans 224 90 0 0 dout_mem0[14]
port 89 nsew signal input
flabel metal2 s 45006 39200 45062 40000 0 FreeSans 224 90 0 0 dout_mem0[15]
port 90 nsew signal input
flabel metal2 s 46846 39200 46902 40000 0 FreeSans 224 90 0 0 dout_mem0[16]
port 91 nsew signal input
flabel metal2 s 48686 39200 48742 40000 0 FreeSans 224 90 0 0 dout_mem0[17]
port 92 nsew signal input
flabel metal2 s 50526 39200 50582 40000 0 FreeSans 224 90 0 0 dout_mem0[18]
port 93 nsew signal input
flabel metal2 s 52366 39200 52422 40000 0 FreeSans 224 90 0 0 dout_mem0[19]
port 94 nsew signal input
flabel metal2 s 10046 39200 10102 40000 0 FreeSans 224 90 0 0 dout_mem0[1]
port 95 nsew signal input
flabel metal2 s 54206 39200 54262 40000 0 FreeSans 224 90 0 0 dout_mem0[20]
port 96 nsew signal input
flabel metal2 s 56046 39200 56102 40000 0 FreeSans 224 90 0 0 dout_mem0[21]
port 97 nsew signal input
flabel metal2 s 57886 39200 57942 40000 0 FreeSans 224 90 0 0 dout_mem0[22]
port 98 nsew signal input
flabel metal2 s 59726 39200 59782 40000 0 FreeSans 224 90 0 0 dout_mem0[23]
port 99 nsew signal input
flabel metal2 s 61566 39200 61622 40000 0 FreeSans 224 90 0 0 dout_mem0[24]
port 100 nsew signal input
flabel metal2 s 63406 39200 63462 40000 0 FreeSans 224 90 0 0 dout_mem0[25]
port 101 nsew signal input
flabel metal2 s 65246 39200 65302 40000 0 FreeSans 224 90 0 0 dout_mem0[26]
port 102 nsew signal input
flabel metal2 s 67086 39200 67142 40000 0 FreeSans 224 90 0 0 dout_mem0[27]
port 103 nsew signal input
flabel metal2 s 68926 39200 68982 40000 0 FreeSans 224 90 0 0 dout_mem0[28]
port 104 nsew signal input
flabel metal2 s 70766 39200 70822 40000 0 FreeSans 224 90 0 0 dout_mem0[29]
port 105 nsew signal input
flabel metal2 s 13726 39200 13782 40000 0 FreeSans 224 90 0 0 dout_mem0[2]
port 106 nsew signal input
flabel metal2 s 72606 39200 72662 40000 0 FreeSans 224 90 0 0 dout_mem0[30]
port 107 nsew signal input
flabel metal2 s 74446 39200 74502 40000 0 FreeSans 224 90 0 0 dout_mem0[31]
port 108 nsew signal input
flabel metal2 s 17406 39200 17462 40000 0 FreeSans 224 90 0 0 dout_mem0[3]
port 109 nsew signal input
flabel metal2 s 21086 39200 21142 40000 0 FreeSans 224 90 0 0 dout_mem0[4]
port 110 nsew signal input
flabel metal2 s 23846 39200 23902 40000 0 FreeSans 224 90 0 0 dout_mem0[5]
port 111 nsew signal input
flabel metal2 s 26606 39200 26662 40000 0 FreeSans 224 90 0 0 dout_mem0[6]
port 112 nsew signal input
flabel metal2 s 29366 39200 29422 40000 0 FreeSans 224 90 0 0 dout_mem0[7]
port 113 nsew signal input
flabel metal2 s 32126 39200 32182 40000 0 FreeSans 224 90 0 0 dout_mem0[8]
port 114 nsew signal input
flabel metal2 s 33966 39200 34022 40000 0 FreeSans 224 90 0 0 dout_mem0[9]
port 115 nsew signal input
flabel metal2 s 79046 39200 79102 40000 0 FreeSans 224 90 0 0 dout_mem1[0]
port 116 nsew signal input
flabel metal2 s 108486 39200 108542 40000 0 FreeSans 224 90 0 0 dout_mem1[10]
port 117 nsew signal input
flabel metal2 s 110326 39200 110382 40000 0 FreeSans 224 90 0 0 dout_mem1[11]
port 118 nsew signal input
flabel metal2 s 112166 39200 112222 40000 0 FreeSans 224 90 0 0 dout_mem1[12]
port 119 nsew signal input
flabel metal2 s 114006 39200 114062 40000 0 FreeSans 224 90 0 0 dout_mem1[13]
port 120 nsew signal input
flabel metal2 s 115846 39200 115902 40000 0 FreeSans 224 90 0 0 dout_mem1[14]
port 121 nsew signal input
flabel metal2 s 117686 39200 117742 40000 0 FreeSans 224 90 0 0 dout_mem1[15]
port 122 nsew signal input
flabel metal2 s 119526 39200 119582 40000 0 FreeSans 224 90 0 0 dout_mem1[16]
port 123 nsew signal input
flabel metal2 s 121366 39200 121422 40000 0 FreeSans 224 90 0 0 dout_mem1[17]
port 124 nsew signal input
flabel metal2 s 123206 39200 123262 40000 0 FreeSans 224 90 0 0 dout_mem1[18]
port 125 nsew signal input
flabel metal2 s 125046 39200 125102 40000 0 FreeSans 224 90 0 0 dout_mem1[19]
port 126 nsew signal input
flabel metal2 s 82726 39200 82782 40000 0 FreeSans 224 90 0 0 dout_mem1[1]
port 127 nsew signal input
flabel metal2 s 126886 39200 126942 40000 0 FreeSans 224 90 0 0 dout_mem1[20]
port 128 nsew signal input
flabel metal2 s 128726 39200 128782 40000 0 FreeSans 224 90 0 0 dout_mem1[21]
port 129 nsew signal input
flabel metal2 s 130566 39200 130622 40000 0 FreeSans 224 90 0 0 dout_mem1[22]
port 130 nsew signal input
flabel metal2 s 132406 39200 132462 40000 0 FreeSans 224 90 0 0 dout_mem1[23]
port 131 nsew signal input
flabel metal2 s 134246 39200 134302 40000 0 FreeSans 224 90 0 0 dout_mem1[24]
port 132 nsew signal input
flabel metal2 s 136086 39200 136142 40000 0 FreeSans 224 90 0 0 dout_mem1[25]
port 133 nsew signal input
flabel metal2 s 137926 39200 137982 40000 0 FreeSans 224 90 0 0 dout_mem1[26]
port 134 nsew signal input
flabel metal2 s 139766 39200 139822 40000 0 FreeSans 224 90 0 0 dout_mem1[27]
port 135 nsew signal input
flabel metal2 s 141606 39200 141662 40000 0 FreeSans 224 90 0 0 dout_mem1[28]
port 136 nsew signal input
flabel metal2 s 143446 39200 143502 40000 0 FreeSans 224 90 0 0 dout_mem1[29]
port 137 nsew signal input
flabel metal2 s 86406 39200 86462 40000 0 FreeSans 224 90 0 0 dout_mem1[2]
port 138 nsew signal input
flabel metal2 s 145286 39200 145342 40000 0 FreeSans 224 90 0 0 dout_mem1[30]
port 139 nsew signal input
flabel metal2 s 147126 39200 147182 40000 0 FreeSans 224 90 0 0 dout_mem1[31]
port 140 nsew signal input
flabel metal2 s 90086 39200 90142 40000 0 FreeSans 224 90 0 0 dout_mem1[3]
port 141 nsew signal input
flabel metal2 s 93766 39200 93822 40000 0 FreeSans 224 90 0 0 dout_mem1[4]
port 142 nsew signal input
flabel metal2 s 96526 39200 96582 40000 0 FreeSans 224 90 0 0 dout_mem1[5]
port 143 nsew signal input
flabel metal2 s 99286 39200 99342 40000 0 FreeSans 224 90 0 0 dout_mem1[6]
port 144 nsew signal input
flabel metal2 s 102046 39200 102102 40000 0 FreeSans 224 90 0 0 dout_mem1[7]
port 145 nsew signal input
flabel metal2 s 104806 39200 104862 40000 0 FreeSans 224 90 0 0 dout_mem1[8]
port 146 nsew signal input
flabel metal2 s 106646 39200 106702 40000 0 FreeSans 224 90 0 0 dout_mem1[9]
port 147 nsew signal input
flabel metal2 s 2502 0 2558 800 0 FreeSans 224 90 0 0 io_wbs_ack
port 148 nsew signal tristate
flabel metal2 s 10782 0 10838 800 0 FreeSans 224 90 0 0 io_wbs_adr[0]
port 149 nsew signal input
flabel metal2 s 57702 0 57758 800 0 FreeSans 224 90 0 0 io_wbs_adr[10]
port 150 nsew signal input
flabel metal2 s 61842 0 61898 800 0 FreeSans 224 90 0 0 io_wbs_adr[11]
port 151 nsew signal input
flabel metal2 s 65982 0 66038 800 0 FreeSans 224 90 0 0 io_wbs_adr[12]
port 152 nsew signal input
flabel metal2 s 70122 0 70178 800 0 FreeSans 224 90 0 0 io_wbs_adr[13]
port 153 nsew signal input
flabel metal2 s 74262 0 74318 800 0 FreeSans 224 90 0 0 io_wbs_adr[14]
port 154 nsew signal input
flabel metal2 s 78402 0 78458 800 0 FreeSans 224 90 0 0 io_wbs_adr[15]
port 155 nsew signal input
flabel metal2 s 82542 0 82598 800 0 FreeSans 224 90 0 0 io_wbs_adr[16]
port 156 nsew signal input
flabel metal2 s 86682 0 86738 800 0 FreeSans 224 90 0 0 io_wbs_adr[17]
port 157 nsew signal input
flabel metal2 s 90822 0 90878 800 0 FreeSans 224 90 0 0 io_wbs_adr[18]
port 158 nsew signal input
flabel metal2 s 94962 0 95018 800 0 FreeSans 224 90 0 0 io_wbs_adr[19]
port 159 nsew signal input
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 io_wbs_adr[1]
port 160 nsew signal input
flabel metal2 s 99102 0 99158 800 0 FreeSans 224 90 0 0 io_wbs_adr[20]
port 161 nsew signal input
flabel metal2 s 103242 0 103298 800 0 FreeSans 224 90 0 0 io_wbs_adr[21]
port 162 nsew signal input
flabel metal2 s 107382 0 107438 800 0 FreeSans 224 90 0 0 io_wbs_adr[22]
port 163 nsew signal input
flabel metal2 s 111522 0 111578 800 0 FreeSans 224 90 0 0 io_wbs_adr[23]
port 164 nsew signal input
flabel metal2 s 115662 0 115718 800 0 FreeSans 224 90 0 0 io_wbs_adr[24]
port 165 nsew signal input
flabel metal2 s 119802 0 119858 800 0 FreeSans 224 90 0 0 io_wbs_adr[25]
port 166 nsew signal input
flabel metal2 s 123942 0 123998 800 0 FreeSans 224 90 0 0 io_wbs_adr[26]
port 167 nsew signal input
flabel metal2 s 128082 0 128138 800 0 FreeSans 224 90 0 0 io_wbs_adr[27]
port 168 nsew signal input
flabel metal2 s 132222 0 132278 800 0 FreeSans 224 90 0 0 io_wbs_adr[28]
port 169 nsew signal input
flabel metal2 s 136362 0 136418 800 0 FreeSans 224 90 0 0 io_wbs_adr[29]
port 170 nsew signal input
flabel metal2 s 21822 0 21878 800 0 FreeSans 224 90 0 0 io_wbs_adr[2]
port 171 nsew signal input
flabel metal2 s 140502 0 140558 800 0 FreeSans 224 90 0 0 io_wbs_adr[30]
port 172 nsew signal input
flabel metal2 s 144642 0 144698 800 0 FreeSans 224 90 0 0 io_wbs_adr[31]
port 173 nsew signal input
flabel metal2 s 27342 0 27398 800 0 FreeSans 224 90 0 0 io_wbs_adr[3]
port 174 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 io_wbs_adr[4]
port 175 nsew signal input
flabel metal2 s 37002 0 37058 800 0 FreeSans 224 90 0 0 io_wbs_adr[5]
port 176 nsew signal input
flabel metal2 s 41142 0 41198 800 0 FreeSans 224 90 0 0 io_wbs_adr[6]
port 177 nsew signal input
flabel metal2 s 45282 0 45338 800 0 FreeSans 224 90 0 0 io_wbs_adr[7]
port 178 nsew signal input
flabel metal2 s 49422 0 49478 800 0 FreeSans 224 90 0 0 io_wbs_adr[8]
port 179 nsew signal input
flabel metal2 s 53562 0 53618 800 0 FreeSans 224 90 0 0 io_wbs_adr[9]
port 180 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 io_wbs_clk
port 181 nsew signal input
flabel metal2 s 5262 0 5318 800 0 FreeSans 224 90 0 0 io_wbs_cyc
port 182 nsew signal input
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 io_wbs_datrd[0]
port 183 nsew signal tristate
flabel metal2 s 59082 0 59138 800 0 FreeSans 224 90 0 0 io_wbs_datrd[10]
port 184 nsew signal tristate
flabel metal2 s 63222 0 63278 800 0 FreeSans 224 90 0 0 io_wbs_datrd[11]
port 185 nsew signal tristate
flabel metal2 s 67362 0 67418 800 0 FreeSans 224 90 0 0 io_wbs_datrd[12]
port 186 nsew signal tristate
flabel metal2 s 71502 0 71558 800 0 FreeSans 224 90 0 0 io_wbs_datrd[13]
port 187 nsew signal tristate
flabel metal2 s 75642 0 75698 800 0 FreeSans 224 90 0 0 io_wbs_datrd[14]
port 188 nsew signal tristate
flabel metal2 s 79782 0 79838 800 0 FreeSans 224 90 0 0 io_wbs_datrd[15]
port 189 nsew signal tristate
flabel metal2 s 83922 0 83978 800 0 FreeSans 224 90 0 0 io_wbs_datrd[16]
port 190 nsew signal tristate
flabel metal2 s 88062 0 88118 800 0 FreeSans 224 90 0 0 io_wbs_datrd[17]
port 191 nsew signal tristate
flabel metal2 s 92202 0 92258 800 0 FreeSans 224 90 0 0 io_wbs_datrd[18]
port 192 nsew signal tristate
flabel metal2 s 96342 0 96398 800 0 FreeSans 224 90 0 0 io_wbs_datrd[19]
port 193 nsew signal tristate
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 io_wbs_datrd[1]
port 194 nsew signal tristate
flabel metal2 s 100482 0 100538 800 0 FreeSans 224 90 0 0 io_wbs_datrd[20]
port 195 nsew signal tristate
flabel metal2 s 104622 0 104678 800 0 FreeSans 224 90 0 0 io_wbs_datrd[21]
port 196 nsew signal tristate
flabel metal2 s 108762 0 108818 800 0 FreeSans 224 90 0 0 io_wbs_datrd[22]
port 197 nsew signal tristate
flabel metal2 s 112902 0 112958 800 0 FreeSans 224 90 0 0 io_wbs_datrd[23]
port 198 nsew signal tristate
flabel metal2 s 117042 0 117098 800 0 FreeSans 224 90 0 0 io_wbs_datrd[24]
port 199 nsew signal tristate
flabel metal2 s 121182 0 121238 800 0 FreeSans 224 90 0 0 io_wbs_datrd[25]
port 200 nsew signal tristate
flabel metal2 s 125322 0 125378 800 0 FreeSans 224 90 0 0 io_wbs_datrd[26]
port 201 nsew signal tristate
flabel metal2 s 129462 0 129518 800 0 FreeSans 224 90 0 0 io_wbs_datrd[27]
port 202 nsew signal tristate
flabel metal2 s 133602 0 133658 800 0 FreeSans 224 90 0 0 io_wbs_datrd[28]
port 203 nsew signal tristate
flabel metal2 s 137742 0 137798 800 0 FreeSans 224 90 0 0 io_wbs_datrd[29]
port 204 nsew signal tristate
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 io_wbs_datrd[2]
port 205 nsew signal tristate
flabel metal2 s 141882 0 141938 800 0 FreeSans 224 90 0 0 io_wbs_datrd[30]
port 206 nsew signal tristate
flabel metal2 s 146022 0 146078 800 0 FreeSans 224 90 0 0 io_wbs_datrd[31]
port 207 nsew signal tristate
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 io_wbs_datrd[3]
port 208 nsew signal tristate
flabel metal2 s 34242 0 34298 800 0 FreeSans 224 90 0 0 io_wbs_datrd[4]
port 209 nsew signal tristate
flabel metal2 s 38382 0 38438 800 0 FreeSans 224 90 0 0 io_wbs_datrd[5]
port 210 nsew signal tristate
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 io_wbs_datrd[6]
port 211 nsew signal tristate
flabel metal2 s 46662 0 46718 800 0 FreeSans 224 90 0 0 io_wbs_datrd[7]
port 212 nsew signal tristate
flabel metal2 s 50802 0 50858 800 0 FreeSans 224 90 0 0 io_wbs_datrd[8]
port 213 nsew signal tristate
flabel metal2 s 54942 0 54998 800 0 FreeSans 224 90 0 0 io_wbs_datrd[9]
port 214 nsew signal tristate
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 io_wbs_datwr[0]
port 215 nsew signal input
flabel metal2 s 60462 0 60518 800 0 FreeSans 224 90 0 0 io_wbs_datwr[10]
port 216 nsew signal input
flabel metal2 s 64602 0 64658 800 0 FreeSans 224 90 0 0 io_wbs_datwr[11]
port 217 nsew signal input
flabel metal2 s 68742 0 68798 800 0 FreeSans 224 90 0 0 io_wbs_datwr[12]
port 218 nsew signal input
flabel metal2 s 72882 0 72938 800 0 FreeSans 224 90 0 0 io_wbs_datwr[13]
port 219 nsew signal input
flabel metal2 s 77022 0 77078 800 0 FreeSans 224 90 0 0 io_wbs_datwr[14]
port 220 nsew signal input
flabel metal2 s 81162 0 81218 800 0 FreeSans 224 90 0 0 io_wbs_datwr[15]
port 221 nsew signal input
flabel metal2 s 85302 0 85358 800 0 FreeSans 224 90 0 0 io_wbs_datwr[16]
port 222 nsew signal input
flabel metal2 s 89442 0 89498 800 0 FreeSans 224 90 0 0 io_wbs_datwr[17]
port 223 nsew signal input
flabel metal2 s 93582 0 93638 800 0 FreeSans 224 90 0 0 io_wbs_datwr[18]
port 224 nsew signal input
flabel metal2 s 97722 0 97778 800 0 FreeSans 224 90 0 0 io_wbs_datwr[19]
port 225 nsew signal input
flabel metal2 s 19062 0 19118 800 0 FreeSans 224 90 0 0 io_wbs_datwr[1]
port 226 nsew signal input
flabel metal2 s 101862 0 101918 800 0 FreeSans 224 90 0 0 io_wbs_datwr[20]
port 227 nsew signal input
flabel metal2 s 106002 0 106058 800 0 FreeSans 224 90 0 0 io_wbs_datwr[21]
port 228 nsew signal input
flabel metal2 s 110142 0 110198 800 0 FreeSans 224 90 0 0 io_wbs_datwr[22]
port 229 nsew signal input
flabel metal2 s 114282 0 114338 800 0 FreeSans 224 90 0 0 io_wbs_datwr[23]
port 230 nsew signal input
flabel metal2 s 118422 0 118478 800 0 FreeSans 224 90 0 0 io_wbs_datwr[24]
port 231 nsew signal input
flabel metal2 s 122562 0 122618 800 0 FreeSans 224 90 0 0 io_wbs_datwr[25]
port 232 nsew signal input
flabel metal2 s 126702 0 126758 800 0 FreeSans 224 90 0 0 io_wbs_datwr[26]
port 233 nsew signal input
flabel metal2 s 130842 0 130898 800 0 FreeSans 224 90 0 0 io_wbs_datwr[27]
port 234 nsew signal input
flabel metal2 s 134982 0 135038 800 0 FreeSans 224 90 0 0 io_wbs_datwr[28]
port 235 nsew signal input
flabel metal2 s 139122 0 139178 800 0 FreeSans 224 90 0 0 io_wbs_datwr[29]
port 236 nsew signal input
flabel metal2 s 24582 0 24638 800 0 FreeSans 224 90 0 0 io_wbs_datwr[2]
port 237 nsew signal input
flabel metal2 s 143262 0 143318 800 0 FreeSans 224 90 0 0 io_wbs_datwr[30]
port 238 nsew signal input
flabel metal2 s 147402 0 147458 800 0 FreeSans 224 90 0 0 io_wbs_datwr[31]
port 239 nsew signal input
flabel metal2 s 30102 0 30158 800 0 FreeSans 224 90 0 0 io_wbs_datwr[3]
port 240 nsew signal input
flabel metal2 s 35622 0 35678 800 0 FreeSans 224 90 0 0 io_wbs_datwr[4]
port 241 nsew signal input
flabel metal2 s 39762 0 39818 800 0 FreeSans 224 90 0 0 io_wbs_datwr[5]
port 242 nsew signal input
flabel metal2 s 43902 0 43958 800 0 FreeSans 224 90 0 0 io_wbs_datwr[6]
port 243 nsew signal input
flabel metal2 s 48042 0 48098 800 0 FreeSans 224 90 0 0 io_wbs_datwr[7]
port 244 nsew signal input
flabel metal2 s 52182 0 52238 800 0 FreeSans 224 90 0 0 io_wbs_datwr[8]
port 245 nsew signal input
flabel metal2 s 56322 0 56378 800 0 FreeSans 224 90 0 0 io_wbs_datwr[9]
port 246 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 io_wbs_rst
port 247 nsew signal input
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 io_wbs_sel[0]
port 248 nsew signal input
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 io_wbs_sel[1]
port 249 nsew signal input
flabel metal2 s 25962 0 26018 800 0 FreeSans 224 90 0 0 io_wbs_sel[2]
port 250 nsew signal input
flabel metal2 s 31482 0 31538 800 0 FreeSans 224 90 0 0 io_wbs_sel[3]
port 251 nsew signal input
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 io_wbs_stb
port 252 nsew signal input
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 io_wbs_we
port 253 nsew signal input
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 254 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 254 nsew power bidirectional
flabel metal4 s 65648 2128 65968 37584 0 FreeSans 1920 90 0 0 vccd1
port 254 nsew power bidirectional
flabel metal4 s 96368 2128 96688 37584 0 FreeSans 1920 90 0 0 vccd1
port 254 nsew power bidirectional
flabel metal4 s 127088 2128 127408 37584 0 FreeSans 1920 90 0 0 vccd1
port 254 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 255 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 37584 0 FreeSans 1920 90 0 0 vssd1
port 255 nsew ground bidirectional
flabel metal4 s 81008 2128 81328 37584 0 FreeSans 1920 90 0 0 vssd1
port 255 nsew ground bidirectional
flabel metal4 s 111728 2128 112048 37584 0 FreeSans 1920 90 0 0 vssd1
port 255 nsew ground bidirectional
flabel metal4 s 142448 2128 142768 37584 0 FreeSans 1920 90 0 0 vssd1
port 255 nsew ground bidirectional
flabel metal2 s 3606 39200 3662 40000 0 FreeSans 224 90 0 0 web_mem0
port 256 nsew signal tristate
flabel metal2 s 76286 39200 76342 40000 0 FreeSans 224 90 0 0 web_mem1
port 257 nsew signal tristate
flabel metal2 s 7286 39200 7342 40000 0 FreeSans 224 90 0 0 wmask_mem0[0]
port 258 nsew signal tristate
flabel metal2 s 10966 39200 11022 40000 0 FreeSans 224 90 0 0 wmask_mem0[1]
port 259 nsew signal tristate
flabel metal2 s 14646 39200 14702 40000 0 FreeSans 224 90 0 0 wmask_mem0[2]
port 260 nsew signal tristate
flabel metal2 s 18326 39200 18382 40000 0 FreeSans 224 90 0 0 wmask_mem0[3]
port 261 nsew signal tristate
flabel metal2 s 79966 39200 80022 40000 0 FreeSans 224 90 0 0 wmask_mem1[0]
port 262 nsew signal tristate
flabel metal2 s 83646 39200 83702 40000 0 FreeSans 224 90 0 0 wmask_mem1[1]
port 263 nsew signal tristate
flabel metal2 s 87326 39200 87382 40000 0 FreeSans 224 90 0 0 wmask_mem1[2]
port 264 nsew signal tristate
flabel metal2 s 91006 39200 91062 40000 0 FreeSans 224 90 0 0 wmask_mem1[3]
port 265 nsew signal tristate
rlabel metal1 74980 37536 74980 37536 0 vccd1
rlabel metal1 74980 36992 74980 36992 0 vssd1
rlabel metal2 6854 3502 6854 3502 0 _000_
rlabel metal2 9430 3366 9430 3366 0 _001_
rlabel metal1 22494 3366 22494 3366 0 _002_
rlabel metal1 21843 3094 21843 3094 0 _003_
rlabel metal1 27232 2822 27232 2822 0 _004_
rlabel metal1 27646 3543 27646 3543 0 _005_
rlabel metal2 33350 3128 33350 3128 0 _006_
rlabel metal2 35926 3400 35926 3400 0 _007_
rlabel metal1 38548 3910 38548 3910 0 _008_
rlabel metal2 39974 3502 39974 3502 0 _009_
rlabel metal1 44719 2346 44719 2346 0 _010_
rlabel metal1 42780 4454 42780 4454 0 _011_
rlabel metal1 49687 2346 49687 2346 0 _012_
rlabel metal2 46230 3128 46230 3128 0 _013_
rlabel metal1 52217 2346 52217 2346 0 _014_
rlabel metal2 51658 3774 51658 3774 0 _015_
rlabel metal1 63204 3978 63204 3978 0 _016_
rlabel metal2 62330 3434 62330 3434 0 _017_
rlabel metal1 61325 3094 61325 3094 0 _018_
rlabel metal1 58788 3978 58788 3978 0 _019_
rlabel metal2 55246 3502 55246 3502 0 _020_
rlabel metal2 56718 2584 56718 2584 0 _021_
rlabel metal1 66516 3910 66516 3910 0 _022_
rlabel metal2 67298 3230 67298 3230 0 _023_
rlabel metal1 69138 3162 69138 3162 0 _024_
rlabel metal1 70695 3094 70695 3094 0 _025_
rlabel metal2 70978 2074 70978 2074 0 _026_
rlabel metal2 79442 4216 79442 4216 0 _027_
rlabel metal1 82945 2346 82945 2346 0 _028_
rlabel metal2 81374 4318 81374 4318 0 _029_
rlabel metal1 80461 2414 80461 2414 0 _030_
rlabel metal1 83513 2414 83513 2414 0 _031_
rlabel metal1 76038 2890 76038 2890 0 _032_
rlabel metal1 74382 3502 74382 3502 0 _033_
rlabel metal1 5481 2346 5481 2346 0 _034_
rlabel metal1 30820 3366 30820 3366 0 _035_
rlabel metal2 7958 2890 7958 2890 0 _036_
rlabel metal2 22310 3128 22310 3128 0 _037_
rlabel metal2 21666 3264 21666 3264 0 _038_
rlabel metal1 26450 2414 26450 2414 0 _039_
rlabel metal1 26864 3570 26864 3570 0 _040_
rlabel metal1 32614 2312 32614 2312 0 _041_
rlabel metal1 34960 2346 34960 2346 0 _042_
rlabel metal2 37766 3128 37766 3128 0 _043_
rlabel metal2 39238 3502 39238 3502 0 _044_
rlabel metal1 42872 3910 42872 3910 0 _045_
rlabel metal2 41906 3740 41906 3740 0 _046_
rlabel metal1 47886 2346 47886 2346 0 _047_
rlabel metal1 46046 2482 46046 2482 0 _048_
rlabel metal1 51244 2482 51244 2482 0 _049_
rlabel metal2 50922 3502 50922 3502 0 _050_
rlabel metal1 63112 3366 63112 3366 0 _051_
rlabel metal1 61548 3366 61548 3366 0 _052_
rlabel metal2 60030 3230 60030 3230 0 _053_
rlabel metal2 58374 3400 58374 3400 0 _054_
rlabel metal2 54602 3230 54602 3230 0 _055_
rlabel metal1 55982 2312 55982 2312 0 _056_
rlabel metal1 65688 2346 65688 2346 0 _057_
rlabel metal2 65550 3502 65550 3502 0 _058_
rlabel metal1 69598 4046 69598 4046 0 _059_
rlabel metal2 70426 3774 70426 3774 0 _060_
rlabel metal1 71208 2346 71208 2346 0 _061_
rlabel metal2 78798 3740 78798 3740 0 _062_
rlabel metal1 81604 2346 81604 2346 0 _063_
rlabel metal1 79488 4182 79488 4182 0 _064_
rlabel metal1 79626 2482 79626 2482 0 _065_
rlabel metal2 80270 3978 80270 3978 0 _066_
rlabel metal1 76544 3366 76544 3366 0 _067_
rlabel metal1 74060 2822 74060 2822 0 _068_
rlabel metal1 79764 37298 79764 37298 0 _069_
rlabel metal2 75762 4828 75762 4828 0 _070_
rlabel metal1 65826 4250 65826 4250 0 _071_
rlabel metal2 74474 3196 74474 3196 0 _072_
rlabel metal2 78246 5236 78246 5236 0 _073_
rlabel metal1 77096 3502 77096 3502 0 _074_
rlabel metal2 82248 31740 82248 31740 0 _075_
rlabel metal2 81742 4148 81742 4148 0 _076_
rlabel metal1 82938 34102 82938 34102 0 _077_
rlabel metal1 82294 3706 82294 3706 0 _078_
rlabel metal2 83122 5814 83122 5814 0 _079_
rlabel metal2 81466 4658 81466 4658 0 _080_
rlabel metal2 81788 16560 81788 16560 0 _081_
rlabel metal1 80868 3706 80868 3706 0 _082_
rlabel metal2 79810 34153 79810 34153 0 _083_
rlabel metal1 78384 4114 78384 4114 0 _084_
rlabel metal1 71622 4114 71622 4114 0 _085_
rlabel via1 69966 3349 69966 3349 0 _086_
rlabel metal2 66286 37264 66286 37264 0 _087_
rlabel metal2 69092 34612 69092 34612 0 _088_
rlabel metal1 69966 3706 69966 3706 0 _089_
rlabel via1 66843 37094 66843 37094 0 _090_
rlabel metal2 68862 3910 68862 3910 0 _091_
rlabel metal2 66056 31740 66056 31740 0 _092_
rlabel metal1 56534 3536 56534 3536 0 _093_
rlabel metal1 65412 4114 65412 4114 0 _094_
rlabel metal2 65642 36652 65642 36652 0 _095_
rlabel metal1 65182 3706 65182 3706 0 _096_
rlabel metal1 58328 4794 58328 4794 0 _097_
rlabel metal2 57454 3910 57454 3910 0 _098_
rlabel metal1 56166 3570 56166 3570 0 _099_
rlabel metal1 54970 3434 54970 3434 0 _100_
rlabel metal1 58788 3094 58788 3094 0 _101_
rlabel metal1 58144 2890 58144 2890 0 _102_
rlabel metal1 60996 37366 60996 37366 0 _103_
rlabel metal1 60398 3502 60398 3502 0 _104_
rlabel metal1 64032 37094 64032 37094 0 _105_
rlabel metal1 62652 2890 62652 2890 0 _106_
rlabel metal1 63710 36550 63710 36550 0 _107_
rlabel metal1 62468 3502 62468 3502 0 _108_
rlabel metal1 43194 36720 43194 36720 0 _109_
rlabel metal1 52946 5338 52946 5338 0 _110_
rlabel metal1 51658 3706 51658 3706 0 _111_
rlabel metal1 53636 3094 53636 3094 0 _112_
rlabel metal1 52578 2890 52578 2890 0 _113_
rlabel metal1 49036 36618 49036 36618 0 _114_
rlabel metal1 41308 4454 41308 4454 0 _115_
rlabel metal2 47058 4284 47058 4284 0 _116_
rlabel metal1 48806 37094 48806 37094 0 _117_
rlabel metal1 46506 3502 46506 3502 0 _118_
rlabel metal1 41446 2618 41446 2618 0 _119_
rlabel metal1 42136 2822 42136 2822 0 _120_
rlabel metal1 43521 37094 43521 37094 0 _121_
rlabel metal2 43838 3910 43838 3910 0 _122_
rlabel metal1 40572 2346 40572 2346 0 _123_
rlabel metal2 40066 3366 40066 3366 0 _124_
rlabel metal1 38272 5338 38272 5338 0 _125_
rlabel metal2 37490 3638 37490 3638 0 _126_
rlabel metal2 36110 4386 36110 4386 0 _127_
rlabel metal1 34178 3468 34178 3468 0 _128_
rlabel metal1 34362 3162 34362 3162 0 _129_
rlabel metal2 33810 3638 33810 3638 0 _130_
rlabel metal1 28106 3094 28106 3094 0 _131_
rlabel metal2 27370 3638 27370 3638 0 _132_
rlabel metal1 28750 36754 28750 36754 0 _133_
rlabel metal1 25806 2992 25806 2992 0 _134_
rlabel metal1 24380 36550 24380 36550 0 _135_
rlabel metal1 21482 3468 21482 3468 0 _136_
rlabel metal1 24371 37094 24371 37094 0 _137_
rlabel metal2 22770 3910 22770 3910 0 _138_
rlabel metal2 6026 3604 6026 3604 0 _139_
rlabel metal2 76130 36346 76130 36346 0 _140_
rlabel metal1 60375 37162 60375 37162 0 _141_
rlabel metal2 6302 3706 6302 3706 0 _142_
rlabel metal1 38134 4114 38134 4114 0 _143_
rlabel metal1 56580 3026 56580 3026 0 _144_
rlabel metal1 79074 5202 79074 5202 0 _145_
rlabel metal1 4692 37094 4692 37094 0 addr_mem0[0]
rlabel metal1 8372 37094 8372 37094 0 addr_mem0[1]
rlabel metal1 12006 37094 12006 37094 0 addr_mem0[2]
rlabel metal1 15686 37094 15686 37094 0 addr_mem0[3]
rlabel metal1 19458 37094 19458 37094 0 addr_mem0[4]
rlabel metal1 22172 37094 22172 37094 0 addr_mem0[5]
rlabel metal1 24932 36346 24932 36346 0 addr_mem0[6]
rlabel metal1 27692 36346 27692 36346 0 addr_mem0[7]
rlabel metal1 30452 36890 30452 36890 0 addr_mem0[8]
rlabel metal1 77556 37094 77556 37094 0 addr_mem1[0]
rlabel metal1 81052 35802 81052 35802 0 addr_mem1[1]
rlabel metal1 85514 37128 85514 37128 0 addr_mem1[2]
rlabel metal1 88734 37094 88734 37094 0 addr_mem1[3]
rlabel metal1 92230 37094 92230 37094 0 addr_mem1[4]
rlabel metal1 95496 37094 95496 37094 0 addr_mem1[5]
rlabel metal1 98164 37094 98164 37094 0 addr_mem1[6]
rlabel metal1 100878 37094 100878 37094 0 addr_mem1[7]
rlabel metal1 103132 36550 103132 36550 0 addr_mem1[8]
rlabel metal2 38226 3264 38226 3264 0 clknet_0_io_wbs_clk
rlabel metal1 38686 4454 38686 4454 0 clknet_2_0__leaf_io_wbs_clk
rlabel metal1 6486 2482 6486 2482 0 clknet_2_1__leaf_io_wbs_clk
rlabel metal1 60950 2550 60950 2550 0 clknet_2_2__leaf_io_wbs_clk
rlabel metal1 59754 3094 59754 3094 0 clknet_2_3__leaf_io_wbs_clk
rlabel metal1 5612 37094 5612 37094 0 din_mem0[0]
rlabel metal1 34316 37094 34316 37094 0 din_mem0[10]
rlabel metal2 36754 38056 36754 38056 0 din_mem0[11]
rlabel metal1 38962 37094 38962 37094 0 din_mem0[12]
rlabel metal1 40342 37094 40342 37094 0 din_mem0[13]
rlabel metal1 42366 36346 42366 36346 0 din_mem0[14]
rlabel metal1 44022 36890 44022 36890 0 din_mem0[15]
rlabel metal1 46046 36618 46046 36618 0 din_mem0[16]
rlabel metal1 47472 37094 47472 37094 0 din_mem0[17]
rlabel metal2 49634 38158 49634 38158 0 din_mem0[18]
rlabel metal2 51474 38158 51474 38158 0 din_mem0[19]
rlabel metal1 9246 37094 9246 37094 0 din_mem0[1]
rlabel metal1 53452 36346 53452 36346 0 din_mem0[20]
rlabel metal1 54970 37094 54970 37094 0 din_mem0[21]
rlabel metal1 56396 37094 56396 37094 0 din_mem0[22]
rlabel metal1 59248 36346 59248 36346 0 din_mem0[23]
rlabel metal1 60490 36890 60490 36890 0 din_mem0[24]
rlabel metal1 62606 36346 62606 36346 0 din_mem0[25]
rlabel metal1 64446 36346 64446 36346 0 din_mem0[26]
rlabel metal1 66332 36890 66332 36890 0 din_mem0[27]
rlabel metal1 68126 36346 68126 36346 0 din_mem0[28]
rlabel metal1 69966 37094 69966 37094 0 din_mem0[29]
rlabel metal1 12926 37094 12926 37094 0 din_mem0[2]
rlabel metal1 72036 37094 72036 37094 0 din_mem0[30]
rlabel metal1 74014 37094 74014 37094 0 din_mem0[31]
rlabel metal1 16790 37094 16790 37094 0 din_mem0[3]
rlabel metal1 20286 37094 20286 37094 0 din_mem0[4]
rlabel metal1 23046 37094 23046 37094 0 din_mem0[5]
rlabel metal1 25806 36346 25806 36346 0 din_mem0[6]
rlabel metal1 28704 36890 28704 36890 0 din_mem0[7]
rlabel metal1 31326 37094 31326 37094 0 din_mem0[8]
rlabel metal1 33212 36890 33212 36890 0 din_mem0[9]
rlabel metal1 78752 36890 78752 36890 0 din_mem1[0]
rlabel metal1 107824 37094 107824 37094 0 din_mem1[10]
rlabel metal1 109618 37094 109618 37094 0 din_mem1[11]
rlabel metal1 112102 37094 112102 37094 0 din_mem1[12]
rlabel metal1 113528 37094 113528 37094 0 din_mem1[13]
rlabel metal1 115368 37094 115368 37094 0 din_mem1[14]
rlabel metal1 117438 37094 117438 37094 0 din_mem1[15]
rlabel metal2 118634 38158 118634 38158 0 din_mem1[16]
rlabel metal1 120980 37434 120980 37434 0 din_mem1[17]
rlabel metal1 123142 37094 123142 37094 0 din_mem1[18]
rlabel metal1 124752 37094 124752 37094 0 din_mem1[19]
rlabel metal1 82616 36550 82616 36550 0 din_mem1[1]
rlabel metal1 126408 37094 126408 37094 0 din_mem1[20]
rlabel metal1 128478 37094 128478 37094 0 din_mem1[21]
rlabel metal1 130088 37094 130088 37094 0 din_mem1[22]
rlabel metal1 131698 37094 131698 37094 0 din_mem1[23]
rlabel metal1 133538 37094 133538 37094 0 din_mem1[24]
rlabel metal2 135194 37551 135194 37551 0 din_mem1[25]
rlabel metal1 137172 37094 137172 37094 0 din_mem1[26]
rlabel metal1 139012 37094 139012 37094 0 din_mem1[27]
rlabel metal1 141128 37094 141128 37094 0 din_mem1[28]
rlabel metal1 142922 37094 142922 37094 0 din_mem1[29]
rlabel metal1 86066 37094 86066 37094 0 din_mem1[2]
rlabel metal1 144578 37094 144578 37094 0 din_mem1[30]
rlabel metal1 146418 37094 146418 37094 0 din_mem1[31]
rlabel metal1 89332 36550 89332 36550 0 din_mem1[3]
rlabel metal1 93058 37094 93058 37094 0 din_mem1[4]
rlabel metal1 95726 36550 95726 36550 0 din_mem1[5]
rlabel metal2 98670 37893 98670 37893 0 din_mem1[6]
rlabel metal1 101292 36550 101292 36550 0 din_mem1[7]
rlabel metal1 104282 37094 104282 37094 0 din_mem1[8]
rlabel metal1 105984 36550 105984 36550 0 din_mem1[9]
rlabel metal1 6486 36754 6486 36754 0 dout_mem0[0]
rlabel metal2 35834 37376 35834 37376 0 dout_mem0[10]
rlabel metal1 37720 36142 37720 36142 0 dout_mem0[11]
rlabel metal2 39514 37784 39514 37784 0 dout_mem0[12]
rlabel metal2 41170 36669 41170 36669 0 dout_mem0[13]
rlabel metal1 44068 35802 44068 35802 0 dout_mem0[14]
rlabel metal1 45172 36754 45172 36754 0 dout_mem0[15]
rlabel metal1 46920 36142 46920 36142 0 dout_mem0[16]
rlabel metal1 49036 36142 49036 36142 0 dout_mem0[17]
rlabel metal2 50600 37196 50600 37196 0 dout_mem0[18]
rlabel metal2 52302 36499 52302 36499 0 dout_mem0[19]
rlabel metal1 10120 37230 10120 37230 0 dout_mem0[1]
rlabel metal1 54970 36720 54970 36720 0 dout_mem0[20]
rlabel metal1 56212 36754 56212 36754 0 dout_mem0[21]
rlabel metal2 58006 36414 58006 36414 0 dout_mem0[22]
rlabel metal1 60628 36142 60628 36142 0 dout_mem0[23]
rlabel metal1 62330 36754 62330 36754 0 dout_mem0[24]
rlabel metal1 63342 36754 63342 36754 0 dout_mem0[25]
rlabel metal1 65320 35666 65320 35666 0 dout_mem0[26]
rlabel metal1 67160 36754 67160 36754 0 dout_mem0[27]
rlabel metal1 69000 36142 69000 36142 0 dout_mem0[28]
rlabel metal1 70840 36754 70840 36754 0 dout_mem0[29]
rlabel metal2 13846 36822 13846 36822 0 dout_mem0[2]
rlabel metal1 72680 36754 72680 36754 0 dout_mem0[30]
rlabel metal1 74520 36142 74520 36142 0 dout_mem0[31]
rlabel metal1 17526 37230 17526 37230 0 dout_mem0[3]
rlabel metal1 21160 36142 21160 36142 0 dout_mem0[4]
rlabel metal1 23598 36754 23598 36754 0 dout_mem0[5]
rlabel metal1 26680 36142 26680 36142 0 dout_mem0[6]
rlabel metal1 29026 37196 29026 37196 0 dout_mem0[7]
rlabel metal1 32200 36142 32200 36142 0 dout_mem0[8]
rlabel metal1 34040 36754 34040 36754 0 dout_mem0[9]
rlabel metal2 80454 37349 80454 37349 0 dout_mem1[0]
rlabel metal1 108560 37230 108560 37230 0 dout_mem1[10]
rlabel metal1 110906 37230 110906 37230 0 dout_mem1[11]
rlabel metal1 112608 37230 112608 37230 0 dout_mem1[12]
rlabel metal1 114402 37230 114402 37230 0 dout_mem1[13]
rlabel metal1 116196 37230 116196 37230 0 dout_mem1[14]
rlabel metal1 117990 37162 117990 37162 0 dout_mem1[15]
rlabel metal1 119738 37230 119738 37230 0 dout_mem1[16]
rlabel metal1 121440 36754 121440 36754 0 dout_mem1[17]
rlabel metal1 123786 37230 123786 37230 0 dout_mem1[18]
rlabel metal1 125488 37230 125488 37230 0 dout_mem1[19]
rlabel metal1 83904 37230 83904 37230 0 dout_mem1[1]
rlabel metal1 127328 37230 127328 37230 0 dout_mem1[20]
rlabel metal1 128938 37230 128938 37230 0 dout_mem1[21]
rlabel metal1 131192 37230 131192 37230 0 dout_mem1[22]
rlabel metal1 132802 37230 132802 37230 0 dout_mem1[23]
rlabel metal1 134320 37230 134320 37230 0 dout_mem1[24]
rlabel metal1 136252 37162 136252 37162 0 dout_mem1[25]
rlabel metal1 138138 37230 138138 37230 0 dout_mem1[26]
rlabel metal1 140162 37230 140162 37230 0 dout_mem1[27]
rlabel metal2 141634 38226 141634 38226 0 dout_mem1[28]
rlabel metal1 143704 37230 143704 37230 0 dout_mem1[29]
rlabel metal1 87216 37230 87216 37230 0 dout_mem1[2]
rlabel metal1 145498 37230 145498 37230 0 dout_mem1[30]
rlabel metal1 147200 37230 147200 37230 0 dout_mem1[31]
rlabel metal1 90436 37230 90436 37230 0 dout_mem1[3]
rlabel metal1 94116 37230 94116 37230 0 dout_mem1[4]
rlabel metal1 96876 37230 96876 37230 0 dout_mem1[5]
rlabel metal2 99866 37026 99866 37026 0 dout_mem1[6]
rlabel metal1 102902 37264 102902 37264 0 dout_mem1[7]
rlabel metal1 105064 37230 105064 37230 0 dout_mem1[8]
rlabel metal1 106996 37230 106996 37230 0 dout_mem1[9]
rlabel metal2 2530 1520 2530 1520 0 io_wbs_ack
rlabel metal1 57776 3094 57776 3094 0 io_wbs_adr[10]
rlabel metal1 61916 3026 61916 3026 0 io_wbs_adr[11]
rlabel metal1 21666 2414 21666 2414 0 io_wbs_adr[2]
rlabel metal1 26450 2312 26450 2312 0 io_wbs_adr[3]
rlabel metal1 32982 3434 32982 3434 0 io_wbs_adr[4]
rlabel metal1 37444 4182 37444 4182 0 io_wbs_adr[5]
rlabel metal1 41124 3434 41124 3434 0 io_wbs_adr[6]
rlabel metal2 45356 2244 45356 2244 0 io_wbs_adr[7]
rlabel metal1 49542 4114 49542 4114 0 io_wbs_adr[8]
rlabel metal1 53682 3434 53682 3434 0 io_wbs_adr[9]
rlabel metal2 3910 1860 3910 1860 0 io_wbs_clk
rlabel metal1 5336 3502 5336 3502 0 io_wbs_cyc
rlabel metal2 12190 1520 12190 1520 0 io_wbs_datrd[0]
rlabel metal2 59110 2064 59110 2064 0 io_wbs_datrd[10]
rlabel metal1 63388 3910 63388 3910 0 io_wbs_datrd[11]
rlabel metal1 67574 2822 67574 2822 0 io_wbs_datrd[12]
rlabel metal1 72082 2890 72082 2890 0 io_wbs_datrd[13]
rlabel metal1 75808 2822 75808 2822 0 io_wbs_datrd[14]
rlabel metal1 78936 3162 78936 3162 0 io_wbs_datrd[15]
rlabel metal2 83950 1520 83950 1520 0 io_wbs_datrd[16]
rlabel metal2 88090 1520 88090 1520 0 io_wbs_datrd[17]
rlabel metal2 92230 1520 92230 1520 0 io_wbs_datrd[18]
rlabel metal2 96370 1520 96370 1520 0 io_wbs_datrd[19]
rlabel metal2 17710 1520 17710 1520 0 io_wbs_datrd[1]
rlabel metal2 100510 1520 100510 1520 0 io_wbs_datrd[20]
rlabel metal2 104650 1520 104650 1520 0 io_wbs_datrd[21]
rlabel metal2 108790 1656 108790 1656 0 io_wbs_datrd[22]
rlabel metal2 112930 1520 112930 1520 0 io_wbs_datrd[23]
rlabel metal2 117070 1520 117070 1520 0 io_wbs_datrd[24]
rlabel metal2 121210 1520 121210 1520 0 io_wbs_datrd[25]
rlabel metal2 125350 1520 125350 1520 0 io_wbs_datrd[26]
rlabel metal2 129490 959 129490 959 0 io_wbs_datrd[27]
rlabel metal2 133630 1520 133630 1520 0 io_wbs_datrd[28]
rlabel metal2 137770 1520 137770 1520 0 io_wbs_datrd[29]
rlabel metal1 23322 3910 23322 3910 0 io_wbs_datrd[2]
rlabel metal2 141910 1520 141910 1520 0 io_wbs_datrd[30]
rlabel metal2 146050 1520 146050 1520 0 io_wbs_datrd[31]
rlabel metal1 28888 3638 28888 3638 0 io_wbs_datrd[3]
rlabel metal2 34270 2336 34270 2336 0 io_wbs_datrd[4]
rlabel metal2 38410 2064 38410 2064 0 io_wbs_datrd[5]
rlabel metal2 42550 1520 42550 1520 0 io_wbs_datrd[6]
rlabel metal1 46828 2822 46828 2822 0 io_wbs_datrd[7]
rlabel metal2 50830 2064 50830 2064 0 io_wbs_datrd[8]
rlabel metal2 54970 1656 54970 1656 0 io_wbs_datrd[9]
rlabel metal1 13616 2278 13616 2278 0 io_wbs_datwr[0]
rlabel metal1 60582 4114 60582 4114 0 io_wbs_datwr[10]
rlabel metal1 64492 3094 64492 3094 0 io_wbs_datwr[11]
rlabel metal2 68770 1554 68770 1554 0 io_wbs_datwr[12]
rlabel metal1 72956 3366 72956 3366 0 io_wbs_datwr[13]
rlabel metal1 77188 3026 77188 3026 0 io_wbs_datwr[14]
rlabel metal1 83214 3026 83214 3026 0 io_wbs_datwr[15]
rlabel metal1 85468 2346 85468 2346 0 io_wbs_datwr[16]
rlabel metal1 89562 2346 89562 2346 0 io_wbs_datwr[17]
rlabel metal1 94047 2346 94047 2346 0 io_wbs_datwr[18]
rlabel metal1 97842 2346 97842 2346 0 io_wbs_datwr[19]
rlabel metal1 18998 2278 18998 2278 0 io_wbs_datwr[1]
rlabel metal1 101982 2346 101982 2346 0 io_wbs_datwr[20]
rlabel metal1 106122 2346 106122 2346 0 io_wbs_datwr[21]
rlabel metal2 110446 2023 110446 2023 0 io_wbs_datwr[22]
rlabel metal1 114264 2278 114264 2278 0 io_wbs_datwr[23]
rlabel metal1 118542 2346 118542 2346 0 io_wbs_datwr[24]
rlabel metal1 122682 2346 122682 2346 0 io_wbs_datwr[25]
rlabel metal1 126822 2346 126822 2346 0 io_wbs_datwr[26]
rlabel metal1 130962 2346 130962 2346 0 io_wbs_datwr[27]
rlabel metal1 134918 2278 134918 2278 0 io_wbs_datwr[28]
rlabel metal1 139196 2414 139196 2414 0 io_wbs_datwr[29]
rlabel metal2 24886 2159 24886 2159 0 io_wbs_datwr[2]
rlabel metal1 143382 2346 143382 2346 0 io_wbs_datwr[30]
rlabel metal1 147522 2346 147522 2346 0 io_wbs_datwr[31]
rlabel metal1 30544 3094 30544 3094 0 io_wbs_datwr[3]
rlabel metal1 35742 4182 35742 4182 0 io_wbs_datwr[4]
rlabel metal1 39652 3366 39652 3366 0 io_wbs_datwr[5]
rlabel metal1 43838 3910 43838 3910 0 io_wbs_datwr[6]
rlabel metal2 48070 1761 48070 1761 0 io_wbs_datwr[7]
rlabel metal1 52762 4182 52762 4182 0 io_wbs_datwr[8]
rlabel metal1 56442 4182 56442 4182 0 io_wbs_datwr[9]
rlabel metal2 6670 2132 6670 2132 0 io_wbs_rst
rlabel metal1 15088 2414 15088 2414 0 io_wbs_sel[0]
rlabel metal1 20516 2346 20516 2346 0 io_wbs_sel[1]
rlabel metal1 25898 2346 25898 2346 0 io_wbs_sel[2]
rlabel metal2 31510 1761 31510 1761 0 io_wbs_sel[3]
rlabel metal1 8188 3026 8188 3026 0 io_wbs_stb
rlabel metal1 9568 2414 9568 2414 0 io_wbs_we
rlabel metal2 22770 36703 22770 36703 0 net1
rlabel metal1 51060 36278 51060 36278 0 net10
rlabel metal1 146234 36754 146234 36754 0 net100
rlabel metal1 24150 36108 24150 36108 0 net101
rlabel metal2 23966 36992 23966 36992 0 net102
rlabel metal1 40066 35462 40066 35462 0 net103
rlabel metal1 43654 36108 43654 36108 0 net104
rlabel metal2 47242 36482 47242 36482 0 net105
rlabel metal1 53176 4114 53176 4114 0 net106
rlabel metal1 56672 4114 56672 4114 0 net107
rlabel metal2 6762 3196 6762 3196 0 net108
rlabel metal1 9292 36550 9292 36550 0 net109
rlabel metal2 58098 36584 58098 36584 0 net11
rlabel metal1 20194 36074 20194 36074 0 net110
rlabel metal1 25576 37094 25576 37094 0 net111
rlabel metal2 31142 36924 31142 36924 0 net112
rlabel metal1 6992 3162 6992 3162 0 net113
rlabel metal1 9476 2618 9476 2618 0 net114
rlabel metal2 4922 37026 4922 37026 0 net115
rlabel metal2 25162 37468 25162 37468 0 net116
rlabel metal2 12282 37060 12282 37060 0 net117
rlabel metal1 16928 36550 16928 36550 0 net118
rlabel metal3 22172 37264 22172 37264 0 net119
rlabel metal2 10350 36618 10350 36618 0 net12
rlabel metal1 22402 37298 22402 37298 0 net120
rlabel metal1 25208 35802 25208 35802 0 net121
rlabel metal1 29578 35530 29578 35530 0 net122
rlabel metal1 30728 36346 30728 36346 0 net123
rlabel metal2 53774 36193 53774 36193 0 net124
rlabel metal2 30038 36499 30038 36499 0 net125
rlabel metal2 33626 37570 33626 37570 0 net126
rlabel metal2 38870 35428 38870 35428 0 net127
rlabel metal2 41998 35309 41998 35309 0 net128
rlabel metal2 45402 37604 45402 37604 0 net129
rlabel metal2 55154 36414 55154 36414 0 net13
rlabel metal1 50692 36754 50692 36754 0 net130
rlabel metal2 54418 35768 54418 35768 0 net131
rlabel metal1 103040 36346 103040 36346 0 net132
rlabel metal1 6210 37230 6210 37230 0 net133
rlabel metal1 37973 35734 37973 35734 0 net134
rlabel metal2 63710 35564 63710 35564 0 net135
rlabel metal2 39422 38250 39422 38250 0 net136
rlabel metal2 40066 36618 40066 36618 0 net137
rlabel metal2 42642 37740 42642 37740 0 net138
rlabel metal1 44068 36754 44068 36754 0 net139
rlabel metal1 56626 36550 56626 36550 0 net14
rlabel metal2 46322 37978 46322 37978 0 net140
rlabel metal2 46966 38080 46966 38080 0 net141
rlabel metal2 49818 38046 49818 38046 0 net142
rlabel metal2 51198 37604 51198 37604 0 net143
rlabel metal2 9798 37060 9798 37060 0 net144
rlabel metal2 101982 37672 101982 37672 0 net145
rlabel metal1 105340 36822 105340 36822 0 net146
rlabel metal1 56120 37230 56120 37230 0 net147
rlabel metal1 59892 36142 59892 36142 0 net148
rlabel metal2 60122 37672 60122 37672 0 net149
rlabel metal1 61088 36006 61088 36006 0 net15
rlabel metal2 62882 37298 62882 37298 0 net150
rlabel metal2 64722 37230 64722 37230 0 net151
rlabel metal2 130318 37332 130318 37332 0 net152
rlabel metal2 68402 36924 68402 36924 0 net153
rlabel metal2 70518 36482 70518 36482 0 net154
rlabel metal1 23874 37128 23874 37128 0 net155
rlabel metal2 105938 35564 105938 35564 0 net156
rlabel metal1 74658 37162 74658 37162 0 net157
rlabel metal2 17342 37060 17342 37060 0 net158
rlabel metal2 20654 37060 20654 37060 0 net159
rlabel metal1 61732 36278 61732 36278 0 net16
rlabel metal2 23322 37145 23322 37145 0 net160
rlabel metal2 42918 36295 42918 36295 0 net161
rlabel metal2 29118 35734 29118 35734 0 net162
rlabel metal1 31464 37230 31464 37230 0 net163
rlabel metal2 55614 36958 55614 36958 0 net164
rlabel metal2 46230 35462 46230 35462 0 net165
rlabel metal1 107732 36346 107732 36346 0 net166
rlabel metal2 109618 35258 109618 35258 0 net167
rlabel metal2 112194 34952 112194 34952 0 net168
rlabel metal2 75854 35734 75854 35734 0 net169
rlabel metal2 71346 36856 71346 36856 0 net17
rlabel metal1 105754 36176 105754 36176 0 net170
rlabel metal2 99498 36720 99498 36720 0 net171
rlabel metal2 86434 36414 86434 36414 0 net172
rlabel metal2 90482 36040 90482 36040 0 net173
rlabel metal2 95082 38148 95082 38148 0 net174
rlabel metal2 99498 37638 99498 37638 0 net175
rlabel metal2 21390 35292 21390 35292 0 net176
rlabel metal1 126500 37230 126500 37230 0 net177
rlabel metal2 128386 36839 128386 36839 0 net178
rlabel metal2 129582 36703 129582 36703 0 net179
rlabel metal2 79166 37060 79166 37060 0 net18
rlabel metal2 131698 36737 131698 36737 0 net180
rlabel metal2 133538 37026 133538 37026 0 net181
rlabel metal2 134458 36958 134458 36958 0 net182
rlabel metal2 136022 37060 136022 37060 0 net183
rlabel metal1 138414 36890 138414 36890 0 net184
rlabel metal1 141266 37196 141266 37196 0 net185
rlabel metal2 143106 37060 143106 37060 0 net186
rlabel metal2 25990 35054 25990 35054 0 net187
rlabel metal1 144210 36890 144210 36890 0 net188
rlabel metal2 146326 37060 146326 37060 0 net189
rlabel metal2 81466 36346 81466 36346 0 net19
rlabel metal2 31786 35547 31786 35547 0 net190
rlabel metal2 37214 35513 37214 35513 0 net191
rlabel metal2 41354 35071 41354 35071 0 net192
rlabel metal2 44850 34680 44850 34680 0 net193
rlabel metal1 101016 36754 101016 36754 0 net194
rlabel metal2 104466 36890 104466 36890 0 net195
rlabel metal2 106398 36550 106398 36550 0 net196
rlabel metal1 4462 2618 4462 2618 0 net197
rlabel metal1 21712 2278 21712 2278 0 net198
rlabel metal1 55338 4114 55338 4114 0 net199
rlabel metal2 39974 36295 39974 36295 0 net2
rlabel metal2 73002 36890 73002 36890 0 net20
rlabel metal2 48162 4828 48162 4828 0 net200
rlabel metal2 53314 3400 53314 3400 0 net201
rlabel metal2 57730 3570 57730 3570 0 net202
rlabel metal1 65044 2618 65044 2618 0 net203
rlabel metal1 63158 2618 63158 2618 0 net204
rlabel metal2 81374 2448 81374 2448 0 net205
rlabel metal2 59846 1938 59846 1938 0 net206
rlabel metal2 56074 2414 56074 2414 0 net207
rlabel metal2 57454 2176 57454 2176 0 net208
rlabel metal1 21988 2958 21988 2958 0 net209
rlabel metal1 70794 36312 70794 36312 0 net21
rlabel metal2 100050 2108 100050 2108 0 net210
rlabel metal1 79810 3672 79810 3672 0 net211
rlabel metal2 109066 2006 109066 2006 0 net212
rlabel metal1 78982 3978 78982 3978 0 net213
rlabel metal2 116702 2040 116702 2040 0 net214
rlabel metal1 121026 2414 121026 2414 0 net215
rlabel metal2 83030 1904 83030 1904 0 net216
rlabel metal2 117254 3230 117254 3230 0 net217
rlabel metal1 83536 2550 83536 2550 0 net218
rlabel metal2 137310 2856 137310 2856 0 net219
rlabel metal2 71070 36380 71070 36380 0 net22
rlabel metal1 28796 3094 28796 3094 0 net220
rlabel metal1 77924 3366 77924 3366 0 net221
rlabel metal1 76360 3502 76360 3502 0 net222
rlabel metal1 28428 3366 28428 3366 0 net223
rlabel metal2 34178 3638 34178 3638 0 net224
rlabel metal1 36892 2618 36892 2618 0 net225
rlabel metal2 39238 2788 39238 2788 0 net226
rlabel metal1 40572 2414 40572 2414 0 net227
rlabel metal1 44298 2618 44298 2618 0 net228
rlabel metal2 51934 2958 51934 2958 0 net229
rlabel metal1 16054 36618 16054 36618 0 net23
rlabel metal2 4554 37128 4554 37128 0 net230
rlabel metal2 76314 36550 76314 36550 0 net231
rlabel metal2 8234 37060 8234 37060 0 net232
rlabel metal1 11178 37196 11178 37196 0 net233
rlabel metal1 25024 36550 25024 36550 0 net234
rlabel metal2 19090 37060 19090 37060 0 net235
rlabel metal1 44298 35156 44298 35156 0 net236
rlabel metal2 22218 37842 22218 37842 0 net237
rlabel metal2 26542 35020 26542 35020 0 net238
rlabel metal2 32522 34952 32522 34952 0 net239
rlabel metal1 73830 36890 73830 36890 0 net24
rlabel metal2 2806 37859 2806 37859 0 net240
rlabel metal1 75072 36618 75072 36618 0 net241
rlabel metal1 75164 36346 75164 36346 0 net25
rlabel metal1 25898 36720 25898 36720 0 net26
rlabel metal1 24058 36040 24058 36040 0 net27
rlabel metal2 23966 36380 23966 36380 0 net28
rlabel metal1 28474 36040 28474 36040 0 net29
rlabel metal1 39698 36312 39698 36312 0 net3
rlabel metal2 29670 36992 29670 36992 0 net30
rlabel metal2 41538 36652 41538 36652 0 net31
rlabel metal1 42872 36890 42872 36890 0 net32
rlabel metal1 24610 36278 24610 36278 0 net33
rlabel metal2 48162 34170 48162 34170 0 net34
rlabel metal2 48070 37468 48070 37468 0 net35
rlabel metal2 53222 37740 53222 37740 0 net36
rlabel metal2 51566 34510 51566 34510 0 net37
rlabel metal2 116242 37536 116242 37536 0 net38
rlabel metal2 118082 38182 118082 38182 0 net39
rlabel metal2 42090 36278 42090 36278 0 net4
rlabel metal2 120106 37978 120106 37978 0 net40
rlabel metal1 58466 36686 58466 36686 0 net41
rlabel metal1 57408 37094 57408 37094 0 net42
rlabel metal1 125948 37434 125948 37434 0 net43
rlabel metal2 24518 36873 24518 36873 0 net44
rlabel metal1 123234 36584 123234 36584 0 net45
rlabel metal2 129306 36057 129306 36057 0 net46
rlabel metal2 130502 36550 130502 36550 0 net47
rlabel metal2 132894 37145 132894 37145 0 net48
rlabel metal2 134550 36125 134550 36125 0 net49
rlabel metal1 41630 36244 41630 36244 0 net5
rlabel metal1 80224 36890 80224 36890 0 net50
rlabel metal1 138046 37332 138046 37332 0 net51
rlabel metal2 140714 36176 140714 36176 0 net52
rlabel metal1 99498 37128 99498 37128 0 net53
rlabel metal2 144026 35734 144026 35734 0 net54
rlabel metal1 28106 37264 28106 37264 0 net55
rlabel metal2 137310 36550 137310 36550 0 net56
rlabel metal2 147430 35088 147430 35088 0 net57
rlabel metal1 28612 36686 28612 36686 0 net58
rlabel metal2 35558 37978 35558 37978 0 net59
rlabel metal1 63158 34918 63158 34918 0 net6
rlabel metal3 45540 37128 45540 37128 0 net60
rlabel metal2 100234 36873 100234 36873 0 net61
rlabel metal2 102718 36601 102718 36601 0 net62
rlabel metal1 43608 37162 43608 37162 0 net63
rlabel metal2 43102 36737 43102 36737 0 net64
rlabel metal1 57178 35462 57178 35462 0 net65
rlabel metal1 25162 37162 25162 37162 0 net66
rlabel metal1 43562 36040 43562 36040 0 net67
rlabel metal1 26680 36550 26680 36550 0 net68
rlabel metal1 32798 36754 32798 36754 0 net69
rlabel metal1 46138 36550 46138 36550 0 net7
rlabel metal1 37720 4114 37720 4114 0 net70
rlabel metal1 41216 35462 41216 35462 0 net71
rlabel metal1 44574 37264 44574 37264 0 net72
rlabel metal1 49542 36074 49542 36074 0 net73
rlabel metal1 54004 35462 54004 35462 0 net74
rlabel metal2 5750 3264 5750 3264 0 net75
rlabel via2 45310 35989 45310 35989 0 net76
rlabel metal1 60490 35496 60490 35496 0 net77
rlabel metal1 64998 36006 64998 36006 0 net78
rlabel metal2 69230 34986 69230 34986 0 net79
rlabel metal2 58742 36720 58742 36720 0 net8
rlabel metal1 74428 24174 74428 24174 0 net80
rlabel metal1 77878 5542 77878 5542 0 net81
rlabel metal2 83076 26220 83076 26220 0 net82
rlabel metal1 85468 36006 85468 36006 0 net83
rlabel metal1 89976 36006 89976 36006 0 net84
rlabel metal1 94530 36006 94530 36006 0 net85
rlabel metal1 97934 2618 97934 2618 0 net86
rlabel metal1 19872 2550 19872 2550 0 net87
rlabel metal1 102212 36550 102212 36550 0 net88
rlabel metal1 107180 36754 107180 36754 0 net89
rlabel metal1 49542 36244 49542 36244 0 net9
rlabel metal1 110446 36550 110446 36550 0 net90
rlabel metal1 114908 2618 114908 2618 0 net91
rlabel metal2 132066 36516 132066 36516 0 net92
rlabel metal1 122820 36550 122820 36550 0 net93
rlabel metal1 135378 36754 135378 36754 0 net94
rlabel metal2 137678 36380 137678 36380 0 net95
rlabel metal1 137540 2550 137540 2550 0 net96
rlabel metal1 140392 2618 140392 2618 0 net97
rlabel metal1 25806 36788 25806 36788 0 net98
rlabel metal1 107364 36346 107364 36346 0 net99
rlabel metal1 5750 2312 5750 2312 0 operation
rlabel metal2 31786 16014 31786 16014 0 web_mem
rlabel metal1 3726 36890 3726 36890 0 web_mem0
rlabel metal1 76452 36890 76452 36890 0 web_mem1
rlabel metal1 7406 37094 7406 37094 0 wmask_mem0[0]
rlabel metal2 10994 38158 10994 38158 0 wmask_mem0[1]
rlabel metal1 14766 37094 14766 37094 0 wmask_mem0[2]
rlabel metal1 18446 37094 18446 37094 0 wmask_mem0[3]
rlabel metal2 79994 38617 79994 38617 0 wmask_mem1[0]
rlabel metal1 83858 36550 83858 36550 0 wmask_mem1[1]
rlabel metal1 87676 37094 87676 37094 0 wmask_mem1[2]
rlabel metal1 91448 37094 91448 37094 0 wmask_mem1[3]
<< properties >>
string FIXED_BBOX 0 0 150000 40000
<< end >>
