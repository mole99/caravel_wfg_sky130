VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wfg_top
  CLASS BLOCK ;
  FOREIGN wfg_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 750.000 BY 550.000 ;
  PIN addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END addr1[0]
  PIN addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END addr1[1]
  PIN addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END addr1[2]
  PIN addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END addr1[3]
  PIN addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END addr1[4]
  PIN addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END addr1[5]
  PIN addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END addr1[6]
  PIN addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END addr1[7]
  PIN addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END addr1[8]
  PIN addr1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END addr1[9]
  PIN csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END csb1
  PIN dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END dout1[0]
  PIN dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END dout1[10]
  PIN dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END dout1[11]
  PIN dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END dout1[12]
  PIN dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 4.000 312.080 ;
    END
  END dout1[13]
  PIN dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END dout1[14]
  PIN dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END dout1[15]
  PIN dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.200 4.000 348.800 ;
    END
  END dout1[16]
  PIN dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END dout1[17]
  PIN dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END dout1[18]
  PIN dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END dout1[19]
  PIN dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END dout1[1]
  PIN dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END dout1[20]
  PIN dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 4.000 410.000 ;
    END
  END dout1[21]
  PIN dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END dout1[22]
  PIN dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.880 4.000 434.480 ;
    END
  END dout1[23]
  PIN dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.120 4.000 446.720 ;
    END
  END dout1[24]
  PIN dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 458.360 4.000 458.960 ;
    END
  END dout1[25]
  PIN dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END dout1[26]
  PIN dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END dout1[27]
  PIN dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.080 4.000 495.680 ;
    END
  END dout1[28]
  PIN dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END dout1[29]
  PIN dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END dout1[2]
  PIN dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.560 4.000 520.160 ;
    END
  END dout1[30]
  PIN dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.800 4.000 532.400 ;
    END
  END dout1[31]
  PIN dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END dout1[3]
  PIN dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END dout1[4]
  PIN dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END dout1[5]
  PIN dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END dout1[6]
  PIN dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END dout1[7]
  PIN dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END dout1[8]
  PIN dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END dout1[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 546.000 576.290 550.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 546.000 737.290 550.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 546.000 592.390 550.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.210 546.000 608.490 550.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.310 546.000 624.590 550.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.410 546.000 640.690 550.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.510 546.000 656.790 550.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.610 546.000 672.890 550.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.710 546.000 688.990 550.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.810 546.000 705.090 550.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.910 546.000 721.190 550.000 ;
    END
  END io_oeb[9]
  PIN io_wbs_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END io_wbs_ack
  PIN io_wbs_adr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END io_wbs_adr[0]
  PIN io_wbs_adr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
    END
  END io_wbs_adr[10]
  PIN io_wbs_adr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END io_wbs_adr[11]
  PIN io_wbs_adr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 4.000 ;
    END
  END io_wbs_adr[12]
  PIN io_wbs_adr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 0.000 337.090 4.000 ;
    END
  END io_wbs_adr[13]
  PIN io_wbs_adr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END io_wbs_adr[14]
  PIN io_wbs_adr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END io_wbs_adr[15]
  PIN io_wbs_adr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 0.000 399.190 4.000 ;
    END
  END io_wbs_adr[16]
  PIN io_wbs_adr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.610 0.000 419.890 4.000 ;
    END
  END io_wbs_adr[17]
  PIN io_wbs_adr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 0.000 440.590 4.000 ;
    END
  END io_wbs_adr[18]
  PIN io_wbs_adr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 4.000 ;
    END
  END io_wbs_adr[19]
  PIN io_wbs_adr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END io_wbs_adr[1]
  PIN io_wbs_adr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 0.000 481.990 4.000 ;
    END
  END io_wbs_adr[20]
  PIN io_wbs_adr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END io_wbs_adr[21]
  PIN io_wbs_adr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.110 0.000 523.390 4.000 ;
    END
  END io_wbs_adr[22]
  PIN io_wbs_adr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 0.000 544.090 4.000 ;
    END
  END io_wbs_adr[23]
  PIN io_wbs_adr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 0.000 564.790 4.000 ;
    END
  END io_wbs_adr[24]
  PIN io_wbs_adr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 4.000 ;
    END
  END io_wbs_adr[25]
  PIN io_wbs_adr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 0.000 606.190 4.000 ;
    END
  END io_wbs_adr[26]
  PIN io_wbs_adr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.610 0.000 626.890 4.000 ;
    END
  END io_wbs_adr[27]
  PIN io_wbs_adr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 0.000 647.590 4.000 ;
    END
  END io_wbs_adr[28]
  PIN io_wbs_adr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.010 0.000 668.290 4.000 ;
    END
  END io_wbs_adr[29]
  PIN io_wbs_adr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END io_wbs_adr[2]
  PIN io_wbs_adr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.710 0.000 688.990 4.000 ;
    END
  END io_wbs_adr[30]
  PIN io_wbs_adr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.410 0.000 709.690 4.000 ;
    END
  END io_wbs_adr[31]
  PIN io_wbs_adr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END io_wbs_adr[3]
  PIN io_wbs_adr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END io_wbs_adr[4]
  PIN io_wbs_adr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END io_wbs_adr[5]
  PIN io_wbs_adr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END io_wbs_adr[6]
  PIN io_wbs_adr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END io_wbs_adr[7]
  PIN io_wbs_adr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 0.000 233.590 4.000 ;
    END
  END io_wbs_adr[8]
  PIN io_wbs_adr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END io_wbs_adr[9]
  PIN io_wbs_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END io_wbs_clk
  PIN io_wbs_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END io_wbs_cyc
  PIN io_wbs_datrd[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END io_wbs_datrd[0]
  PIN io_wbs_datrd[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 4.000 ;
    END
  END io_wbs_datrd[10]
  PIN io_wbs_datrd[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 4.000 ;
    END
  END io_wbs_datrd[11]
  PIN io_wbs_datrd[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 4.000 ;
    END
  END io_wbs_datrd[12]
  PIN io_wbs_datrd[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 4.000 ;
    END
  END io_wbs_datrd[13]
  PIN io_wbs_datrd[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END io_wbs_datrd[14]
  PIN io_wbs_datrd[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 0.000 385.390 4.000 ;
    END
  END io_wbs_datrd[15]
  PIN io_wbs_datrd[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END io_wbs_datrd[16]
  PIN io_wbs_datrd[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 0.000 426.790 4.000 ;
    END
  END io_wbs_datrd[17]
  PIN io_wbs_datrd[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 0.000 447.490 4.000 ;
    END
  END io_wbs_datrd[18]
  PIN io_wbs_datrd[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 0.000 468.190 4.000 ;
    END
  END io_wbs_datrd[19]
  PIN io_wbs_datrd[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 4.000 ;
    END
  END io_wbs_datrd[1]
  PIN io_wbs_datrd[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 0.000 488.890 4.000 ;
    END
  END io_wbs_datrd[20]
  PIN io_wbs_datrd[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 0.000 509.590 4.000 ;
    END
  END io_wbs_datrd[21]
  PIN io_wbs_datrd[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 0.000 530.290 4.000 ;
    END
  END io_wbs_datrd[22]
  PIN io_wbs_datrd[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 0.000 550.990 4.000 ;
    END
  END io_wbs_datrd[23]
  PIN io_wbs_datrd[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 0.000 571.690 4.000 ;
    END
  END io_wbs_datrd[24]
  PIN io_wbs_datrd[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 0.000 592.390 4.000 ;
    END
  END io_wbs_datrd[25]
  PIN io_wbs_datrd[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 0.000 613.090 4.000 ;
    END
  END io_wbs_datrd[26]
  PIN io_wbs_datrd[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.510 0.000 633.790 4.000 ;
    END
  END io_wbs_datrd[27]
  PIN io_wbs_datrd[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.210 0.000 654.490 4.000 ;
    END
  END io_wbs_datrd[28]
  PIN io_wbs_datrd[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 0.000 675.190 4.000 ;
    END
  END io_wbs_datrd[29]
  PIN io_wbs_datrd[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END io_wbs_datrd[2]
  PIN io_wbs_datrd[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END io_wbs_datrd[30]
  PIN io_wbs_datrd[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.310 0.000 716.590 4.000 ;
    END
  END io_wbs_datrd[31]
  PIN io_wbs_datrd[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END io_wbs_datrd[3]
  PIN io_wbs_datrd[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END io_wbs_datrd[4]
  PIN io_wbs_datrd[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 4.000 ;
    END
  END io_wbs_datrd[5]
  PIN io_wbs_datrd[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END io_wbs_datrd[6]
  PIN io_wbs_datrd[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 0.000 219.790 4.000 ;
    END
  END io_wbs_datrd[7]
  PIN io_wbs_datrd[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 4.000 ;
    END
  END io_wbs_datrd[8]
  PIN io_wbs_datrd[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END io_wbs_datrd[9]
  PIN io_wbs_datwr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 4.000 ;
    END
  END io_wbs_datwr[0]
  PIN io_wbs_datwr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END io_wbs_datwr[10]
  PIN io_wbs_datwr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END io_wbs_datwr[11]
  PIN io_wbs_datwr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 0.000 330.190 4.000 ;
    END
  END io_wbs_datwr[12]
  PIN io_wbs_datwr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END io_wbs_datwr[13]
  PIN io_wbs_datwr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 0.000 371.590 4.000 ;
    END
  END io_wbs_datwr[14]
  PIN io_wbs_datwr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END io_wbs_datwr[15]
  PIN io_wbs_datwr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 0.000 412.990 4.000 ;
    END
  END io_wbs_datwr[16]
  PIN io_wbs_datwr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 0.000 433.690 4.000 ;
    END
  END io_wbs_datwr[17]
  PIN io_wbs_datwr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END io_wbs_datwr[18]
  PIN io_wbs_datwr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.810 0.000 475.090 4.000 ;
    END
  END io_wbs_datwr[19]
  PIN io_wbs_datwr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END io_wbs_datwr[1]
  PIN io_wbs_datwr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 0.000 495.790 4.000 ;
    END
  END io_wbs_datwr[20]
  PIN io_wbs_datwr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 0.000 516.490 4.000 ;
    END
  END io_wbs_datwr[21]
  PIN io_wbs_datwr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 0.000 537.190 4.000 ;
    END
  END io_wbs_datwr[22]
  PIN io_wbs_datwr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.610 0.000 557.890 4.000 ;
    END
  END io_wbs_datwr[23]
  PIN io_wbs_datwr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 0.000 578.590 4.000 ;
    END
  END io_wbs_datwr[24]
  PIN io_wbs_datwr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END io_wbs_datwr[25]
  PIN io_wbs_datwr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 0.000 619.990 4.000 ;
    END
  END io_wbs_datwr[26]
  PIN io_wbs_datwr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.410 0.000 640.690 4.000 ;
    END
  END io_wbs_datwr[27]
  PIN io_wbs_datwr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.110 0.000 661.390 4.000 ;
    END
  END io_wbs_datwr[28]
  PIN io_wbs_datwr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.810 0.000 682.090 4.000 ;
    END
  END io_wbs_datwr[29]
  PIN io_wbs_datwr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END io_wbs_datwr[2]
  PIN io_wbs_datwr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 0.000 702.790 4.000 ;
    END
  END io_wbs_datwr[30]
  PIN io_wbs_datwr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.210 0.000 723.490 4.000 ;
    END
  END io_wbs_datwr[31]
  PIN io_wbs_datwr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END io_wbs_datwr[3]
  PIN io_wbs_datwr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END io_wbs_datwr[4]
  PIN io_wbs_datwr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END io_wbs_datwr[5]
  PIN io_wbs_datwr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END io_wbs_datwr[6]
  PIN io_wbs_datwr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END io_wbs_datwr[7]
  PIN io_wbs_datwr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 4.000 ;
    END
  END io_wbs_datwr[8]
  PIN io_wbs_datwr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 4.000 ;
    END
  END io_wbs_datwr[9]
  PIN io_wbs_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END io_wbs_rst
  PIN io_wbs_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END io_wbs_stb
  PIN io_wbs_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END io_wbs_we
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 538.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 538.800 ;
    END
  END vssd1
  PIN wfg_drive_pat_dout_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 546.000 61.090 550.000 ;
    END
  END wfg_drive_pat_dout_o[0]
  PIN wfg_drive_pat_dout_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 546.000 222.090 550.000 ;
    END
  END wfg_drive_pat_dout_o[10]
  PIN wfg_drive_pat_dout_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 546.000 238.190 550.000 ;
    END
  END wfg_drive_pat_dout_o[11]
  PIN wfg_drive_pat_dout_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 546.000 254.290 550.000 ;
    END
  END wfg_drive_pat_dout_o[12]
  PIN wfg_drive_pat_dout_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 546.000 270.390 550.000 ;
    END
  END wfg_drive_pat_dout_o[13]
  PIN wfg_drive_pat_dout_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 546.000 286.490 550.000 ;
    END
  END wfg_drive_pat_dout_o[14]
  PIN wfg_drive_pat_dout_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 546.000 302.590 550.000 ;
    END
  END wfg_drive_pat_dout_o[15]
  PIN wfg_drive_pat_dout_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 546.000 318.690 550.000 ;
    END
  END wfg_drive_pat_dout_o[16]
  PIN wfg_drive_pat_dout_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.510 546.000 334.790 550.000 ;
    END
  END wfg_drive_pat_dout_o[17]
  PIN wfg_drive_pat_dout_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 546.000 350.890 550.000 ;
    END
  END wfg_drive_pat_dout_o[18]
  PIN wfg_drive_pat_dout_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 546.000 366.990 550.000 ;
    END
  END wfg_drive_pat_dout_o[19]
  PIN wfg_drive_pat_dout_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 546.000 77.190 550.000 ;
    END
  END wfg_drive_pat_dout_o[1]
  PIN wfg_drive_pat_dout_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 546.000 383.090 550.000 ;
    END
  END wfg_drive_pat_dout_o[20]
  PIN wfg_drive_pat_dout_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 546.000 399.190 550.000 ;
    END
  END wfg_drive_pat_dout_o[21]
  PIN wfg_drive_pat_dout_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.010 546.000 415.290 550.000 ;
    END
  END wfg_drive_pat_dout_o[22]
  PIN wfg_drive_pat_dout_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.110 546.000 431.390 550.000 ;
    END
  END wfg_drive_pat_dout_o[23]
  PIN wfg_drive_pat_dout_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 546.000 447.490 550.000 ;
    END
  END wfg_drive_pat_dout_o[24]
  PIN wfg_drive_pat_dout_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.310 546.000 463.590 550.000 ;
    END
  END wfg_drive_pat_dout_o[25]
  PIN wfg_drive_pat_dout_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 546.000 479.690 550.000 ;
    END
  END wfg_drive_pat_dout_o[26]
  PIN wfg_drive_pat_dout_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 546.000 495.790 550.000 ;
    END
  END wfg_drive_pat_dout_o[27]
  PIN wfg_drive_pat_dout_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.610 546.000 511.890 550.000 ;
    END
  END wfg_drive_pat_dout_o[28]
  PIN wfg_drive_pat_dout_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.710 546.000 527.990 550.000 ;
    END
  END wfg_drive_pat_dout_o[29]
  PIN wfg_drive_pat_dout_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 546.000 93.290 550.000 ;
    END
  END wfg_drive_pat_dout_o[2]
  PIN wfg_drive_pat_dout_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 546.000 544.090 550.000 ;
    END
  END wfg_drive_pat_dout_o[30]
  PIN wfg_drive_pat_dout_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.910 546.000 560.190 550.000 ;
    END
  END wfg_drive_pat_dout_o[31]
  PIN wfg_drive_pat_dout_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 546.000 109.390 550.000 ;
    END
  END wfg_drive_pat_dout_o[3]
  PIN wfg_drive_pat_dout_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 546.000 125.490 550.000 ;
    END
  END wfg_drive_pat_dout_o[4]
  PIN wfg_drive_pat_dout_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 546.000 141.590 550.000 ;
    END
  END wfg_drive_pat_dout_o[5]
  PIN wfg_drive_pat_dout_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 546.000 157.690 550.000 ;
    END
  END wfg_drive_pat_dout_o[6]
  PIN wfg_drive_pat_dout_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 546.000 173.790 550.000 ;
    END
  END wfg_drive_pat_dout_o[7]
  PIN wfg_drive_pat_dout_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 546.000 189.890 550.000 ;
    END
  END wfg_drive_pat_dout_o[8]
  PIN wfg_drive_pat_dout_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 546.000 205.990 550.000 ;
    END
  END wfg_drive_pat_dout_o[9]
  PIN wfg_drive_spi_cs_no
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 546.000 12.790 550.000 ;
    END
  END wfg_drive_spi_cs_no
  PIN wfg_drive_spi_sclk_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 546.000 28.890 550.000 ;
    END
  END wfg_drive_spi_sclk_o
  PIN wfg_drive_spi_sdo_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 546.000 44.990 550.000 ;
    END
  END wfg_drive_spi_sdo_o
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 744.280 538.645 ;
      LAYER met1 ;
        RECT 5.520 7.520 744.280 538.800 ;
      LAYER met2 ;
        RECT 6.990 545.720 12.230 546.000 ;
        RECT 13.070 545.720 28.330 546.000 ;
        RECT 29.170 545.720 44.430 546.000 ;
        RECT 45.270 545.720 60.530 546.000 ;
        RECT 61.370 545.720 76.630 546.000 ;
        RECT 77.470 545.720 92.730 546.000 ;
        RECT 93.570 545.720 108.830 546.000 ;
        RECT 109.670 545.720 124.930 546.000 ;
        RECT 125.770 545.720 141.030 546.000 ;
        RECT 141.870 545.720 157.130 546.000 ;
        RECT 157.970 545.720 173.230 546.000 ;
        RECT 174.070 545.720 189.330 546.000 ;
        RECT 190.170 545.720 205.430 546.000 ;
        RECT 206.270 545.720 221.530 546.000 ;
        RECT 222.370 545.720 237.630 546.000 ;
        RECT 238.470 545.720 253.730 546.000 ;
        RECT 254.570 545.720 269.830 546.000 ;
        RECT 270.670 545.720 285.930 546.000 ;
        RECT 286.770 545.720 302.030 546.000 ;
        RECT 302.870 545.720 318.130 546.000 ;
        RECT 318.970 545.720 334.230 546.000 ;
        RECT 335.070 545.720 350.330 546.000 ;
        RECT 351.170 545.720 366.430 546.000 ;
        RECT 367.270 545.720 382.530 546.000 ;
        RECT 383.370 545.720 398.630 546.000 ;
        RECT 399.470 545.720 414.730 546.000 ;
        RECT 415.570 545.720 430.830 546.000 ;
        RECT 431.670 545.720 446.930 546.000 ;
        RECT 447.770 545.720 463.030 546.000 ;
        RECT 463.870 545.720 479.130 546.000 ;
        RECT 479.970 545.720 495.230 546.000 ;
        RECT 496.070 545.720 511.330 546.000 ;
        RECT 512.170 545.720 527.430 546.000 ;
        RECT 528.270 545.720 543.530 546.000 ;
        RECT 544.370 545.720 559.630 546.000 ;
        RECT 560.470 545.720 575.730 546.000 ;
        RECT 576.570 545.720 591.830 546.000 ;
        RECT 592.670 545.720 607.930 546.000 ;
        RECT 608.770 545.720 624.030 546.000 ;
        RECT 624.870 545.720 640.130 546.000 ;
        RECT 640.970 545.720 656.230 546.000 ;
        RECT 657.070 545.720 672.330 546.000 ;
        RECT 673.170 545.720 688.430 546.000 ;
        RECT 689.270 545.720 704.530 546.000 ;
        RECT 705.370 545.720 720.630 546.000 ;
        RECT 721.470 545.720 736.730 546.000 ;
        RECT 737.570 545.720 738.660 546.000 ;
        RECT 6.990 4.280 738.660 545.720 ;
        RECT 6.990 4.000 26.030 4.280 ;
        RECT 26.870 4.000 32.930 4.280 ;
        RECT 33.770 4.000 39.830 4.280 ;
        RECT 40.670 4.000 46.730 4.280 ;
        RECT 47.570 4.000 53.630 4.280 ;
        RECT 54.470 4.000 60.530 4.280 ;
        RECT 61.370 4.000 67.430 4.280 ;
        RECT 68.270 4.000 74.330 4.280 ;
        RECT 75.170 4.000 81.230 4.280 ;
        RECT 82.070 4.000 88.130 4.280 ;
        RECT 88.970 4.000 95.030 4.280 ;
        RECT 95.870 4.000 101.930 4.280 ;
        RECT 102.770 4.000 108.830 4.280 ;
        RECT 109.670 4.000 115.730 4.280 ;
        RECT 116.570 4.000 122.630 4.280 ;
        RECT 123.470 4.000 129.530 4.280 ;
        RECT 130.370 4.000 136.430 4.280 ;
        RECT 137.270 4.000 143.330 4.280 ;
        RECT 144.170 4.000 150.230 4.280 ;
        RECT 151.070 4.000 157.130 4.280 ;
        RECT 157.970 4.000 164.030 4.280 ;
        RECT 164.870 4.000 170.930 4.280 ;
        RECT 171.770 4.000 177.830 4.280 ;
        RECT 178.670 4.000 184.730 4.280 ;
        RECT 185.570 4.000 191.630 4.280 ;
        RECT 192.470 4.000 198.530 4.280 ;
        RECT 199.370 4.000 205.430 4.280 ;
        RECT 206.270 4.000 212.330 4.280 ;
        RECT 213.170 4.000 219.230 4.280 ;
        RECT 220.070 4.000 226.130 4.280 ;
        RECT 226.970 4.000 233.030 4.280 ;
        RECT 233.870 4.000 239.930 4.280 ;
        RECT 240.770 4.000 246.830 4.280 ;
        RECT 247.670 4.000 253.730 4.280 ;
        RECT 254.570 4.000 260.630 4.280 ;
        RECT 261.470 4.000 267.530 4.280 ;
        RECT 268.370 4.000 274.430 4.280 ;
        RECT 275.270 4.000 281.330 4.280 ;
        RECT 282.170 4.000 288.230 4.280 ;
        RECT 289.070 4.000 295.130 4.280 ;
        RECT 295.970 4.000 302.030 4.280 ;
        RECT 302.870 4.000 308.930 4.280 ;
        RECT 309.770 4.000 315.830 4.280 ;
        RECT 316.670 4.000 322.730 4.280 ;
        RECT 323.570 4.000 329.630 4.280 ;
        RECT 330.470 4.000 336.530 4.280 ;
        RECT 337.370 4.000 343.430 4.280 ;
        RECT 344.270 4.000 350.330 4.280 ;
        RECT 351.170 4.000 357.230 4.280 ;
        RECT 358.070 4.000 364.130 4.280 ;
        RECT 364.970 4.000 371.030 4.280 ;
        RECT 371.870 4.000 377.930 4.280 ;
        RECT 378.770 4.000 384.830 4.280 ;
        RECT 385.670 4.000 391.730 4.280 ;
        RECT 392.570 4.000 398.630 4.280 ;
        RECT 399.470 4.000 405.530 4.280 ;
        RECT 406.370 4.000 412.430 4.280 ;
        RECT 413.270 4.000 419.330 4.280 ;
        RECT 420.170 4.000 426.230 4.280 ;
        RECT 427.070 4.000 433.130 4.280 ;
        RECT 433.970 4.000 440.030 4.280 ;
        RECT 440.870 4.000 446.930 4.280 ;
        RECT 447.770 4.000 453.830 4.280 ;
        RECT 454.670 4.000 460.730 4.280 ;
        RECT 461.570 4.000 467.630 4.280 ;
        RECT 468.470 4.000 474.530 4.280 ;
        RECT 475.370 4.000 481.430 4.280 ;
        RECT 482.270 4.000 488.330 4.280 ;
        RECT 489.170 4.000 495.230 4.280 ;
        RECT 496.070 4.000 502.130 4.280 ;
        RECT 502.970 4.000 509.030 4.280 ;
        RECT 509.870 4.000 515.930 4.280 ;
        RECT 516.770 4.000 522.830 4.280 ;
        RECT 523.670 4.000 529.730 4.280 ;
        RECT 530.570 4.000 536.630 4.280 ;
        RECT 537.470 4.000 543.530 4.280 ;
        RECT 544.370 4.000 550.430 4.280 ;
        RECT 551.270 4.000 557.330 4.280 ;
        RECT 558.170 4.000 564.230 4.280 ;
        RECT 565.070 4.000 571.130 4.280 ;
        RECT 571.970 4.000 578.030 4.280 ;
        RECT 578.870 4.000 584.930 4.280 ;
        RECT 585.770 4.000 591.830 4.280 ;
        RECT 592.670 4.000 598.730 4.280 ;
        RECT 599.570 4.000 605.630 4.280 ;
        RECT 606.470 4.000 612.530 4.280 ;
        RECT 613.370 4.000 619.430 4.280 ;
        RECT 620.270 4.000 626.330 4.280 ;
        RECT 627.170 4.000 633.230 4.280 ;
        RECT 634.070 4.000 640.130 4.280 ;
        RECT 640.970 4.000 647.030 4.280 ;
        RECT 647.870 4.000 653.930 4.280 ;
        RECT 654.770 4.000 660.830 4.280 ;
        RECT 661.670 4.000 667.730 4.280 ;
        RECT 668.570 4.000 674.630 4.280 ;
        RECT 675.470 4.000 681.530 4.280 ;
        RECT 682.370 4.000 688.430 4.280 ;
        RECT 689.270 4.000 695.330 4.280 ;
        RECT 696.170 4.000 702.230 4.280 ;
        RECT 703.070 4.000 709.130 4.280 ;
        RECT 709.970 4.000 716.030 4.280 ;
        RECT 716.870 4.000 722.930 4.280 ;
        RECT 723.770 4.000 738.660 4.280 ;
      LAYER met3 ;
        RECT 4.000 532.800 713.855 538.725 ;
        RECT 4.400 531.400 713.855 532.800 ;
        RECT 4.000 520.560 713.855 531.400 ;
        RECT 4.400 519.160 713.855 520.560 ;
        RECT 4.000 508.320 713.855 519.160 ;
        RECT 4.400 506.920 713.855 508.320 ;
        RECT 4.000 496.080 713.855 506.920 ;
        RECT 4.400 494.680 713.855 496.080 ;
        RECT 4.000 483.840 713.855 494.680 ;
        RECT 4.400 482.440 713.855 483.840 ;
        RECT 4.000 471.600 713.855 482.440 ;
        RECT 4.400 470.200 713.855 471.600 ;
        RECT 4.000 459.360 713.855 470.200 ;
        RECT 4.400 457.960 713.855 459.360 ;
        RECT 4.000 447.120 713.855 457.960 ;
        RECT 4.400 445.720 713.855 447.120 ;
        RECT 4.000 434.880 713.855 445.720 ;
        RECT 4.400 433.480 713.855 434.880 ;
        RECT 4.000 422.640 713.855 433.480 ;
        RECT 4.400 421.240 713.855 422.640 ;
        RECT 4.000 410.400 713.855 421.240 ;
        RECT 4.400 409.000 713.855 410.400 ;
        RECT 4.000 398.160 713.855 409.000 ;
        RECT 4.400 396.760 713.855 398.160 ;
        RECT 4.000 385.920 713.855 396.760 ;
        RECT 4.400 384.520 713.855 385.920 ;
        RECT 4.000 373.680 713.855 384.520 ;
        RECT 4.400 372.280 713.855 373.680 ;
        RECT 4.000 361.440 713.855 372.280 ;
        RECT 4.400 360.040 713.855 361.440 ;
        RECT 4.000 349.200 713.855 360.040 ;
        RECT 4.400 347.800 713.855 349.200 ;
        RECT 4.000 336.960 713.855 347.800 ;
        RECT 4.400 335.560 713.855 336.960 ;
        RECT 4.000 324.720 713.855 335.560 ;
        RECT 4.400 323.320 713.855 324.720 ;
        RECT 4.000 312.480 713.855 323.320 ;
        RECT 4.400 311.080 713.855 312.480 ;
        RECT 4.000 300.240 713.855 311.080 ;
        RECT 4.400 298.840 713.855 300.240 ;
        RECT 4.000 288.000 713.855 298.840 ;
        RECT 4.400 286.600 713.855 288.000 ;
        RECT 4.000 275.760 713.855 286.600 ;
        RECT 4.400 274.360 713.855 275.760 ;
        RECT 4.000 263.520 713.855 274.360 ;
        RECT 4.400 262.120 713.855 263.520 ;
        RECT 4.000 251.280 713.855 262.120 ;
        RECT 4.400 249.880 713.855 251.280 ;
        RECT 4.000 239.040 713.855 249.880 ;
        RECT 4.400 237.640 713.855 239.040 ;
        RECT 4.000 226.800 713.855 237.640 ;
        RECT 4.400 225.400 713.855 226.800 ;
        RECT 4.000 214.560 713.855 225.400 ;
        RECT 4.400 213.160 713.855 214.560 ;
        RECT 4.000 202.320 713.855 213.160 ;
        RECT 4.400 200.920 713.855 202.320 ;
        RECT 4.000 190.080 713.855 200.920 ;
        RECT 4.400 188.680 713.855 190.080 ;
        RECT 4.000 177.840 713.855 188.680 ;
        RECT 4.400 176.440 713.855 177.840 ;
        RECT 4.000 165.600 713.855 176.440 ;
        RECT 4.400 164.200 713.855 165.600 ;
        RECT 4.000 153.360 713.855 164.200 ;
        RECT 4.400 151.960 713.855 153.360 ;
        RECT 4.000 141.120 713.855 151.960 ;
        RECT 4.400 139.720 713.855 141.120 ;
        RECT 4.000 128.880 713.855 139.720 ;
        RECT 4.400 127.480 713.855 128.880 ;
        RECT 4.000 116.640 713.855 127.480 ;
        RECT 4.400 115.240 713.855 116.640 ;
        RECT 4.000 104.400 713.855 115.240 ;
        RECT 4.400 103.000 713.855 104.400 ;
        RECT 4.000 92.160 713.855 103.000 ;
        RECT 4.400 90.760 713.855 92.160 ;
        RECT 4.000 79.920 713.855 90.760 ;
        RECT 4.400 78.520 713.855 79.920 ;
        RECT 4.000 67.680 713.855 78.520 ;
        RECT 4.400 66.280 713.855 67.680 ;
        RECT 4.000 55.440 713.855 66.280 ;
        RECT 4.400 54.040 713.855 55.440 ;
        RECT 4.000 43.200 713.855 54.040 ;
        RECT 4.400 41.800 713.855 43.200 ;
        RECT 4.000 30.960 713.855 41.800 ;
        RECT 4.400 29.560 713.855 30.960 ;
        RECT 4.000 18.720 713.855 29.560 ;
        RECT 4.400 17.320 713.855 18.720 ;
        RECT 4.000 10.715 713.855 17.320 ;
      LAYER met4 ;
        RECT 15.015 12.415 20.640 537.025 ;
        RECT 23.040 12.415 97.440 537.025 ;
        RECT 99.840 12.415 174.240 537.025 ;
        RECT 176.640 12.415 251.040 537.025 ;
        RECT 253.440 12.415 327.840 537.025 ;
        RECT 330.240 12.415 404.640 537.025 ;
        RECT 407.040 12.415 481.440 537.025 ;
        RECT 483.840 12.415 558.240 537.025 ;
        RECT 560.640 12.415 635.040 537.025 ;
        RECT 637.440 12.415 640.025 537.025 ;
  END
END wfg_top
END LIBRARY

